// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Mar 31 2025 15:38:36

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "cemf_module_64ch_main" view "INTERFACE"

module cemf_module_64ch_main (
    clock,
    start0,
    s0,
    intb0,
    dout1,
    csb1,
    sync_50hz,
    sdin1,
    sda,
    s1,
    intb1,
    dout0,
    csb0,
    serial_out_testing,
    sdin0,
    scl,
    s2,
    mcu_sclk,
    frame_sync,
    enable_config,
    elec_config_out,
    stop1,
    s3,
    rst_n,
    cemf_signal,
    trigger1,
    stop0,
    trigger0,
    stop_fpga2,
    sclk0,
    next_sequence,
    start1,
    sclk1,
    mcu_data);

    input clock;
    output start0;
    output s0;
    input intb0;
    output dout1;
    output csb1;
    input sync_50hz;
    input sdin1;
    inout sda;
    output s1;
    input intb1;
    output dout0;
    output csb0;
    output serial_out_testing;
    input sdin0;
    input scl;
    output s2;
    output mcu_sclk;
    output frame_sync;
    output enable_config;
    output elec_config_out;
    output stop1;
    output s3;
    input rst_n;
    input cemf_signal;
    input trigger1;
    output stop0;
    input trigger0;
    output stop_fpga2;
    output sclk0;
    output next_sequence;
    output start1;
    output sclk1;
    output mcu_data;

    wire N__67138;
    wire N__67137;
    wire N__67136;
    wire N__67129;
    wire N__67128;
    wire N__67127;
    wire N__67120;
    wire N__67119;
    wire N__67118;
    wire N__67111;
    wire N__67110;
    wire N__67109;
    wire N__67102;
    wire N__67101;
    wire N__67100;
    wire N__67093;
    wire N__67092;
    wire N__67091;
    wire N__67084;
    wire N__67083;
    wire N__67082;
    wire N__67075;
    wire N__67074;
    wire N__67073;
    wire N__67066;
    wire N__67065;
    wire N__67064;
    wire N__67057;
    wire N__67056;
    wire N__67055;
    wire N__67048;
    wire N__67047;
    wire N__67046;
    wire N__67039;
    wire N__67038;
    wire N__67037;
    wire N__67030;
    wire N__67029;
    wire N__67028;
    wire N__67021;
    wire N__67020;
    wire N__67019;
    wire N__67012;
    wire N__67011;
    wire N__67010;
    wire N__67003;
    wire N__67002;
    wire N__67001;
    wire N__66994;
    wire N__66993;
    wire N__66992;
    wire N__66985;
    wire N__66984;
    wire N__66983;
    wire N__66976;
    wire N__66975;
    wire N__66974;
    wire N__66967;
    wire N__66966;
    wire N__66965;
    wire N__66958;
    wire N__66957;
    wire N__66956;
    wire N__66949;
    wire N__66948;
    wire N__66947;
    wire N__66940;
    wire N__66939;
    wire N__66938;
    wire N__66931;
    wire N__66930;
    wire N__66929;
    wire N__66922;
    wire N__66921;
    wire N__66920;
    wire N__66913;
    wire N__66912;
    wire N__66911;
    wire N__66904;
    wire N__66903;
    wire N__66902;
    wire N__66895;
    wire N__66894;
    wire N__66893;
    wire N__66886;
    wire N__66885;
    wire N__66884;
    wire N__66867;
    wire N__66866;
    wire N__66863;
    wire N__66860;
    wire N__66857;
    wire N__66854;
    wire N__66853;
    wire N__66852;
    wire N__66851;
    wire N__66850;
    wire N__66847;
    wire N__66844;
    wire N__66839;
    wire N__66834;
    wire N__66825;
    wire N__66822;
    wire N__66819;
    wire N__66816;
    wire N__66815;
    wire N__66814;
    wire N__66813;
    wire N__66806;
    wire N__66803;
    wire N__66800;
    wire N__66799;
    wire N__66798;
    wire N__66795;
    wire N__66794;
    wire N__66791;
    wire N__66790;
    wire N__66789;
    wire N__66788;
    wire N__66787;
    wire N__66784;
    wire N__66781;
    wire N__66780;
    wire N__66779;
    wire N__66776;
    wire N__66773;
    wire N__66770;
    wire N__66769;
    wire N__66764;
    wire N__66759;
    wire N__66756;
    wire N__66755;
    wire N__66752;
    wire N__66747;
    wire N__66744;
    wire N__66739;
    wire N__66736;
    wire N__66731;
    wire N__66728;
    wire N__66725;
    wire N__66720;
    wire N__66715;
    wire N__66708;
    wire N__66699;
    wire N__66696;
    wire N__66693;
    wire N__66692;
    wire N__66691;
    wire N__66688;
    wire N__66687;
    wire N__66684;
    wire N__66681;
    wire N__66680;
    wire N__66677;
    wire N__66676;
    wire N__66675;
    wire N__66674;
    wire N__66673;
    wire N__66670;
    wire N__66665;
    wire N__66662;
    wire N__66659;
    wire N__66658;
    wire N__66655;
    wire N__66654;
    wire N__66653;
    wire N__66650;
    wire N__66645;
    wire N__66640;
    wire N__66637;
    wire N__66634;
    wire N__66627;
    wire N__66624;
    wire N__66609;
    wire N__66608;
    wire N__66607;
    wire N__66604;
    wire N__66603;
    wire N__66602;
    wire N__66599;
    wire N__66594;
    wire N__66593;
    wire N__66590;
    wire N__66587;
    wire N__66582;
    wire N__66579;
    wire N__66574;
    wire N__66571;
    wire N__66568;
    wire N__66561;
    wire N__66560;
    wire N__66559;
    wire N__66556;
    wire N__66555;
    wire N__66554;
    wire N__66553;
    wire N__66552;
    wire N__66551;
    wire N__66550;
    wire N__66549;
    wire N__66548;
    wire N__66545;
    wire N__66542;
    wire N__66539;
    wire N__66536;
    wire N__66533;
    wire N__66522;
    wire N__66519;
    wire N__66504;
    wire N__66503;
    wire N__66502;
    wire N__66499;
    wire N__66498;
    wire N__66497;
    wire N__66496;
    wire N__66495;
    wire N__66494;
    wire N__66493;
    wire N__66492;
    wire N__66489;
    wire N__66486;
    wire N__66483;
    wire N__66478;
    wire N__66471;
    wire N__66466;
    wire N__66453;
    wire N__66450;
    wire N__66449;
    wire N__66446;
    wire N__66443;
    wire N__66440;
    wire N__66437;
    wire N__66432;
    wire N__66431;
    wire N__66428;
    wire N__66425;
    wire N__66420;
    wire N__66419;
    wire N__66416;
    wire N__66413;
    wire N__66412;
    wire N__66411;
    wire N__66410;
    wire N__66407;
    wire N__66402;
    wire N__66397;
    wire N__66394;
    wire N__66389;
    wire N__66384;
    wire N__66383;
    wire N__66382;
    wire N__66379;
    wire N__66378;
    wire N__66377;
    wire N__66376;
    wire N__66375;
    wire N__66370;
    wire N__66367;
    wire N__66364;
    wire N__66361;
    wire N__66356;
    wire N__66353;
    wire N__66346;
    wire N__66339;
    wire N__66336;
    wire N__66333;
    wire N__66330;
    wire N__66329;
    wire N__66328;
    wire N__66327;
    wire N__66326;
    wire N__66325;
    wire N__66324;
    wire N__66321;
    wire N__66312;
    wire N__66309;
    wire N__66306;
    wire N__66303;
    wire N__66300;
    wire N__66291;
    wire N__66290;
    wire N__66287;
    wire N__66284;
    wire N__66279;
    wire N__66276;
    wire N__66275;
    wire N__66274;
    wire N__66273;
    wire N__66268;
    wire N__66265;
    wire N__66264;
    wire N__66261;
    wire N__66256;
    wire N__66255;
    wire N__66252;
    wire N__66251;
    wire N__66248;
    wire N__66245;
    wire N__66244;
    wire N__66243;
    wire N__66240;
    wire N__66237;
    wire N__66234;
    wire N__66229;
    wire N__66226;
    wire N__66223;
    wire N__66220;
    wire N__66215;
    wire N__66210;
    wire N__66201;
    wire N__66198;
    wire N__66195;
    wire N__66192;
    wire N__66191;
    wire N__66188;
    wire N__66187;
    wire N__66186;
    wire N__66185;
    wire N__66184;
    wire N__66175;
    wire N__66174;
    wire N__66169;
    wire N__66168;
    wire N__66167;
    wire N__66166;
    wire N__66165;
    wire N__66164;
    wire N__66163;
    wire N__66160;
    wire N__66157;
    wire N__66156;
    wire N__66155;
    wire N__66154;
    wire N__66151;
    wire N__66150;
    wire N__66143;
    wire N__66138;
    wire N__66135;
    wire N__66130;
    wire N__66129;
    wire N__66126;
    wire N__66125;
    wire N__66122;
    wire N__66119;
    wire N__66118;
    wire N__66115;
    wire N__66112;
    wire N__66111;
    wire N__66110;
    wire N__66109;
    wire N__66106;
    wire N__66105;
    wire N__66102;
    wire N__66099;
    wire N__66096;
    wire N__66095;
    wire N__66094;
    wire N__66093;
    wire N__66086;
    wire N__66079;
    wire N__66074;
    wire N__66067;
    wire N__66064;
    wire N__66061;
    wire N__66054;
    wire N__66051;
    wire N__66046;
    wire N__66041;
    wire N__66038;
    wire N__66021;
    wire N__66020;
    wire N__66019;
    wire N__66018;
    wire N__66017;
    wire N__66012;
    wire N__66009;
    wire N__66006;
    wire N__66003;
    wire N__65998;
    wire N__65991;
    wire N__65988;
    wire N__65987;
    wire N__65986;
    wire N__65985;
    wire N__65982;
    wire N__65979;
    wire N__65978;
    wire N__65975;
    wire N__65974;
    wire N__65971;
    wire N__65968;
    wire N__65965;
    wire N__65962;
    wire N__65957;
    wire N__65946;
    wire N__65945;
    wire N__65942;
    wire N__65939;
    wire N__65934;
    wire N__65933;
    wire N__65932;
    wire N__65927;
    wire N__65926;
    wire N__65923;
    wire N__65920;
    wire N__65915;
    wire N__65914;
    wire N__65909;
    wire N__65906;
    wire N__65903;
    wire N__65898;
    wire N__65897;
    wire N__65894;
    wire N__65893;
    wire N__65892;
    wire N__65889;
    wire N__65884;
    wire N__65881;
    wire N__65878;
    wire N__65873;
    wire N__65872;
    wire N__65871;
    wire N__65866;
    wire N__65861;
    wire N__65856;
    wire N__65853;
    wire N__65852;
    wire N__65849;
    wire N__65848;
    wire N__65845;
    wire N__65842;
    wire N__65839;
    wire N__65836;
    wire N__65829;
    wire N__65826;
    wire N__65823;
    wire N__65820;
    wire N__65819;
    wire N__65816;
    wire N__65813;
    wire N__65808;
    wire N__65807;
    wire N__65804;
    wire N__65801;
    wire N__65800;
    wire N__65797;
    wire N__65792;
    wire N__65787;
    wire N__65784;
    wire N__65783;
    wire N__65780;
    wire N__65777;
    wire N__65772;
    wire N__65769;
    wire N__65768;
    wire N__65767;
    wire N__65764;
    wire N__65761;
    wire N__65758;
    wire N__65755;
    wire N__65754;
    wire N__65753;
    wire N__65752;
    wire N__65751;
    wire N__65750;
    wire N__65749;
    wire N__65748;
    wire N__65747;
    wire N__65746;
    wire N__65745;
    wire N__65744;
    wire N__65743;
    wire N__65742;
    wire N__65741;
    wire N__65740;
    wire N__65739;
    wire N__65738;
    wire N__65737;
    wire N__65736;
    wire N__65735;
    wire N__65734;
    wire N__65733;
    wire N__65732;
    wire N__65731;
    wire N__65730;
    wire N__65729;
    wire N__65728;
    wire N__65727;
    wire N__65726;
    wire N__65725;
    wire N__65724;
    wire N__65723;
    wire N__65722;
    wire N__65721;
    wire N__65720;
    wire N__65719;
    wire N__65718;
    wire N__65717;
    wire N__65716;
    wire N__65715;
    wire N__65714;
    wire N__65713;
    wire N__65710;
    wire N__65707;
    wire N__65706;
    wire N__65705;
    wire N__65704;
    wire N__65703;
    wire N__65702;
    wire N__65701;
    wire N__65700;
    wire N__65699;
    wire N__65698;
    wire N__65697;
    wire N__65696;
    wire N__65695;
    wire N__65694;
    wire N__65693;
    wire N__65692;
    wire N__65691;
    wire N__65690;
    wire N__65689;
    wire N__65688;
    wire N__65687;
    wire N__65686;
    wire N__65685;
    wire N__65684;
    wire N__65683;
    wire N__65682;
    wire N__65681;
    wire N__65680;
    wire N__65679;
    wire N__65678;
    wire N__65677;
    wire N__65676;
    wire N__65675;
    wire N__65674;
    wire N__65673;
    wire N__65672;
    wire N__65671;
    wire N__65670;
    wire N__65669;
    wire N__65668;
    wire N__65667;
    wire N__65666;
    wire N__65665;
    wire N__65664;
    wire N__65663;
    wire N__65662;
    wire N__65661;
    wire N__65660;
    wire N__65659;
    wire N__65658;
    wire N__65657;
    wire N__65656;
    wire N__65655;
    wire N__65654;
    wire N__65653;
    wire N__65652;
    wire N__65651;
    wire N__65650;
    wire N__65649;
    wire N__65648;
    wire N__65647;
    wire N__65646;
    wire N__65645;
    wire N__65644;
    wire N__65643;
    wire N__65642;
    wire N__65641;
    wire N__65640;
    wire N__65639;
    wire N__65638;
    wire N__65637;
    wire N__65636;
    wire N__65635;
    wire N__65634;
    wire N__65633;
    wire N__65632;
    wire N__65631;
    wire N__65630;
    wire N__65629;
    wire N__65628;
    wire N__65627;
    wire N__65626;
    wire N__65625;
    wire N__65624;
    wire N__65623;
    wire N__65622;
    wire N__65621;
    wire N__65620;
    wire N__65619;
    wire N__65618;
    wire N__65617;
    wire N__65616;
    wire N__65615;
    wire N__65614;
    wire N__65613;
    wire N__65612;
    wire N__65611;
    wire N__65610;
    wire N__65609;
    wire N__65608;
    wire N__65607;
    wire N__65606;
    wire N__65605;
    wire N__65604;
    wire N__65603;
    wire N__65602;
    wire N__65601;
    wire N__65600;
    wire N__65599;
    wire N__65598;
    wire N__65597;
    wire N__65596;
    wire N__65595;
    wire N__65594;
    wire N__65593;
    wire N__65592;
    wire N__65591;
    wire N__65590;
    wire N__65589;
    wire N__65588;
    wire N__65587;
    wire N__65586;
    wire N__65585;
    wire N__65584;
    wire N__65583;
    wire N__65582;
    wire N__65581;
    wire N__65580;
    wire N__65579;
    wire N__65578;
    wire N__65577;
    wire N__65576;
    wire N__65575;
    wire N__65574;
    wire N__65573;
    wire N__65572;
    wire N__65571;
    wire N__65570;
    wire N__65569;
    wire N__65568;
    wire N__65567;
    wire N__65566;
    wire N__65565;
    wire N__65564;
    wire N__65563;
    wire N__65562;
    wire N__65561;
    wire N__65560;
    wire N__65559;
    wire N__65558;
    wire N__65557;
    wire N__65556;
    wire N__65555;
    wire N__65554;
    wire N__65553;
    wire N__65552;
    wire N__65551;
    wire N__65550;
    wire N__65549;
    wire N__65548;
    wire N__65547;
    wire N__65546;
    wire N__65545;
    wire N__65544;
    wire N__65543;
    wire N__65542;
    wire N__65541;
    wire N__65540;
    wire N__65539;
    wire N__65538;
    wire N__65537;
    wire N__65536;
    wire N__65535;
    wire N__65534;
    wire N__65533;
    wire N__65532;
    wire N__65531;
    wire N__65530;
    wire N__65529;
    wire N__65528;
    wire N__65527;
    wire N__65526;
    wire N__65525;
    wire N__65524;
    wire N__65523;
    wire N__65522;
    wire N__65521;
    wire N__65520;
    wire N__65519;
    wire N__65518;
    wire N__65517;
    wire N__65516;
    wire N__65515;
    wire N__65514;
    wire N__65513;
    wire N__65034;
    wire N__65031;
    wire N__65028;
    wire N__65027;
    wire N__65026;
    wire N__65025;
    wire N__65024;
    wire N__65023;
    wire N__65022;
    wire N__65021;
    wire N__65020;
    wire N__65019;
    wire N__65018;
    wire N__65017;
    wire N__65016;
    wire N__65015;
    wire N__65014;
    wire N__65013;
    wire N__65012;
    wire N__65011;
    wire N__65010;
    wire N__65009;
    wire N__65008;
    wire N__65007;
    wire N__65006;
    wire N__65005;
    wire N__65004;
    wire N__65003;
    wire N__65002;
    wire N__65001;
    wire N__65000;
    wire N__64999;
    wire N__64998;
    wire N__64997;
    wire N__64996;
    wire N__64995;
    wire N__64994;
    wire N__64993;
    wire N__64992;
    wire N__64991;
    wire N__64990;
    wire N__64989;
    wire N__64988;
    wire N__64987;
    wire N__64986;
    wire N__64985;
    wire N__64984;
    wire N__64983;
    wire N__64982;
    wire N__64981;
    wire N__64980;
    wire N__64979;
    wire N__64978;
    wire N__64977;
    wire N__64976;
    wire N__64975;
    wire N__64974;
    wire N__64973;
    wire N__64972;
    wire N__64971;
    wire N__64970;
    wire N__64969;
    wire N__64968;
    wire N__64967;
    wire N__64966;
    wire N__64965;
    wire N__64964;
    wire N__64963;
    wire N__64830;
    wire N__64827;
    wire N__64824;
    wire N__64821;
    wire N__64818;
    wire N__64815;
    wire N__64812;
    wire N__64809;
    wire N__64806;
    wire N__64803;
    wire N__64802;
    wire N__64801;
    wire N__64798;
    wire N__64795;
    wire N__64794;
    wire N__64791;
    wire N__64790;
    wire N__64789;
    wire N__64788;
    wire N__64787;
    wire N__64784;
    wire N__64781;
    wire N__64778;
    wire N__64775;
    wire N__64772;
    wire N__64769;
    wire N__64766;
    wire N__64763;
    wire N__64756;
    wire N__64751;
    wire N__64748;
    wire N__64737;
    wire N__64734;
    wire N__64731;
    wire N__64728;
    wire N__64725;
    wire N__64722;
    wire N__64721;
    wire N__64716;
    wire N__64713;
    wire N__64712;
    wire N__64709;
    wire N__64708;
    wire N__64707;
    wire N__64706;
    wire N__64705;
    wire N__64704;
    wire N__64701;
    wire N__64698;
    wire N__64697;
    wire N__64696;
    wire N__64693;
    wire N__64688;
    wire N__64687;
    wire N__64686;
    wire N__64685;
    wire N__64680;
    wire N__64679;
    wire N__64674;
    wire N__64669;
    wire N__64664;
    wire N__64657;
    wire N__64654;
    wire N__64651;
    wire N__64648;
    wire N__64641;
    wire N__64638;
    wire N__64629;
    wire N__64626;
    wire N__64623;
    wire N__64620;
    wire N__64617;
    wire N__64614;
    wire N__64611;
    wire N__64608;
    wire N__64605;
    wire N__64602;
    wire N__64599;
    wire N__64596;
    wire N__64593;
    wire N__64590;
    wire N__64587;
    wire N__64584;
    wire N__64583;
    wire N__64582;
    wire N__64581;
    wire N__64578;
    wire N__64577;
    wire N__64576;
    wire N__64575;
    wire N__64574;
    wire N__64573;
    wire N__64572;
    wire N__64571;
    wire N__64570;
    wire N__64561;
    wire N__64552;
    wire N__64551;
    wire N__64542;
    wire N__64539;
    wire N__64536;
    wire N__64533;
    wire N__64526;
    wire N__64523;
    wire N__64518;
    wire N__64515;
    wire N__64512;
    wire N__64509;
    wire N__64506;
    wire N__64503;
    wire N__64500;
    wire N__64497;
    wire N__64496;
    wire N__64493;
    wire N__64490;
    wire N__64485;
    wire N__64482;
    wire N__64479;
    wire N__64476;
    wire N__64473;
    wire N__64472;
    wire N__64469;
    wire N__64466;
    wire N__64465;
    wire N__64462;
    wire N__64459;
    wire N__64458;
    wire N__64457;
    wire N__64454;
    wire N__64449;
    wire N__64444;
    wire N__64437;
    wire N__64434;
    wire N__64433;
    wire N__64432;
    wire N__64429;
    wire N__64426;
    wire N__64425;
    wire N__64422;
    wire N__64421;
    wire N__64420;
    wire N__64417;
    wire N__64414;
    wire N__64411;
    wire N__64408;
    wire N__64407;
    wire N__64406;
    wire N__64401;
    wire N__64398;
    wire N__64393;
    wire N__64390;
    wire N__64385;
    wire N__64374;
    wire N__64371;
    wire N__64368;
    wire N__64365;
    wire N__64362;
    wire N__64359;
    wire N__64356;
    wire N__64355;
    wire N__64352;
    wire N__64349;
    wire N__64344;
    wire N__64343;
    wire N__64340;
    wire N__64337;
    wire N__64334;
    wire N__64331;
    wire N__64328;
    wire N__64323;
    wire N__64320;
    wire N__64317;
    wire N__64316;
    wire N__64313;
    wire N__64312;
    wire N__64309;
    wire N__64306;
    wire N__64303;
    wire N__64300;
    wire N__64299;
    wire N__64296;
    wire N__64293;
    wire N__64290;
    wire N__64287;
    wire N__64284;
    wire N__64281;
    wire N__64274;
    wire N__64269;
    wire N__64268;
    wire N__64267;
    wire N__64266;
    wire N__64265;
    wire N__64262;
    wire N__64261;
    wire N__64260;
    wire N__64259;
    wire N__64256;
    wire N__64253;
    wire N__64252;
    wire N__64251;
    wire N__64250;
    wire N__64249;
    wire N__64248;
    wire N__64247;
    wire N__64246;
    wire N__64245;
    wire N__64244;
    wire N__64243;
    wire N__64240;
    wire N__64237;
    wire N__64236;
    wire N__64235;
    wire N__64234;
    wire N__64231;
    wire N__64230;
    wire N__64229;
    wire N__64228;
    wire N__64225;
    wire N__64220;
    wire N__64219;
    wire N__64218;
    wire N__64217;
    wire N__64216;
    wire N__64215;
    wire N__64214;
    wire N__64213;
    wire N__64210;
    wire N__64209;
    wire N__64208;
    wire N__64207;
    wire N__64206;
    wire N__64205;
    wire N__64204;
    wire N__64203;
    wire N__64202;
    wire N__64201;
    wire N__64198;
    wire N__64193;
    wire N__64190;
    wire N__64175;
    wire N__64174;
    wire N__64173;
    wire N__64172;
    wire N__64169;
    wire N__64166;
    wire N__64161;
    wire N__64158;
    wire N__64157;
    wire N__64154;
    wire N__64153;
    wire N__64152;
    wire N__64149;
    wire N__64144;
    wire N__64139;
    wire N__64124;
    wire N__64121;
    wire N__64118;
    wire N__64117;
    wire N__64100;
    wire N__64095;
    wire N__64092;
    wire N__64089;
    wire N__64082;
    wire N__64081;
    wire N__64078;
    wire N__64075;
    wire N__64074;
    wire N__64073;
    wire N__64072;
    wire N__64071;
    wire N__64070;
    wire N__64069;
    wire N__64068;
    wire N__64067;
    wire N__64066;
    wire N__64061;
    wire N__64058;
    wire N__64055;
    wire N__64050;
    wire N__64043;
    wire N__64038;
    wire N__64033;
    wire N__64028;
    wire N__64021;
    wire N__64018;
    wire N__64013;
    wire N__64010;
    wire N__64007;
    wire N__64000;
    wire N__63991;
    wire N__63988;
    wire N__63977;
    wire N__63970;
    wire N__63951;
    wire N__63948;
    wire N__63945;
    wire N__63944;
    wire N__63941;
    wire N__63940;
    wire N__63939;
    wire N__63936;
    wire N__63933;
    wire N__63930;
    wire N__63927;
    wire N__63924;
    wire N__63923;
    wire N__63918;
    wire N__63915;
    wire N__63914;
    wire N__63911;
    wire N__63910;
    wire N__63909;
    wire N__63906;
    wire N__63905;
    wire N__63902;
    wire N__63899;
    wire N__63896;
    wire N__63893;
    wire N__63890;
    wire N__63887;
    wire N__63884;
    wire N__63881;
    wire N__63878;
    wire N__63873;
    wire N__63870;
    wire N__63867;
    wire N__63864;
    wire N__63859;
    wire N__63854;
    wire N__63851;
    wire N__63844;
    wire N__63837;
    wire N__63834;
    wire N__63831;
    wire N__63828;
    wire N__63827;
    wire N__63826;
    wire N__63823;
    wire N__63822;
    wire N__63819;
    wire N__63816;
    wire N__63813;
    wire N__63810;
    wire N__63809;
    wire N__63806;
    wire N__63803;
    wire N__63800;
    wire N__63799;
    wire N__63796;
    wire N__63793;
    wire N__63790;
    wire N__63789;
    wire N__63786;
    wire N__63785;
    wire N__63782;
    wire N__63779;
    wire N__63776;
    wire N__63775;
    wire N__63770;
    wire N__63767;
    wire N__63764;
    wire N__63761;
    wire N__63756;
    wire N__63753;
    wire N__63750;
    wire N__63747;
    wire N__63742;
    wire N__63739;
    wire N__63736;
    wire N__63733;
    wire N__63730;
    wire N__63727;
    wire N__63724;
    wire N__63719;
    wire N__63708;
    wire N__63705;
    wire N__63702;
    wire N__63701;
    wire N__63698;
    wire N__63697;
    wire N__63694;
    wire N__63691;
    wire N__63688;
    wire N__63687;
    wire N__63684;
    wire N__63681;
    wire N__63678;
    wire N__63677;
    wire N__63674;
    wire N__63671;
    wire N__63670;
    wire N__63665;
    wire N__63662;
    wire N__63661;
    wire N__63658;
    wire N__63657;
    wire N__63654;
    wire N__63651;
    wire N__63646;
    wire N__63645;
    wire N__63642;
    wire N__63639;
    wire N__63636;
    wire N__63633;
    wire N__63630;
    wire N__63627;
    wire N__63624;
    wire N__63621;
    wire N__63612;
    wire N__63609;
    wire N__63606;
    wire N__63603;
    wire N__63600;
    wire N__63591;
    wire N__63588;
    wire N__63585;
    wire N__63584;
    wire N__63583;
    wire N__63582;
    wire N__63581;
    wire N__63580;
    wire N__63577;
    wire N__63574;
    wire N__63569;
    wire N__63568;
    wire N__63565;
    wire N__63562;
    wire N__63559;
    wire N__63556;
    wire N__63553;
    wire N__63550;
    wire N__63547;
    wire N__63544;
    wire N__63543;
    wire N__63540;
    wire N__63537;
    wire N__63532;
    wire N__63527;
    wire N__63526;
    wire N__63523;
    wire N__63520;
    wire N__63517;
    wire N__63514;
    wire N__63511;
    wire N__63508;
    wire N__63503;
    wire N__63498;
    wire N__63489;
    wire N__63486;
    wire N__63483;
    wire N__63482;
    wire N__63481;
    wire N__63478;
    wire N__63477;
    wire N__63476;
    wire N__63473;
    wire N__63472;
    wire N__63471;
    wire N__63468;
    wire N__63467;
    wire N__63464;
    wire N__63461;
    wire N__63458;
    wire N__63455;
    wire N__63452;
    wire N__63449;
    wire N__63448;
    wire N__63445;
    wire N__63442;
    wire N__63439;
    wire N__63436;
    wire N__63433;
    wire N__63430;
    wire N__63427;
    wire N__63424;
    wire N__63421;
    wire N__63418;
    wire N__63407;
    wire N__63400;
    wire N__63397;
    wire N__63394;
    wire N__63391;
    wire N__63384;
    wire N__63383;
    wire N__63382;
    wire N__63381;
    wire N__63380;
    wire N__63379;
    wire N__63378;
    wire N__63377;
    wire N__63376;
    wire N__63359;
    wire N__63356;
    wire N__63355;
    wire N__63354;
    wire N__63353;
    wire N__63352;
    wire N__63351;
    wire N__63350;
    wire N__63349;
    wire N__63348;
    wire N__63347;
    wire N__63346;
    wire N__63345;
    wire N__63344;
    wire N__63343;
    wire N__63342;
    wire N__63341;
    wire N__63338;
    wire N__63327;
    wire N__63310;
    wire N__63303;
    wire N__63302;
    wire N__63301;
    wire N__63300;
    wire N__63299;
    wire N__63298;
    wire N__63297;
    wire N__63296;
    wire N__63295;
    wire N__63294;
    wire N__63293;
    wire N__63292;
    wire N__63285;
    wire N__63282;
    wire N__63281;
    wire N__63278;
    wire N__63275;
    wire N__63274;
    wire N__63273;
    wire N__63270;
    wire N__63255;
    wire N__63252;
    wire N__63247;
    wire N__63246;
    wire N__63243;
    wire N__63238;
    wire N__63235;
    wire N__63232;
    wire N__63231;
    wire N__63230;
    wire N__63225;
    wire N__63222;
    wire N__63219;
    wire N__63216;
    wire N__63211;
    wire N__63202;
    wire N__63199;
    wire N__63198;
    wire N__63197;
    wire N__63194;
    wire N__63191;
    wire N__63188;
    wire N__63183;
    wire N__63180;
    wire N__63175;
    wire N__63170;
    wire N__63163;
    wire N__63156;
    wire N__63153;
    wire N__63150;
    wire N__63149;
    wire N__63146;
    wire N__63145;
    wire N__63144;
    wire N__63141;
    wire N__63138;
    wire N__63135;
    wire N__63134;
    wire N__63131;
    wire N__63128;
    wire N__63123;
    wire N__63120;
    wire N__63119;
    wire N__63118;
    wire N__63115;
    wire N__63110;
    wire N__63107;
    wire N__63104;
    wire N__63103;
    wire N__63102;
    wire N__63099;
    wire N__63094;
    wire N__63091;
    wire N__63088;
    wire N__63083;
    wire N__63080;
    wire N__63077;
    wire N__63074;
    wire N__63071;
    wire N__63068;
    wire N__63065;
    wire N__63062;
    wire N__63059;
    wire N__63054;
    wire N__63045;
    wire N__63042;
    wire N__63039;
    wire N__63036;
    wire N__63033;
    wire N__63030;
    wire N__63029;
    wire N__63026;
    wire N__63025;
    wire N__63022;
    wire N__63019;
    wire N__63016;
    wire N__63015;
    wire N__63012;
    wire N__63007;
    wire N__63004;
    wire N__63003;
    wire N__63002;
    wire N__62999;
    wire N__62994;
    wire N__62991;
    wire N__62988;
    wire N__62985;
    wire N__62980;
    wire N__62977;
    wire N__62974;
    wire N__62971;
    wire N__62968;
    wire N__62961;
    wire N__62960;
    wire N__62959;
    wire N__62958;
    wire N__62957;
    wire N__62956;
    wire N__62955;
    wire N__62954;
    wire N__62953;
    wire N__62952;
    wire N__62951;
    wire N__62950;
    wire N__62949;
    wire N__62948;
    wire N__62947;
    wire N__62946;
    wire N__62945;
    wire N__62944;
    wire N__62943;
    wire N__62942;
    wire N__62941;
    wire N__62940;
    wire N__62939;
    wire N__62938;
    wire N__62937;
    wire N__62936;
    wire N__62935;
    wire N__62934;
    wire N__62933;
    wire N__62932;
    wire N__62931;
    wire N__62930;
    wire N__62929;
    wire N__62928;
    wire N__62927;
    wire N__62926;
    wire N__62925;
    wire N__62924;
    wire N__62923;
    wire N__62922;
    wire N__62921;
    wire N__62920;
    wire N__62919;
    wire N__62918;
    wire N__62917;
    wire N__62916;
    wire N__62915;
    wire N__62914;
    wire N__62913;
    wire N__62912;
    wire N__62911;
    wire N__62910;
    wire N__62909;
    wire N__62908;
    wire N__62907;
    wire N__62906;
    wire N__62905;
    wire N__62904;
    wire N__62903;
    wire N__62902;
    wire N__62901;
    wire N__62900;
    wire N__62899;
    wire N__62898;
    wire N__62897;
    wire N__62896;
    wire N__62895;
    wire N__62894;
    wire N__62893;
    wire N__62892;
    wire N__62891;
    wire N__62890;
    wire N__62889;
    wire N__62888;
    wire N__62887;
    wire N__62886;
    wire N__62885;
    wire N__62884;
    wire N__62883;
    wire N__62882;
    wire N__62881;
    wire N__62880;
    wire N__62879;
    wire N__62878;
    wire N__62877;
    wire N__62876;
    wire N__62875;
    wire N__62874;
    wire N__62873;
    wire N__62872;
    wire N__62871;
    wire N__62870;
    wire N__62869;
    wire N__62868;
    wire N__62867;
    wire N__62866;
    wire N__62865;
    wire N__62864;
    wire N__62863;
    wire N__62862;
    wire N__62861;
    wire N__62860;
    wire N__62859;
    wire N__62858;
    wire N__62857;
    wire N__62856;
    wire N__62855;
    wire N__62854;
    wire N__62853;
    wire N__62852;
    wire N__62851;
    wire N__62850;
    wire N__62849;
    wire N__62848;
    wire N__62847;
    wire N__62846;
    wire N__62845;
    wire N__62844;
    wire N__62843;
    wire N__62842;
    wire N__62841;
    wire N__62840;
    wire N__62839;
    wire N__62838;
    wire N__62837;
    wire N__62836;
    wire N__62835;
    wire N__62834;
    wire N__62833;
    wire N__62832;
    wire N__62831;
    wire N__62830;
    wire N__62829;
    wire N__62828;
    wire N__62827;
    wire N__62826;
    wire N__62825;
    wire N__62824;
    wire N__62823;
    wire N__62822;
    wire N__62821;
    wire N__62820;
    wire N__62819;
    wire N__62818;
    wire N__62817;
    wire N__62816;
    wire N__62815;
    wire N__62814;
    wire N__62813;
    wire N__62812;
    wire N__62811;
    wire N__62810;
    wire N__62809;
    wire N__62808;
    wire N__62807;
    wire N__62806;
    wire N__62805;
    wire N__62804;
    wire N__62487;
    wire N__62484;
    wire N__62481;
    wire N__62480;
    wire N__62479;
    wire N__62476;
    wire N__62473;
    wire N__62472;
    wire N__62469;
    wire N__62466;
    wire N__62463;
    wire N__62460;
    wire N__62457;
    wire N__62456;
    wire N__62455;
    wire N__62452;
    wire N__62447;
    wire N__62444;
    wire N__62441;
    wire N__62438;
    wire N__62433;
    wire N__62428;
    wire N__62421;
    wire N__62420;
    wire N__62417;
    wire N__62414;
    wire N__62411;
    wire N__62406;
    wire N__62403;
    wire N__62402;
    wire N__62399;
    wire N__62396;
    wire N__62393;
    wire N__62390;
    wire N__62387;
    wire N__62382;
    wire N__62379;
    wire N__62376;
    wire N__62373;
    wire N__62370;
    wire N__62369;
    wire N__62368;
    wire N__62367;
    wire N__62364;
    wire N__62361;
    wire N__62358;
    wire N__62357;
    wire N__62356;
    wire N__62353;
    wire N__62350;
    wire N__62347;
    wire N__62344;
    wire N__62341;
    wire N__62338;
    wire N__62337;
    wire N__62336;
    wire N__62333;
    wire N__62330;
    wire N__62327;
    wire N__62320;
    wire N__62317;
    wire N__62314;
    wire N__62311;
    wire N__62306;
    wire N__62303;
    wire N__62300;
    wire N__62295;
    wire N__62292;
    wire N__62289;
    wire N__62286;
    wire N__62281;
    wire N__62276;
    wire N__62271;
    wire N__62268;
    wire N__62265;
    wire N__62264;
    wire N__62263;
    wire N__62262;
    wire N__62261;
    wire N__62260;
    wire N__62259;
    wire N__62256;
    wire N__62253;
    wire N__62250;
    wire N__62247;
    wire N__62246;
    wire N__62243;
    wire N__62240;
    wire N__62237;
    wire N__62234;
    wire N__62231;
    wire N__62226;
    wire N__62223;
    wire N__62218;
    wire N__62215;
    wire N__62212;
    wire N__62209;
    wire N__62206;
    wire N__62197;
    wire N__62190;
    wire N__62187;
    wire N__62184;
    wire N__62183;
    wire N__62180;
    wire N__62179;
    wire N__62176;
    wire N__62173;
    wire N__62170;
    wire N__62169;
    wire N__62166;
    wire N__62165;
    wire N__62160;
    wire N__62157;
    wire N__62154;
    wire N__62151;
    wire N__62148;
    wire N__62147;
    wire N__62144;
    wire N__62139;
    wire N__62136;
    wire N__62133;
    wire N__62132;
    wire N__62129;
    wire N__62126;
    wire N__62125;
    wire N__62120;
    wire N__62117;
    wire N__62114;
    wire N__62111;
    wire N__62108;
    wire N__62105;
    wire N__62102;
    wire N__62097;
    wire N__62090;
    wire N__62087;
    wire N__62084;
    wire N__62079;
    wire N__62076;
    wire N__62073;
    wire N__62072;
    wire N__62071;
    wire N__62070;
    wire N__62067;
    wire N__62064;
    wire N__62061;
    wire N__62060;
    wire N__62059;
    wire N__62056;
    wire N__62051;
    wire N__62048;
    wire N__62045;
    wire N__62044;
    wire N__62041;
    wire N__62038;
    wire N__62033;
    wire N__62028;
    wire N__62025;
    wire N__62024;
    wire N__62019;
    wire N__62016;
    wire N__62013;
    wire N__62010;
    wire N__62007;
    wire N__62004;
    wire N__62001;
    wire N__61994;
    wire N__61989;
    wire N__61986;
    wire N__61983;
    wire N__61980;
    wire N__61977;
    wire N__61974;
    wire N__61971;
    wire N__61970;
    wire N__61969;
    wire N__61968;
    wire N__61965;
    wire N__61964;
    wire N__61963;
    wire N__61960;
    wire N__61959;
    wire N__61956;
    wire N__61953;
    wire N__61950;
    wire N__61947;
    wire N__61944;
    wire N__61943;
    wire N__61940;
    wire N__61937;
    wire N__61934;
    wire N__61931;
    wire N__61930;
    wire N__61927;
    wire N__61922;
    wire N__61919;
    wire N__61910;
    wire N__61907;
    wire N__61904;
    wire N__61901;
    wire N__61898;
    wire N__61895;
    wire N__61890;
    wire N__61887;
    wire N__61878;
    wire N__61875;
    wire N__61872;
    wire N__61871;
    wire N__61868;
    wire N__61867;
    wire N__61864;
    wire N__61863;
    wire N__61862;
    wire N__61861;
    wire N__61860;
    wire N__61859;
    wire N__61856;
    wire N__61853;
    wire N__61850;
    wire N__61847;
    wire N__61844;
    wire N__61841;
    wire N__61838;
    wire N__61835;
    wire N__61832;
    wire N__61827;
    wire N__61824;
    wire N__61821;
    wire N__61820;
    wire N__61817;
    wire N__61814;
    wire N__61811;
    wire N__61808;
    wire N__61803;
    wire N__61800;
    wire N__61797;
    wire N__61794;
    wire N__61791;
    wire N__61788;
    wire N__61785;
    wire N__61782;
    wire N__61779;
    wire N__61776;
    wire N__61773;
    wire N__61766;
    wire N__61759;
    wire N__61752;
    wire N__61749;
    wire N__61746;
    wire N__61745;
    wire N__61742;
    wire N__61739;
    wire N__61738;
    wire N__61737;
    wire N__61734;
    wire N__61731;
    wire N__61730;
    wire N__61729;
    wire N__61726;
    wire N__61723;
    wire N__61720;
    wire N__61719;
    wire N__61716;
    wire N__61713;
    wire N__61712;
    wire N__61711;
    wire N__61708;
    wire N__61705;
    wire N__61700;
    wire N__61697;
    wire N__61694;
    wire N__61691;
    wire N__61688;
    wire N__61685;
    wire N__61682;
    wire N__61675;
    wire N__61670;
    wire N__61667;
    wire N__61662;
    wire N__61659;
    wire N__61656;
    wire N__61647;
    wire N__61646;
    wire N__61645;
    wire N__61644;
    wire N__61641;
    wire N__61640;
    wire N__61639;
    wire N__61636;
    wire N__61633;
    wire N__61632;
    wire N__61631;
    wire N__61628;
    wire N__61625;
    wire N__61622;
    wire N__61619;
    wire N__61614;
    wire N__61613;
    wire N__61610;
    wire N__61607;
    wire N__61604;
    wire N__61599;
    wire N__61596;
    wire N__61593;
    wire N__61590;
    wire N__61587;
    wire N__61580;
    wire N__61575;
    wire N__61572;
    wire N__61569;
    wire N__61566;
    wire N__61559;
    wire N__61554;
    wire N__61551;
    wire N__61548;
    wire N__61547;
    wire N__61546;
    wire N__61545;
    wire N__61544;
    wire N__61541;
    wire N__61538;
    wire N__61535;
    wire N__61532;
    wire N__61531;
    wire N__61530;
    wire N__61527;
    wire N__61526;
    wire N__61525;
    wire N__61522;
    wire N__61517;
    wire N__61514;
    wire N__61511;
    wire N__61508;
    wire N__61505;
    wire N__61502;
    wire N__61499;
    wire N__61494;
    wire N__61491;
    wire N__61486;
    wire N__61483;
    wire N__61478;
    wire N__61473;
    wire N__61468;
    wire N__61461;
    wire N__61458;
    wire N__61455;
    wire N__61452;
    wire N__61449;
    wire N__61448;
    wire N__61447;
    wire N__61444;
    wire N__61441;
    wire N__61438;
    wire N__61437;
    wire N__61436;
    wire N__61435;
    wire N__61434;
    wire N__61431;
    wire N__61428;
    wire N__61425;
    wire N__61422;
    wire N__61421;
    wire N__61418;
    wire N__61415;
    wire N__61412;
    wire N__61407;
    wire N__61406;
    wire N__61401;
    wire N__61398;
    wire N__61395;
    wire N__61390;
    wire N__61387;
    wire N__61384;
    wire N__61381;
    wire N__61376;
    wire N__61371;
    wire N__61362;
    wire N__61359;
    wire N__61356;
    wire N__61355;
    wire N__61354;
    wire N__61353;
    wire N__61352;
    wire N__61349;
    wire N__61348;
    wire N__61345;
    wire N__61342;
    wire N__61339;
    wire N__61336;
    wire N__61333;
    wire N__61330;
    wire N__61327;
    wire N__61320;
    wire N__61319;
    wire N__61318;
    wire N__61311;
    wire N__61310;
    wire N__61307;
    wire N__61304;
    wire N__61301;
    wire N__61298;
    wire N__61295;
    wire N__61290;
    wire N__61287;
    wire N__61284;
    wire N__61281;
    wire N__61276;
    wire N__61273;
    wire N__61270;
    wire N__61267;
    wire N__61260;
    wire N__61257;
    wire N__61254;
    wire N__61253;
    wire N__61252;
    wire N__61249;
    wire N__61248;
    wire N__61247;
    wire N__61246;
    wire N__61243;
    wire N__61242;
    wire N__61239;
    wire N__61236;
    wire N__61233;
    wire N__61230;
    wire N__61229;
    wire N__61226;
    wire N__61223;
    wire N__61220;
    wire N__61217;
    wire N__61212;
    wire N__61209;
    wire N__61206;
    wire N__61203;
    wire N__61200;
    wire N__61197;
    wire N__61194;
    wire N__61193;
    wire N__61188;
    wire N__61185;
    wire N__61182;
    wire N__61177;
    wire N__61174;
    wire N__61171;
    wire N__61166;
    wire N__61163;
    wire N__61158;
    wire N__61155;
    wire N__61152;
    wire N__61149;
    wire N__61146;
    wire N__61137;
    wire N__61134;
    wire N__61131;
    wire N__61130;
    wire N__61127;
    wire N__61126;
    wire N__61125;
    wire N__61124;
    wire N__61121;
    wire N__61118;
    wire N__61117;
    wire N__61114;
    wire N__61113;
    wire N__61110;
    wire N__61107;
    wire N__61104;
    wire N__61103;
    wire N__61100;
    wire N__61097;
    wire N__61094;
    wire N__61091;
    wire N__61088;
    wire N__61085;
    wire N__61082;
    wire N__61079;
    wire N__61076;
    wire N__61073;
    wire N__61070;
    wire N__61063;
    wire N__61060;
    wire N__61057;
    wire N__61054;
    wire N__61051;
    wire N__61048;
    wire N__61045;
    wire N__61038;
    wire N__61033;
    wire N__61026;
    wire N__61023;
    wire N__61020;
    wire N__61019;
    wire N__61018;
    wire N__61015;
    wire N__61014;
    wire N__61013;
    wire N__61010;
    wire N__61007;
    wire N__61004;
    wire N__61001;
    wire N__61000;
    wire N__60997;
    wire N__60994;
    wire N__60991;
    wire N__60988;
    wire N__60985;
    wire N__60982;
    wire N__60981;
    wire N__60980;
    wire N__60977;
    wire N__60972;
    wire N__60967;
    wire N__60964;
    wire N__60961;
    wire N__60958;
    wire N__60955;
    wire N__60952;
    wire N__60949;
    wire N__60946;
    wire N__60939;
    wire N__60934;
    wire N__60927;
    wire N__60924;
    wire N__60921;
    wire N__60918;
    wire N__60915;
    wire N__60914;
    wire N__60913;
    wire N__60912;
    wire N__60909;
    wire N__60906;
    wire N__60905;
    wire N__60902;
    wire N__60901;
    wire N__60898;
    wire N__60897;
    wire N__60892;
    wire N__60889;
    wire N__60886;
    wire N__60883;
    wire N__60880;
    wire N__60877;
    wire N__60872;
    wire N__60869;
    wire N__60866;
    wire N__60863;
    wire N__60860;
    wire N__60857;
    wire N__60850;
    wire N__60849;
    wire N__60846;
    wire N__60843;
    wire N__60840;
    wire N__60837;
    wire N__60834;
    wire N__60829;
    wire N__60822;
    wire N__60819;
    wire N__60816;
    wire N__60813;
    wire N__60810;
    wire N__60807;
    wire N__60806;
    wire N__60805;
    wire N__60802;
    wire N__60799;
    wire N__60798;
    wire N__60797;
    wire N__60794;
    wire N__60791;
    wire N__60788;
    wire N__60787;
    wire N__60786;
    wire N__60783;
    wire N__60780;
    wire N__60777;
    wire N__60776;
    wire N__60771;
    wire N__60768;
    wire N__60765;
    wire N__60762;
    wire N__60759;
    wire N__60756;
    wire N__60753;
    wire N__60746;
    wire N__60743;
    wire N__60740;
    wire N__60737;
    wire N__60734;
    wire N__60731;
    wire N__60728;
    wire N__60723;
    wire N__60714;
    wire N__60711;
    wire N__60710;
    wire N__60709;
    wire N__60706;
    wire N__60703;
    wire N__60700;
    wire N__60697;
    wire N__60694;
    wire N__60691;
    wire N__60688;
    wire N__60683;
    wire N__60678;
    wire N__60675;
    wire N__60672;
    wire N__60669;
    wire N__60666;
    wire N__60663;
    wire N__60660;
    wire N__60657;
    wire N__60654;
    wire N__60651;
    wire N__60648;
    wire N__60645;
    wire N__60642;
    wire N__60641;
    wire N__60640;
    wire N__60637;
    wire N__60634;
    wire N__60631;
    wire N__60626;
    wire N__60623;
    wire N__60618;
    wire N__60617;
    wire N__60616;
    wire N__60615;
    wire N__60614;
    wire N__60613;
    wire N__60612;
    wire N__60609;
    wire N__60606;
    wire N__60605;
    wire N__60604;
    wire N__60599;
    wire N__60598;
    wire N__60597;
    wire N__60592;
    wire N__60591;
    wire N__60590;
    wire N__60589;
    wire N__60586;
    wire N__60581;
    wire N__60578;
    wire N__60575;
    wire N__60572;
    wire N__60569;
    wire N__60566;
    wire N__60565;
    wire N__60562;
    wire N__60559;
    wire N__60558;
    wire N__60557;
    wire N__60552;
    wire N__60549;
    wire N__60544;
    wire N__60541;
    wire N__60540;
    wire N__60535;
    wire N__60532;
    wire N__60529;
    wire N__60524;
    wire N__60521;
    wire N__60518;
    wire N__60517;
    wire N__60516;
    wire N__60515;
    wire N__60512;
    wire N__60507;
    wire N__60504;
    wire N__60501;
    wire N__60496;
    wire N__60489;
    wire N__60486;
    wire N__60483;
    wire N__60478;
    wire N__60475;
    wire N__60474;
    wire N__60473;
    wire N__60472;
    wire N__60469;
    wire N__60464;
    wire N__60461;
    wire N__60456;
    wire N__60451;
    wire N__60448;
    wire N__60445;
    wire N__60440;
    wire N__60435;
    wire N__60430;
    wire N__60427;
    wire N__60420;
    wire N__60411;
    wire N__60408;
    wire N__60405;
    wire N__60402;
    wire N__60399;
    wire N__60396;
    wire N__60393;
    wire N__60390;
    wire N__60387;
    wire N__60386;
    wire N__60385;
    wire N__60384;
    wire N__60383;
    wire N__60382;
    wire N__60381;
    wire N__60380;
    wire N__60379;
    wire N__60378;
    wire N__60377;
    wire N__60376;
    wire N__60375;
    wire N__60374;
    wire N__60369;
    wire N__60364;
    wire N__60359;
    wire N__60358;
    wire N__60357;
    wire N__60356;
    wire N__60355;
    wire N__60354;
    wire N__60353;
    wire N__60350;
    wire N__60347;
    wire N__60346;
    wire N__60345;
    wire N__60340;
    wire N__60335;
    wire N__60330;
    wire N__60329;
    wire N__60328;
    wire N__60325;
    wire N__60320;
    wire N__60317;
    wire N__60312;
    wire N__60307;
    wire N__60304;
    wire N__60299;
    wire N__60294;
    wire N__60287;
    wire N__60282;
    wire N__60277;
    wire N__60272;
    wire N__60269;
    wire N__60266;
    wire N__60263;
    wire N__60260;
    wire N__60257;
    wire N__60254;
    wire N__60249;
    wire N__60246;
    wire N__60243;
    wire N__60240;
    wire N__60235;
    wire N__60230;
    wire N__60219;
    wire N__60216;
    wire N__60213;
    wire N__60210;
    wire N__60207;
    wire N__60206;
    wire N__60205;
    wire N__60204;
    wire N__60203;
    wire N__60202;
    wire N__60197;
    wire N__60196;
    wire N__60195;
    wire N__60194;
    wire N__60193;
    wire N__60188;
    wire N__60187;
    wire N__60186;
    wire N__60181;
    wire N__60178;
    wire N__60173;
    wire N__60168;
    wire N__60167;
    wire N__60166;
    wire N__60165;
    wire N__60164;
    wire N__60163;
    wire N__60162;
    wire N__60159;
    wire N__60158;
    wire N__60157;
    wire N__60152;
    wire N__60151;
    wire N__60150;
    wire N__60149;
    wire N__60148;
    wire N__60145;
    wire N__60138;
    wire N__60133;
    wire N__60128;
    wire N__60127;
    wire N__60122;
    wire N__60119;
    wire N__60114;
    wire N__60111;
    wire N__60106;
    wire N__60101;
    wire N__60098;
    wire N__60093;
    wire N__60090;
    wire N__60087;
    wire N__60084;
    wire N__60081;
    wire N__60078;
    wire N__60073;
    wire N__60070;
    wire N__60063;
    wire N__60060;
    wire N__60057;
    wire N__60054;
    wire N__60051;
    wire N__60046;
    wire N__60041;
    wire N__60030;
    wire N__60027;
    wire N__60024;
    wire N__60023;
    wire N__60022;
    wire N__60019;
    wire N__60018;
    wire N__60017;
    wire N__60016;
    wire N__60013;
    wire N__60010;
    wire N__60009;
    wire N__60006;
    wire N__60005;
    wire N__60004;
    wire N__60001;
    wire N__59998;
    wire N__59995;
    wire N__59994;
    wire N__59991;
    wire N__59988;
    wire N__59985;
    wire N__59984;
    wire N__59981;
    wire N__59978;
    wire N__59975;
    wire N__59972;
    wire N__59969;
    wire N__59966;
    wire N__59963;
    wire N__59958;
    wire N__59955;
    wire N__59952;
    wire N__59947;
    wire N__59944;
    wire N__59941;
    wire N__59940;
    wire N__59935;
    wire N__59932;
    wire N__59929;
    wire N__59926;
    wire N__59923;
    wire N__59920;
    wire N__59917;
    wire N__59914;
    wire N__59911;
    wire N__59906;
    wire N__59901;
    wire N__59896;
    wire N__59893;
    wire N__59888;
    wire N__59885;
    wire N__59882;
    wire N__59879;
    wire N__59874;
    wire N__59865;
    wire N__59864;
    wire N__59863;
    wire N__59860;
    wire N__59857;
    wire N__59854;
    wire N__59853;
    wire N__59852;
    wire N__59851;
    wire N__59850;
    wire N__59845;
    wire N__59844;
    wire N__59841;
    wire N__59838;
    wire N__59835;
    wire N__59834;
    wire N__59831;
    wire N__59828;
    wire N__59825;
    wire N__59822;
    wire N__59817;
    wire N__59814;
    wire N__59811;
    wire N__59808;
    wire N__59805;
    wire N__59802;
    wire N__59797;
    wire N__59794;
    wire N__59791;
    wire N__59788;
    wire N__59783;
    wire N__59780;
    wire N__59775;
    wire N__59772;
    wire N__59763;
    wire N__59760;
    wire N__59757;
    wire N__59754;
    wire N__59751;
    wire N__59748;
    wire N__59745;
    wire N__59742;
    wire N__59739;
    wire N__59736;
    wire N__59733;
    wire N__59730;
    wire N__59729;
    wire N__59728;
    wire N__59727;
    wire N__59726;
    wire N__59723;
    wire N__59720;
    wire N__59719;
    wire N__59718;
    wire N__59717;
    wire N__59716;
    wire N__59715;
    wire N__59714;
    wire N__59713;
    wire N__59712;
    wire N__59711;
    wire N__59710;
    wire N__59709;
    wire N__59708;
    wire N__59707;
    wire N__59706;
    wire N__59705;
    wire N__59704;
    wire N__59703;
    wire N__59702;
    wire N__59699;
    wire N__59698;
    wire N__59697;
    wire N__59696;
    wire N__59695;
    wire N__59690;
    wire N__59677;
    wire N__59676;
    wire N__59675;
    wire N__59674;
    wire N__59673;
    wire N__59672;
    wire N__59671;
    wire N__59654;
    wire N__59653;
    wire N__59652;
    wire N__59651;
    wire N__59650;
    wire N__59649;
    wire N__59648;
    wire N__59647;
    wire N__59646;
    wire N__59645;
    wire N__59644;
    wire N__59643;
    wire N__59642;
    wire N__59641;
    wire N__59640;
    wire N__59639;
    wire N__59638;
    wire N__59637;
    wire N__59636;
    wire N__59635;
    wire N__59634;
    wire N__59633;
    wire N__59632;
    wire N__59625;
    wire N__59608;
    wire N__59607;
    wire N__59606;
    wire N__59605;
    wire N__59604;
    wire N__59603;
    wire N__59602;
    wire N__59601;
    wire N__59600;
    wire N__59599;
    wire N__59598;
    wire N__59597;
    wire N__59596;
    wire N__59595;
    wire N__59594;
    wire N__59593;
    wire N__59592;
    wire N__59591;
    wire N__59590;
    wire N__59589;
    wire N__59588;
    wire N__59587;
    wire N__59582;
    wire N__59569;
    wire N__59566;
    wire N__59559;
    wire N__59558;
    wire N__59557;
    wire N__59556;
    wire N__59555;
    wire N__59554;
    wire N__59553;
    wire N__59552;
    wire N__59551;
    wire N__59550;
    wire N__59549;
    wire N__59548;
    wire N__59547;
    wire N__59546;
    wire N__59545;
    wire N__59544;
    wire N__59543;
    wire N__59542;
    wire N__59541;
    wire N__59524;
    wire N__59517;
    wire N__59516;
    wire N__59515;
    wire N__59514;
    wire N__59513;
    wire N__59512;
    wire N__59511;
    wire N__59510;
    wire N__59509;
    wire N__59508;
    wire N__59507;
    wire N__59506;
    wire N__59505;
    wire N__59504;
    wire N__59487;
    wire N__59482;
    wire N__59465;
    wire N__59460;
    wire N__59449;
    wire N__59448;
    wire N__59447;
    wire N__59446;
    wire N__59445;
    wire N__59444;
    wire N__59443;
    wire N__59442;
    wire N__59441;
    wire N__59440;
    wire N__59439;
    wire N__59438;
    wire N__59437;
    wire N__59436;
    wire N__59435;
    wire N__59434;
    wire N__59433;
    wire N__59432;
    wire N__59431;
    wire N__59430;
    wire N__59429;
    wire N__59428;
    wire N__59427;
    wire N__59426;
    wire N__59425;
    wire N__59424;
    wire N__59423;
    wire N__59422;
    wire N__59421;
    wire N__59420;
    wire N__59419;
    wire N__59418;
    wire N__59417;
    wire N__59416;
    wire N__59415;
    wire N__59414;
    wire N__59413;
    wire N__59412;
    wire N__59399;
    wire N__59394;
    wire N__59389;
    wire N__59388;
    wire N__59387;
    wire N__59386;
    wire N__59385;
    wire N__59384;
    wire N__59383;
    wire N__59382;
    wire N__59381;
    wire N__59374;
    wire N__59371;
    wire N__59368;
    wire N__59365;
    wire N__59348;
    wire N__59345;
    wire N__59342;
    wire N__59339;
    wire N__59336;
    wire N__59335;
    wire N__59334;
    wire N__59333;
    wire N__59328;
    wire N__59311;
    wire N__59308;
    wire N__59299;
    wire N__59294;
    wire N__59287;
    wire N__59284;
    wire N__59281;
    wire N__59278;
    wire N__59277;
    wire N__59276;
    wire N__59275;
    wire N__59272;
    wire N__59269;
    wire N__59262;
    wire N__59245;
    wire N__59240;
    wire N__59223;
    wire N__59216;
    wire N__59199;
    wire N__59194;
    wire N__59191;
    wire N__59190;
    wire N__59189;
    wire N__59188;
    wire N__59187;
    wire N__59186;
    wire N__59185;
    wire N__59184;
    wire N__59183;
    wire N__59180;
    wire N__59171;
    wire N__59166;
    wire N__59165;
    wire N__59164;
    wire N__59163;
    wire N__59162;
    wire N__59161;
    wire N__59160;
    wire N__59157;
    wire N__59150;
    wire N__59149;
    wire N__59148;
    wire N__59147;
    wire N__59146;
    wire N__59145;
    wire N__59144;
    wire N__59143;
    wire N__59142;
    wire N__59141;
    wire N__59140;
    wire N__59139;
    wire N__59134;
    wire N__59119;
    wire N__59106;
    wire N__59093;
    wire N__59090;
    wire N__59085;
    wire N__59082;
    wire N__59071;
    wire N__59068;
    wire N__59051;
    wire N__59046;
    wire N__59043;
    wire N__59038;
    wire N__59035;
    wire N__59032;
    wire N__59029;
    wire N__59026;
    wire N__59025;
    wire N__59024;
    wire N__59023;
    wire N__59020;
    wire N__59017;
    wire N__59016;
    wire N__59015;
    wire N__59014;
    wire N__59013;
    wire N__59012;
    wire N__59011;
    wire N__59010;
    wire N__58993;
    wire N__58988;
    wire N__58985;
    wire N__58978;
    wire N__58971;
    wire N__58964;
    wire N__58955;
    wire N__58940;
    wire N__58935;
    wire N__58926;
    wire N__58919;
    wire N__58916;
    wire N__58909;
    wire N__58902;
    wire N__58897;
    wire N__58884;
    wire N__58881;
    wire N__58880;
    wire N__58879;
    wire N__58876;
    wire N__58873;
    wire N__58870;
    wire N__58869;
    wire N__58868;
    wire N__58867;
    wire N__58862;
    wire N__58859;
    wire N__58856;
    wire N__58853;
    wire N__58850;
    wire N__58843;
    wire N__58840;
    wire N__58837;
    wire N__58834;
    wire N__58831;
    wire N__58828;
    wire N__58825;
    wire N__58818;
    wire N__58815;
    wire N__58812;
    wire N__58809;
    wire N__58806;
    wire N__58803;
    wire N__58800;
    wire N__58797;
    wire N__58796;
    wire N__58795;
    wire N__58792;
    wire N__58789;
    wire N__58788;
    wire N__58787;
    wire N__58784;
    wire N__58783;
    wire N__58780;
    wire N__58779;
    wire N__58776;
    wire N__58773;
    wire N__58770;
    wire N__58767;
    wire N__58766;
    wire N__58763;
    wire N__58760;
    wire N__58757;
    wire N__58750;
    wire N__58749;
    wire N__58746;
    wire N__58743;
    wire N__58738;
    wire N__58733;
    wire N__58730;
    wire N__58727;
    wire N__58724;
    wire N__58721;
    wire N__58716;
    wire N__58707;
    wire N__58704;
    wire N__58701;
    wire N__58700;
    wire N__58697;
    wire N__58696;
    wire N__58693;
    wire N__58692;
    wire N__58691;
    wire N__58688;
    wire N__58685;
    wire N__58684;
    wire N__58681;
    wire N__58678;
    wire N__58675;
    wire N__58670;
    wire N__58667;
    wire N__58666;
    wire N__58661;
    wire N__58660;
    wire N__58657;
    wire N__58652;
    wire N__58649;
    wire N__58646;
    wire N__58643;
    wire N__58638;
    wire N__58635;
    wire N__58634;
    wire N__58629;
    wire N__58626;
    wire N__58623;
    wire N__58620;
    wire N__58617;
    wire N__58612;
    wire N__58609;
    wire N__58602;
    wire N__58599;
    wire N__58596;
    wire N__58595;
    wire N__58594;
    wire N__58593;
    wire N__58592;
    wire N__58591;
    wire N__58590;
    wire N__58589;
    wire N__58586;
    wire N__58583;
    wire N__58580;
    wire N__58577;
    wire N__58574;
    wire N__58571;
    wire N__58568;
    wire N__58565;
    wire N__58562;
    wire N__58561;
    wire N__58556;
    wire N__58553;
    wire N__58550;
    wire N__58545;
    wire N__58540;
    wire N__58537;
    wire N__58534;
    wire N__58531;
    wire N__58524;
    wire N__58521;
    wire N__58518;
    wire N__58515;
    wire N__58512;
    wire N__58509;
    wire N__58500;
    wire N__58499;
    wire N__58498;
    wire N__58497;
    wire N__58496;
    wire N__58493;
    wire N__58490;
    wire N__58489;
    wire N__58486;
    wire N__58483;
    wire N__58480;
    wire N__58477;
    wire N__58474;
    wire N__58473;
    wire N__58470;
    wire N__58465;
    wire N__58462;
    wire N__58459;
    wire N__58456;
    wire N__58455;
    wire N__58452;
    wire N__58449;
    wire N__58444;
    wire N__58441;
    wire N__58440;
    wire N__58437;
    wire N__58434;
    wire N__58431;
    wire N__58428;
    wire N__58425;
    wire N__58422;
    wire N__58419;
    wire N__58416;
    wire N__58413;
    wire N__58406;
    wire N__58403;
    wire N__58400;
    wire N__58395;
    wire N__58386;
    wire N__58383;
    wire N__58380;
    wire N__58377;
    wire N__58376;
    wire N__58373;
    wire N__58370;
    wire N__58365;
    wire N__58364;
    wire N__58361;
    wire N__58358;
    wire N__58357;
    wire N__58352;
    wire N__58351;
    wire N__58350;
    wire N__58349;
    wire N__58348;
    wire N__58345;
    wire N__58342;
    wire N__58339;
    wire N__58336;
    wire N__58333;
    wire N__58332;
    wire N__58329;
    wire N__58326;
    wire N__58323;
    wire N__58316;
    wire N__58313;
    wire N__58310;
    wire N__58307;
    wire N__58302;
    wire N__58299;
    wire N__58296;
    wire N__58293;
    wire N__58290;
    wire N__58287;
    wire N__58284;
    wire N__58281;
    wire N__58276;
    wire N__58269;
    wire N__58266;
    wire N__58263;
    wire N__58260;
    wire N__58257;
    wire N__58256;
    wire N__58253;
    wire N__58250;
    wire N__58247;
    wire N__58246;
    wire N__58243;
    wire N__58240;
    wire N__58237;
    wire N__58232;
    wire N__58227;
    wire N__58224;
    wire N__58223;
    wire N__58220;
    wire N__58217;
    wire N__58212;
    wire N__58211;
    wire N__58208;
    wire N__58205;
    wire N__58200;
    wire N__58199;
    wire N__58198;
    wire N__58197;
    wire N__58196;
    wire N__58191;
    wire N__58190;
    wire N__58187;
    wire N__58186;
    wire N__58185;
    wire N__58184;
    wire N__58183;
    wire N__58182;
    wire N__58181;
    wire N__58180;
    wire N__58179;
    wire N__58174;
    wire N__58171;
    wire N__58166;
    wire N__58165;
    wire N__58160;
    wire N__58159;
    wire N__58158;
    wire N__58157;
    wire N__58156;
    wire N__58153;
    wire N__58148;
    wire N__58143;
    wire N__58140;
    wire N__58135;
    wire N__58132;
    wire N__58129;
    wire N__58126;
    wire N__58121;
    wire N__58120;
    wire N__58117;
    wire N__58114;
    wire N__58113;
    wire N__58112;
    wire N__58111;
    wire N__58110;
    wire N__58105;
    wire N__58102;
    wire N__58099;
    wire N__58094;
    wire N__58089;
    wire N__58086;
    wire N__58083;
    wire N__58078;
    wire N__58073;
    wire N__58068;
    wire N__58065;
    wire N__58060;
    wire N__58057;
    wire N__58050;
    wire N__58045;
    wire N__58038;
    wire N__58035;
    wire N__58032;
    wire N__58027;
    wire N__58024;
    wire N__58017;
    wire N__58016;
    wire N__58015;
    wire N__58014;
    wire N__58013;
    wire N__58008;
    wire N__58007;
    wire N__58006;
    wire N__58005;
    wire N__58004;
    wire N__58001;
    wire N__57996;
    wire N__57993;
    wire N__57992;
    wire N__57991;
    wire N__57990;
    wire N__57989;
    wire N__57988;
    wire N__57987;
    wire N__57982;
    wire N__57981;
    wire N__57980;
    wire N__57979;
    wire N__57978;
    wire N__57973;
    wire N__57970;
    wire N__57967;
    wire N__57964;
    wire N__57959;
    wire N__57954;
    wire N__57949;
    wire N__57946;
    wire N__57943;
    wire N__57942;
    wire N__57941;
    wire N__57936;
    wire N__57935;
    wire N__57932;
    wire N__57927;
    wire N__57926;
    wire N__57923;
    wire N__57918;
    wire N__57915;
    wire N__57914;
    wire N__57911;
    wire N__57906;
    wire N__57901;
    wire N__57898;
    wire N__57895;
    wire N__57890;
    wire N__57887;
    wire N__57880;
    wire N__57877;
    wire N__57872;
    wire N__57869;
    wire N__57866;
    wire N__57861;
    wire N__57852;
    wire N__57849;
    wire N__57846;
    wire N__57841;
    wire N__57834;
    wire N__57833;
    wire N__57830;
    wire N__57827;
    wire N__57826;
    wire N__57823;
    wire N__57820;
    wire N__57817;
    wire N__57814;
    wire N__57811;
    wire N__57808;
    wire N__57801;
    wire N__57800;
    wire N__57799;
    wire N__57796;
    wire N__57793;
    wire N__57790;
    wire N__57787;
    wire N__57784;
    wire N__57781;
    wire N__57778;
    wire N__57775;
    wire N__57772;
    wire N__57769;
    wire N__57764;
    wire N__57761;
    wire N__57758;
    wire N__57753;
    wire N__57750;
    wire N__57747;
    wire N__57744;
    wire N__57743;
    wire N__57740;
    wire N__57737;
    wire N__57736;
    wire N__57731;
    wire N__57728;
    wire N__57723;
    wire N__57720;
    wire N__57719;
    wire N__57718;
    wire N__57715;
    wire N__57710;
    wire N__57705;
    wire N__57702;
    wire N__57699;
    wire N__57696;
    wire N__57693;
    wire N__57690;
    wire N__57687;
    wire N__57686;
    wire N__57685;
    wire N__57682;
    wire N__57679;
    wire N__57676;
    wire N__57671;
    wire N__57668;
    wire N__57665;
    wire N__57662;
    wire N__57659;
    wire N__57656;
    wire N__57653;
    wire N__57650;
    wire N__57645;
    wire N__57642;
    wire N__57639;
    wire N__57636;
    wire N__57633;
    wire N__57632;
    wire N__57629;
    wire N__57628;
    wire N__57627;
    wire N__57624;
    wire N__57621;
    wire N__57620;
    wire N__57619;
    wire N__57618;
    wire N__57615;
    wire N__57612;
    wire N__57609;
    wire N__57608;
    wire N__57605;
    wire N__57602;
    wire N__57601;
    wire N__57598;
    wire N__57595;
    wire N__57592;
    wire N__57589;
    wire N__57586;
    wire N__57583;
    wire N__57580;
    wire N__57577;
    wire N__57574;
    wire N__57571;
    wire N__57568;
    wire N__57561;
    wire N__57558;
    wire N__57555;
    wire N__57540;
    wire N__57537;
    wire N__57536;
    wire N__57535;
    wire N__57534;
    wire N__57531;
    wire N__57528;
    wire N__57525;
    wire N__57524;
    wire N__57521;
    wire N__57520;
    wire N__57513;
    wire N__57510;
    wire N__57509;
    wire N__57506;
    wire N__57503;
    wire N__57500;
    wire N__57497;
    wire N__57496;
    wire N__57493;
    wire N__57490;
    wire N__57487;
    wire N__57482;
    wire N__57479;
    wire N__57476;
    wire N__57475;
    wire N__57472;
    wire N__57469;
    wire N__57464;
    wire N__57461;
    wire N__57458;
    wire N__57453;
    wire N__57450;
    wire N__57447;
    wire N__57444;
    wire N__57435;
    wire N__57432;
    wire N__57429;
    wire N__57426;
    wire N__57423;
    wire N__57420;
    wire N__57419;
    wire N__57418;
    wire N__57415;
    wire N__57414;
    wire N__57413;
    wire N__57412;
    wire N__57409;
    wire N__57406;
    wire N__57403;
    wire N__57400;
    wire N__57397;
    wire N__57394;
    wire N__57393;
    wire N__57392;
    wire N__57389;
    wire N__57386;
    wire N__57383;
    wire N__57380;
    wire N__57375;
    wire N__57374;
    wire N__57371;
    wire N__57368;
    wire N__57361;
    wire N__57356;
    wire N__57353;
    wire N__57350;
    wire N__57343;
    wire N__57340;
    wire N__57337;
    wire N__57330;
    wire N__57327;
    wire N__57324;
    wire N__57323;
    wire N__57320;
    wire N__57319;
    wire N__57316;
    wire N__57313;
    wire N__57310;
    wire N__57307;
    wire N__57300;
    wire N__57297;
    wire N__57294;
    wire N__57291;
    wire N__57288;
    wire N__57287;
    wire N__57284;
    wire N__57281;
    wire N__57278;
    wire N__57275;
    wire N__57272;
    wire N__57267;
    wire N__57264;
    wire N__57261;
    wire N__57258;
    wire N__57255;
    wire N__57252;
    wire N__57249;
    wire N__57248;
    wire N__57243;
    wire N__57242;
    wire N__57239;
    wire N__57238;
    wire N__57237;
    wire N__57234;
    wire N__57231;
    wire N__57228;
    wire N__57227;
    wire N__57224;
    wire N__57223;
    wire N__57220;
    wire N__57217;
    wire N__57216;
    wire N__57213;
    wire N__57210;
    wire N__57209;
    wire N__57208;
    wire N__57205;
    wire N__57202;
    wire N__57197;
    wire N__57194;
    wire N__57191;
    wire N__57188;
    wire N__57185;
    wire N__57182;
    wire N__57179;
    wire N__57176;
    wire N__57173;
    wire N__57170;
    wire N__57167;
    wire N__57150;
    wire N__57147;
    wire N__57146;
    wire N__57143;
    wire N__57138;
    wire N__57135;
    wire N__57132;
    wire N__57131;
    wire N__57128;
    wire N__57125;
    wire N__57124;
    wire N__57123;
    wire N__57120;
    wire N__57117;
    wire N__57114;
    wire N__57111;
    wire N__57104;
    wire N__57101;
    wire N__57098;
    wire N__57093;
    wire N__57090;
    wire N__57089;
    wire N__57086;
    wire N__57083;
    wire N__57082;
    wire N__57079;
    wire N__57076;
    wire N__57073;
    wire N__57066;
    wire N__57063;
    wire N__57060;
    wire N__57057;
    wire N__57056;
    wire N__57053;
    wire N__57050;
    wire N__57047;
    wire N__57044;
    wire N__57041;
    wire N__57036;
    wire N__57033;
    wire N__57030;
    wire N__57029;
    wire N__57028;
    wire N__57023;
    wire N__57020;
    wire N__57015;
    wire N__57014;
    wire N__57013;
    wire N__57012;
    wire N__57009;
    wire N__57006;
    wire N__57003;
    wire N__57002;
    wire N__56999;
    wire N__56996;
    wire N__56995;
    wire N__56994;
    wire N__56993;
    wire N__56990;
    wire N__56985;
    wire N__56980;
    wire N__56973;
    wire N__56964;
    wire N__56961;
    wire N__56958;
    wire N__56955;
    wire N__56952;
    wire N__56949;
    wire N__56948;
    wire N__56947;
    wire N__56946;
    wire N__56943;
    wire N__56940;
    wire N__56935;
    wire N__56932;
    wire N__56929;
    wire N__56926;
    wire N__56921;
    wire N__56916;
    wire N__56915;
    wire N__56910;
    wire N__56909;
    wire N__56908;
    wire N__56905;
    wire N__56902;
    wire N__56899;
    wire N__56896;
    wire N__56889;
    wire N__56886;
    wire N__56885;
    wire N__56882;
    wire N__56879;
    wire N__56878;
    wire N__56873;
    wire N__56870;
    wire N__56869;
    wire N__56868;
    wire N__56863;
    wire N__56858;
    wire N__56853;
    wire N__56850;
    wire N__56847;
    wire N__56844;
    wire N__56843;
    wire N__56840;
    wire N__56837;
    wire N__56834;
    wire N__56829;
    wire N__56828;
    wire N__56825;
    wire N__56822;
    wire N__56819;
    wire N__56818;
    wire N__56817;
    wire N__56816;
    wire N__56815;
    wire N__56812;
    wire N__56809;
    wire N__56806;
    wire N__56799;
    wire N__56796;
    wire N__56787;
    wire N__56784;
    wire N__56781;
    wire N__56778;
    wire N__56775;
    wire N__56772;
    wire N__56771;
    wire N__56770;
    wire N__56767;
    wire N__56762;
    wire N__56757;
    wire N__56754;
    wire N__56751;
    wire N__56748;
    wire N__56745;
    wire N__56742;
    wire N__56739;
    wire N__56736;
    wire N__56733;
    wire N__56730;
    wire N__56729;
    wire N__56728;
    wire N__56727;
    wire N__56726;
    wire N__56725;
    wire N__56722;
    wire N__56719;
    wire N__56718;
    wire N__56713;
    wire N__56708;
    wire N__56705;
    wire N__56702;
    wire N__56701;
    wire N__56700;
    wire N__56697;
    wire N__56692;
    wire N__56687;
    wire N__56684;
    wire N__56681;
    wire N__56670;
    wire N__56667;
    wire N__56664;
    wire N__56661;
    wire N__56660;
    wire N__56657;
    wire N__56654;
    wire N__56651;
    wire N__56650;
    wire N__56649;
    wire N__56646;
    wire N__56643;
    wire N__56638;
    wire N__56631;
    wire N__56628;
    wire N__56627;
    wire N__56622;
    wire N__56621;
    wire N__56620;
    wire N__56617;
    wire N__56612;
    wire N__56607;
    wire N__56606;
    wire N__56601;
    wire N__56598;
    wire N__56595;
    wire N__56594;
    wire N__56593;
    wire N__56592;
    wire N__56591;
    wire N__56588;
    wire N__56585;
    wire N__56584;
    wire N__56583;
    wire N__56578;
    wire N__56575;
    wire N__56574;
    wire N__56569;
    wire N__56564;
    wire N__56561;
    wire N__56560;
    wire N__56559;
    wire N__56554;
    wire N__56549;
    wire N__56546;
    wire N__56543;
    wire N__56540;
    wire N__56537;
    wire N__56534;
    wire N__56529;
    wire N__56520;
    wire N__56517;
    wire N__56516;
    wire N__56513;
    wire N__56512;
    wire N__56511;
    wire N__56508;
    wire N__56505;
    wire N__56500;
    wire N__56493;
    wire N__56490;
    wire N__56489;
    wire N__56486;
    wire N__56483;
    wire N__56480;
    wire N__56477;
    wire N__56472;
    wire N__56469;
    wire N__56468;
    wire N__56465;
    wire N__56462;
    wire N__56459;
    wire N__56456;
    wire N__56453;
    wire N__56448;
    wire N__56447;
    wire N__56446;
    wire N__56443;
    wire N__56442;
    wire N__56441;
    wire N__56440;
    wire N__56439;
    wire N__56434;
    wire N__56431;
    wire N__56428;
    wire N__56425;
    wire N__56422;
    wire N__56419;
    wire N__56416;
    wire N__56411;
    wire N__56408;
    wire N__56407;
    wire N__56406;
    wire N__56403;
    wire N__56394;
    wire N__56389;
    wire N__56384;
    wire N__56379;
    wire N__56376;
    wire N__56373;
    wire N__56370;
    wire N__56367;
    wire N__56364;
    wire N__56361;
    wire N__56360;
    wire N__56359;
    wire N__56358;
    wire N__56357;
    wire N__56354;
    wire N__56353;
    wire N__56352;
    wire N__56351;
    wire N__56350;
    wire N__56347;
    wire N__56340;
    wire N__56337;
    wire N__56336;
    wire N__56333;
    wire N__56330;
    wire N__56327;
    wire N__56324;
    wire N__56317;
    wire N__56312;
    wire N__56309;
    wire N__56308;
    wire N__56299;
    wire N__56296;
    wire N__56293;
    wire N__56290;
    wire N__56283;
    wire N__56280;
    wire N__56277;
    wire N__56274;
    wire N__56271;
    wire N__56268;
    wire N__56265;
    wire N__56262;
    wire N__56259;
    wire N__56256;
    wire N__56253;
    wire N__56250;
    wire N__56249;
    wire N__56248;
    wire N__56247;
    wire N__56246;
    wire N__56245;
    wire N__56242;
    wire N__56239;
    wire N__56236;
    wire N__56233;
    wire N__56232;
    wire N__56229;
    wire N__56226;
    wire N__56223;
    wire N__56216;
    wire N__56213;
    wire N__56210;
    wire N__56207;
    wire N__56204;
    wire N__56201;
    wire N__56198;
    wire N__56195;
    wire N__56186;
    wire N__56181;
    wire N__56180;
    wire N__56177;
    wire N__56174;
    wire N__56173;
    wire N__56170;
    wire N__56167;
    wire N__56164;
    wire N__56159;
    wire N__56154;
    wire N__56151;
    wire N__56148;
    wire N__56147;
    wire N__56146;
    wire N__56145;
    wire N__56144;
    wire N__56141;
    wire N__56138;
    wire N__56131;
    wire N__56130;
    wire N__56129;
    wire N__56128;
    wire N__56127;
    wire N__56124;
    wire N__56123;
    wire N__56122;
    wire N__56119;
    wire N__56116;
    wire N__56113;
    wire N__56110;
    wire N__56105;
    wire N__56102;
    wire N__56099;
    wire N__56096;
    wire N__56093;
    wire N__56088;
    wire N__56081;
    wire N__56070;
    wire N__56069;
    wire N__56066;
    wire N__56063;
    wire N__56058;
    wire N__56057;
    wire N__56056;
    wire N__56053;
    wire N__56050;
    wire N__56047;
    wire N__56040;
    wire N__56037;
    wire N__56036;
    wire N__56031;
    wire N__56028;
    wire N__56027;
    wire N__56022;
    wire N__56019;
    wire N__56016;
    wire N__56013;
    wire N__56010;
    wire N__56007;
    wire N__56004;
    wire N__56001;
    wire N__55998;
    wire N__55995;
    wire N__55992;
    wire N__55989;
    wire N__55988;
    wire N__55983;
    wire N__55982;
    wire N__55979;
    wire N__55976;
    wire N__55971;
    wire N__55968;
    wire N__55965;
    wire N__55964;
    wire N__55961;
    wire N__55960;
    wire N__55957;
    wire N__55954;
    wire N__55951;
    wire N__55944;
    wire N__55943;
    wire N__55940;
    wire N__55937;
    wire N__55934;
    wire N__55929;
    wire N__55928;
    wire N__55927;
    wire N__55924;
    wire N__55921;
    wire N__55920;
    wire N__55917;
    wire N__55916;
    wire N__55913;
    wire N__55910;
    wire N__55907;
    wire N__55904;
    wire N__55901;
    wire N__55896;
    wire N__55893;
    wire N__55890;
    wire N__55887;
    wire N__55884;
    wire N__55875;
    wire N__55872;
    wire N__55869;
    wire N__55868;
    wire N__55865;
    wire N__55864;
    wire N__55863;
    wire N__55862;
    wire N__55861;
    wire N__55858;
    wire N__55857;
    wire N__55856;
    wire N__55855;
    wire N__55854;
    wire N__55853;
    wire N__55850;
    wire N__55847;
    wire N__55844;
    wire N__55841;
    wire N__55838;
    wire N__55835;
    wire N__55824;
    wire N__55817;
    wire N__55808;
    wire N__55805;
    wire N__55800;
    wire N__55797;
    wire N__55796;
    wire N__55795;
    wire N__55794;
    wire N__55791;
    wire N__55788;
    wire N__55785;
    wire N__55782;
    wire N__55775;
    wire N__55770;
    wire N__55767;
    wire N__55764;
    wire N__55761;
    wire N__55758;
    wire N__55755;
    wire N__55752;
    wire N__55749;
    wire N__55746;
    wire N__55745;
    wire N__55744;
    wire N__55743;
    wire N__55742;
    wire N__55741;
    wire N__55740;
    wire N__55735;
    wire N__55728;
    wire N__55727;
    wire N__55726;
    wire N__55725;
    wire N__55724;
    wire N__55723;
    wire N__55722;
    wire N__55717;
    wire N__55712;
    wire N__55707;
    wire N__55702;
    wire N__55697;
    wire N__55696;
    wire N__55695;
    wire N__55694;
    wire N__55693;
    wire N__55690;
    wire N__55689;
    wire N__55688;
    wire N__55687;
    wire N__55686;
    wire N__55683;
    wire N__55680;
    wire N__55675;
    wire N__55670;
    wire N__55665;
    wire N__55662;
    wire N__55653;
    wire N__55652;
    wire N__55651;
    wire N__55650;
    wire N__55645;
    wire N__55640;
    wire N__55637;
    wire N__55632;
    wire N__55625;
    wire N__55622;
    wire N__55619;
    wire N__55612;
    wire N__55609;
    wire N__55606;
    wire N__55603;
    wire N__55596;
    wire N__55593;
    wire N__55590;
    wire N__55587;
    wire N__55584;
    wire N__55581;
    wire N__55578;
    wire N__55575;
    wire N__55572;
    wire N__55571;
    wire N__55570;
    wire N__55567;
    wire N__55564;
    wire N__55563;
    wire N__55560;
    wire N__55559;
    wire N__55558;
    wire N__55555;
    wire N__55552;
    wire N__55549;
    wire N__55546;
    wire N__55543;
    wire N__55540;
    wire N__55539;
    wire N__55538;
    wire N__55531;
    wire N__55526;
    wire N__55523;
    wire N__55522;
    wire N__55521;
    wire N__55518;
    wire N__55515;
    wire N__55512;
    wire N__55507;
    wire N__55504;
    wire N__55501;
    wire N__55498;
    wire N__55495;
    wire N__55492;
    wire N__55489;
    wire N__55484;
    wire N__55481;
    wire N__55478;
    wire N__55475;
    wire N__55472;
    wire N__55467;
    wire N__55460;
    wire N__55455;
    wire N__55454;
    wire N__55453;
    wire N__55452;
    wire N__55451;
    wire N__55450;
    wire N__55449;
    wire N__55448;
    wire N__55447;
    wire N__55446;
    wire N__55445;
    wire N__55444;
    wire N__55439;
    wire N__55438;
    wire N__55435;
    wire N__55432;
    wire N__55431;
    wire N__55430;
    wire N__55429;
    wire N__55428;
    wire N__55427;
    wire N__55424;
    wire N__55423;
    wire N__55420;
    wire N__55417;
    wire N__55410;
    wire N__55409;
    wire N__55406;
    wire N__55403;
    wire N__55400;
    wire N__55399;
    wire N__55396;
    wire N__55391;
    wire N__55388;
    wire N__55387;
    wire N__55386;
    wire N__55383;
    wire N__55376;
    wire N__55373;
    wire N__55370;
    wire N__55367;
    wire N__55362;
    wire N__55359;
    wire N__55352;
    wire N__55351;
    wire N__55348;
    wire N__55345;
    wire N__55342;
    wire N__55339;
    wire N__55336;
    wire N__55333;
    wire N__55328;
    wire N__55319;
    wire N__55314;
    wire N__55311;
    wire N__55306;
    wire N__55303;
    wire N__55296;
    wire N__55291;
    wire N__55288;
    wire N__55283;
    wire N__55278;
    wire N__55275;
    wire N__55272;
    wire N__55263;
    wire N__55262;
    wire N__55259;
    wire N__55258;
    wire N__55257;
    wire N__55256;
    wire N__55255;
    wire N__55254;
    wire N__55251;
    wire N__55250;
    wire N__55249;
    wire N__55246;
    wire N__55239;
    wire N__55236;
    wire N__55233;
    wire N__55232;
    wire N__55231;
    wire N__55230;
    wire N__55229;
    wire N__55228;
    wire N__55225;
    wire N__55222;
    wire N__55221;
    wire N__55218;
    wire N__55217;
    wire N__55212;
    wire N__55209;
    wire N__55206;
    wire N__55199;
    wire N__55198;
    wire N__55193;
    wire N__55192;
    wire N__55187;
    wire N__55184;
    wire N__55183;
    wire N__55180;
    wire N__55177;
    wire N__55174;
    wire N__55167;
    wire N__55164;
    wire N__55163;
    wire N__55160;
    wire N__55157;
    wire N__55156;
    wire N__55155;
    wire N__55154;
    wire N__55151;
    wire N__55148;
    wire N__55145;
    wire N__55140;
    wire N__55135;
    wire N__55132;
    wire N__55129;
    wire N__55126;
    wire N__55123;
    wire N__55120;
    wire N__55117;
    wire N__55114;
    wire N__55113;
    wire N__55110;
    wire N__55105;
    wire N__55098;
    wire N__55085;
    wire N__55082;
    wire N__55079;
    wire N__55076;
    wire N__55069;
    wire N__55062;
    wire N__55059;
    wire N__55058;
    wire N__55057;
    wire N__55056;
    wire N__55055;
    wire N__55054;
    wire N__55053;
    wire N__55052;
    wire N__55049;
    wire N__55046;
    wire N__55043;
    wire N__55040;
    wire N__55037;
    wire N__55036;
    wire N__55035;
    wire N__55032;
    wire N__55031;
    wire N__55030;
    wire N__55029;
    wire N__55026;
    wire N__55023;
    wire N__55022;
    wire N__55021;
    wire N__55020;
    wire N__55019;
    wire N__55014;
    wire N__55011;
    wire N__55010;
    wire N__55005;
    wire N__55002;
    wire N__55001;
    wire N__54998;
    wire N__54995;
    wire N__54992;
    wire N__54989;
    wire N__54986;
    wire N__54979;
    wire N__54976;
    wire N__54973;
    wire N__54970;
    wire N__54967;
    wire N__54964;
    wire N__54963;
    wire N__54960;
    wire N__54955;
    wire N__54954;
    wire N__54953;
    wire N__54950;
    wire N__54947;
    wire N__54944;
    wire N__54939;
    wire N__54930;
    wire N__54929;
    wire N__54928;
    wire N__54925;
    wire N__54920;
    wire N__54917;
    wire N__54914;
    wire N__54911;
    wire N__54908;
    wire N__54905;
    wire N__54902;
    wire N__54893;
    wire N__54888;
    wire N__54885;
    wire N__54882;
    wire N__54879;
    wire N__54874;
    wire N__54871;
    wire N__54862;
    wire N__54859;
    wire N__54854;
    wire N__54851;
    wire N__54846;
    wire N__54837;
    wire N__54836;
    wire N__54835;
    wire N__54834;
    wire N__54833;
    wire N__54832;
    wire N__54829;
    wire N__54826;
    wire N__54825;
    wire N__54822;
    wire N__54821;
    wire N__54820;
    wire N__54819;
    wire N__54818;
    wire N__54817;
    wire N__54816;
    wire N__54813;
    wire N__54810;
    wire N__54807;
    wire N__54806;
    wire N__54803;
    wire N__54802;
    wire N__54799;
    wire N__54798;
    wire N__54795;
    wire N__54792;
    wire N__54789;
    wire N__54784;
    wire N__54783;
    wire N__54782;
    wire N__54781;
    wire N__54780;
    wire N__54775;
    wire N__54772;
    wire N__54769;
    wire N__54764;
    wire N__54761;
    wire N__54758;
    wire N__54757;
    wire N__54756;
    wire N__54753;
    wire N__54750;
    wire N__54747;
    wire N__54744;
    wire N__54737;
    wire N__54736;
    wire N__54735;
    wire N__54732;
    wire N__54729;
    wire N__54724;
    wire N__54721;
    wire N__54712;
    wire N__54709;
    wire N__54706;
    wire N__54703;
    wire N__54698;
    wire N__54691;
    wire N__54686;
    wire N__54675;
    wire N__54672;
    wire N__54669;
    wire N__54660;
    wire N__54657;
    wire N__54654;
    wire N__54649;
    wire N__54646;
    wire N__54639;
    wire N__54638;
    wire N__54635;
    wire N__54634;
    wire N__54631;
    wire N__54628;
    wire N__54623;
    wire N__54620;
    wire N__54617;
    wire N__54614;
    wire N__54611;
    wire N__54606;
    wire N__54603;
    wire N__54600;
    wire N__54599;
    wire N__54598;
    wire N__54595;
    wire N__54592;
    wire N__54589;
    wire N__54586;
    wire N__54581;
    wire N__54576;
    wire N__54573;
    wire N__54570;
    wire N__54567;
    wire N__54564;
    wire N__54561;
    wire N__54558;
    wire N__54555;
    wire N__54552;
    wire N__54549;
    wire N__54546;
    wire N__54543;
    wire N__54540;
    wire N__54537;
    wire N__54534;
    wire N__54531;
    wire N__54528;
    wire N__54525;
    wire N__54524;
    wire N__54523;
    wire N__54522;
    wire N__54521;
    wire N__54520;
    wire N__54519;
    wire N__54518;
    wire N__54517;
    wire N__54516;
    wire N__54515;
    wire N__54514;
    wire N__54513;
    wire N__54512;
    wire N__54511;
    wire N__54510;
    wire N__54509;
    wire N__54508;
    wire N__54507;
    wire N__54506;
    wire N__54505;
    wire N__54504;
    wire N__54503;
    wire N__54502;
    wire N__54501;
    wire N__54500;
    wire N__54499;
    wire N__54498;
    wire N__54497;
    wire N__54496;
    wire N__54495;
    wire N__54494;
    wire N__54429;
    wire N__54426;
    wire N__54423;
    wire N__54420;
    wire N__54419;
    wire N__54416;
    wire N__54413;
    wire N__54410;
    wire N__54405;
    wire N__54404;
    wire N__54403;
    wire N__54402;
    wire N__54399;
    wire N__54398;
    wire N__54395;
    wire N__54392;
    wire N__54389;
    wire N__54384;
    wire N__54381;
    wire N__54380;
    wire N__54373;
    wire N__54370;
    wire N__54367;
    wire N__54364;
    wire N__54359;
    wire N__54356;
    wire N__54351;
    wire N__54348;
    wire N__54345;
    wire N__54344;
    wire N__54343;
    wire N__54342;
    wire N__54339;
    wire N__54338;
    wire N__54337;
    wire N__54336;
    wire N__54335;
    wire N__54334;
    wire N__54331;
    wire N__54326;
    wire N__54323;
    wire N__54320;
    wire N__54315;
    wire N__54312;
    wire N__54309;
    wire N__54306;
    wire N__54303;
    wire N__54300;
    wire N__54293;
    wire N__54290;
    wire N__54289;
    wire N__54288;
    wire N__54285;
    wire N__54282;
    wire N__54277;
    wire N__54274;
    wire N__54269;
    wire N__54258;
    wire N__54255;
    wire N__54252;
    wire N__54251;
    wire N__54248;
    wire N__54245;
    wire N__54240;
    wire N__54237;
    wire N__54234;
    wire N__54231;
    wire N__54228;
    wire N__54225;
    wire N__54222;
    wire N__54219;
    wire N__54216;
    wire N__54213;
    wire N__54210;
    wire N__54207;
    wire N__54206;
    wire N__54203;
    wire N__54200;
    wire N__54197;
    wire N__54194;
    wire N__54193;
    wire N__54190;
    wire N__54187;
    wire N__54184;
    wire N__54177;
    wire N__54174;
    wire N__54171;
    wire N__54168;
    wire N__54165;
    wire N__54162;
    wire N__54159;
    wire N__54156;
    wire N__54153;
    wire N__54152;
    wire N__54149;
    wire N__54146;
    wire N__54143;
    wire N__54142;
    wire N__54139;
    wire N__54136;
    wire N__54133;
    wire N__54130;
    wire N__54123;
    wire N__54120;
    wire N__54119;
    wire N__54118;
    wire N__54115;
    wire N__54114;
    wire N__54113;
    wire N__54112;
    wire N__54109;
    wire N__54106;
    wire N__54103;
    wire N__54100;
    wire N__54097;
    wire N__54094;
    wire N__54091;
    wire N__54086;
    wire N__54083;
    wire N__54080;
    wire N__54077;
    wire N__54074;
    wire N__54071;
    wire N__54068;
    wire N__54065;
    wire N__54060;
    wire N__54057;
    wire N__54048;
    wire N__54045;
    wire N__54042;
    wire N__54039;
    wire N__54036;
    wire N__54033;
    wire N__54030;
    wire N__54027;
    wire N__54024;
    wire N__54021;
    wire N__54018;
    wire N__54015;
    wire N__54012;
    wire N__54009;
    wire N__54006;
    wire N__54005;
    wire N__54004;
    wire N__54003;
    wire N__54002;
    wire N__54001;
    wire N__53998;
    wire N__53995;
    wire N__53994;
    wire N__53993;
    wire N__53992;
    wire N__53991;
    wire N__53988;
    wire N__53985;
    wire N__53980;
    wire N__53979;
    wire N__53978;
    wire N__53977;
    wire N__53976;
    wire N__53973;
    wire N__53970;
    wire N__53969;
    wire N__53968;
    wire N__53967;
    wire N__53966;
    wire N__53963;
    wire N__53962;
    wire N__53961;
    wire N__53960;
    wire N__53959;
    wire N__53956;
    wire N__53953;
    wire N__53950;
    wire N__53949;
    wire N__53948;
    wire N__53945;
    wire N__53942;
    wire N__53939;
    wire N__53934;
    wire N__53931;
    wire N__53928;
    wire N__53925;
    wire N__53922;
    wire N__53919;
    wire N__53914;
    wire N__53911;
    wire N__53908;
    wire N__53905;
    wire N__53902;
    wire N__53899;
    wire N__53896;
    wire N__53893;
    wire N__53888;
    wire N__53885;
    wire N__53882;
    wire N__53879;
    wire N__53874;
    wire N__53871;
    wire N__53868;
    wire N__53865;
    wire N__53858;
    wire N__53853;
    wire N__53832;
    wire N__53827;
    wire N__53824;
    wire N__53819;
    wire N__53816;
    wire N__53813;
    wire N__53810;
    wire N__53805;
    wire N__53802;
    wire N__53793;
    wire N__53792;
    wire N__53789;
    wire N__53788;
    wire N__53785;
    wire N__53782;
    wire N__53779;
    wire N__53776;
    wire N__53773;
    wire N__53770;
    wire N__53767;
    wire N__53764;
    wire N__53761;
    wire N__53756;
    wire N__53753;
    wire N__53750;
    wire N__53745;
    wire N__53742;
    wire N__53739;
    wire N__53736;
    wire N__53733;
    wire N__53730;
    wire N__53727;
    wire N__53724;
    wire N__53721;
    wire N__53720;
    wire N__53719;
    wire N__53718;
    wire N__53717;
    wire N__53716;
    wire N__53715;
    wire N__53714;
    wire N__53713;
    wire N__53712;
    wire N__53709;
    wire N__53704;
    wire N__53701;
    wire N__53696;
    wire N__53695;
    wire N__53694;
    wire N__53693;
    wire N__53692;
    wire N__53691;
    wire N__53690;
    wire N__53689;
    wire N__53684;
    wire N__53679;
    wire N__53676;
    wire N__53675;
    wire N__53674;
    wire N__53673;
    wire N__53672;
    wire N__53671;
    wire N__53670;
    wire N__53669;
    wire N__53666;
    wire N__53661;
    wire N__53656;
    wire N__53651;
    wire N__53648;
    wire N__53643;
    wire N__53640;
    wire N__53637;
    wire N__53634;
    wire N__53629;
    wire N__53626;
    wire N__53623;
    wire N__53620;
    wire N__53615;
    wire N__53610;
    wire N__53607;
    wire N__53596;
    wire N__53593;
    wire N__53588;
    wire N__53585;
    wire N__53578;
    wire N__53573;
    wire N__53568;
    wire N__53565;
    wire N__53562;
    wire N__53559;
    wire N__53556;
    wire N__53547;
    wire N__53544;
    wire N__53541;
    wire N__53538;
    wire N__53535;
    wire N__53532;
    wire N__53529;
    wire N__53526;
    wire N__53525;
    wire N__53524;
    wire N__53521;
    wire N__53518;
    wire N__53515;
    wire N__53512;
    wire N__53509;
    wire N__53504;
    wire N__53501;
    wire N__53496;
    wire N__53493;
    wire N__53490;
    wire N__53487;
    wire N__53484;
    wire N__53481;
    wire N__53478;
    wire N__53475;
    wire N__53472;
    wire N__53469;
    wire N__53466;
    wire N__53463;
    wire N__53460;
    wire N__53457;
    wire N__53454;
    wire N__53451;
    wire N__53448;
    wire N__53445;
    wire N__53442;
    wire N__53439;
    wire N__53436;
    wire N__53433;
    wire N__53430;
    wire N__53427;
    wire N__53424;
    wire N__53421;
    wire N__53420;
    wire N__53419;
    wire N__53416;
    wire N__53413;
    wire N__53410;
    wire N__53407;
    wire N__53404;
    wire N__53401;
    wire N__53398;
    wire N__53393;
    wire N__53390;
    wire N__53387;
    wire N__53382;
    wire N__53379;
    wire N__53376;
    wire N__53375;
    wire N__53372;
    wire N__53371;
    wire N__53368;
    wire N__53365;
    wire N__53362;
    wire N__53359;
    wire N__53356;
    wire N__53351;
    wire N__53348;
    wire N__53345;
    wire N__53340;
    wire N__53337;
    wire N__53334;
    wire N__53331;
    wire N__53330;
    wire N__53329;
    wire N__53328;
    wire N__53325;
    wire N__53324;
    wire N__53323;
    wire N__53320;
    wire N__53319;
    wire N__53318;
    wire N__53317;
    wire N__53316;
    wire N__53315;
    wire N__53314;
    wire N__53311;
    wire N__53310;
    wire N__53307;
    wire N__53306;
    wire N__53303;
    wire N__53300;
    wire N__53297;
    wire N__53296;
    wire N__53293;
    wire N__53290;
    wire N__53287;
    wire N__53286;
    wire N__53283;
    wire N__53282;
    wire N__53281;
    wire N__53278;
    wire N__53275;
    wire N__53272;
    wire N__53271;
    wire N__53270;
    wire N__53267;
    wire N__53266;
    wire N__53263;
    wire N__53262;
    wire N__53259;
    wire N__53258;
    wire N__53257;
    wire N__53256;
    wire N__53253;
    wire N__53250;
    wire N__53247;
    wire N__53244;
    wire N__53241;
    wire N__53238;
    wire N__53235;
    wire N__53232;
    wire N__53229;
    wire N__53226;
    wire N__53223;
    wire N__53220;
    wire N__53217;
    wire N__53214;
    wire N__53211;
    wire N__53208;
    wire N__53205;
    wire N__53202;
    wire N__53199;
    wire N__53196;
    wire N__53195;
    wire N__53194;
    wire N__53191;
    wire N__53188;
    wire N__53185;
    wire N__53182;
    wire N__53181;
    wire N__53180;
    wire N__53179;
    wire N__53176;
    wire N__53175;
    wire N__53172;
    wire N__53167;
    wire N__53162;
    wire N__53157;
    wire N__53154;
    wire N__53147;
    wire N__53142;
    wire N__53137;
    wire N__53130;
    wire N__53127;
    wire N__53124;
    wire N__53119;
    wire N__53116;
    wire N__53111;
    wire N__53108;
    wire N__53097;
    wire N__53090;
    wire N__53087;
    wire N__53082;
    wire N__53075;
    wire N__53068;
    wire N__53059;
    wire N__53056;
    wire N__53053;
    wire N__53048;
    wire N__53043;
    wire N__53034;
    wire N__53031;
    wire N__53028;
    wire N__53025;
    wire N__53022;
    wire N__53019;
    wire N__53016;
    wire N__53015;
    wire N__53014;
    wire N__53013;
    wire N__53012;
    wire N__53011;
    wire N__53010;
    wire N__53009;
    wire N__53008;
    wire N__53005;
    wire N__53004;
    wire N__53001;
    wire N__53000;
    wire N__52999;
    wire N__52998;
    wire N__52995;
    wire N__52994;
    wire N__52991;
    wire N__52990;
    wire N__52989;
    wire N__52988;
    wire N__52987;
    wire N__52984;
    wire N__52983;
    wire N__52982;
    wire N__52979;
    wire N__52976;
    wire N__52973;
    wire N__52970;
    wire N__52967;
    wire N__52964;
    wire N__52961;
    wire N__52958;
    wire N__52955;
    wire N__52952;
    wire N__52949;
    wire N__52946;
    wire N__52943;
    wire N__52940;
    wire N__52937;
    wire N__52934;
    wire N__52931;
    wire N__52928;
    wire N__52927;
    wire N__52926;
    wire N__52925;
    wire N__52924;
    wire N__52923;
    wire N__52922;
    wire N__52919;
    wire N__52916;
    wire N__52911;
    wire N__52908;
    wire N__52905;
    wire N__52904;
    wire N__52903;
    wire N__52902;
    wire N__52901;
    wire N__52894;
    wire N__52885;
    wire N__52882;
    wire N__52877;
    wire N__52872;
    wire N__52867;
    wire N__52854;
    wire N__52847;
    wire N__52842;
    wire N__52833;
    wire N__52830;
    wire N__52827;
    wire N__52816;
    wire N__52803;
    wire N__52800;
    wire N__52797;
    wire N__52794;
    wire N__52791;
    wire N__52788;
    wire N__52785;
    wire N__52782;
    wire N__52781;
    wire N__52780;
    wire N__52779;
    wire N__52776;
    wire N__52773;
    wire N__52772;
    wire N__52771;
    wire N__52770;
    wire N__52769;
    wire N__52768;
    wire N__52765;
    wire N__52762;
    wire N__52761;
    wire N__52760;
    wire N__52757;
    wire N__52756;
    wire N__52755;
    wire N__52752;
    wire N__52749;
    wire N__52746;
    wire N__52745;
    wire N__52744;
    wire N__52743;
    wire N__52742;
    wire N__52741;
    wire N__52740;
    wire N__52739;
    wire N__52738;
    wire N__52737;
    wire N__52736;
    wire N__52733;
    wire N__52730;
    wire N__52727;
    wire N__52722;
    wire N__52719;
    wire N__52716;
    wire N__52713;
    wire N__52710;
    wire N__52707;
    wire N__52702;
    wire N__52701;
    wire N__52700;
    wire N__52697;
    wire N__52694;
    wire N__52691;
    wire N__52688;
    wire N__52685;
    wire N__52682;
    wire N__52677;
    wire N__52676;
    wire N__52675;
    wire N__52674;
    wire N__52673;
    wire N__52672;
    wire N__52669;
    wire N__52666;
    wire N__52663;
    wire N__52660;
    wire N__52657;
    wire N__52648;
    wire N__52643;
    wire N__52640;
    wire N__52637;
    wire N__52634;
    wire N__52631;
    wire N__52626;
    wire N__52621;
    wire N__52614;
    wire N__52611;
    wire N__52608;
    wire N__52605;
    wire N__52602;
    wire N__52599;
    wire N__52592;
    wire N__52585;
    wire N__52578;
    wire N__52567;
    wire N__52548;
    wire N__52545;
    wire N__52542;
    wire N__52539;
    wire N__52536;
    wire N__52533;
    wire N__52530;
    wire N__52527;
    wire N__52526;
    wire N__52525;
    wire N__52524;
    wire N__52523;
    wire N__52522;
    wire N__52521;
    wire N__52520;
    wire N__52517;
    wire N__52514;
    wire N__52513;
    wire N__52512;
    wire N__52509;
    wire N__52506;
    wire N__52503;
    wire N__52500;
    wire N__52497;
    wire N__52496;
    wire N__52495;
    wire N__52494;
    wire N__52493;
    wire N__52492;
    wire N__52489;
    wire N__52488;
    wire N__52487;
    wire N__52486;
    wire N__52485;
    wire N__52484;
    wire N__52481;
    wire N__52478;
    wire N__52475;
    wire N__52472;
    wire N__52471;
    wire N__52468;
    wire N__52463;
    wire N__52458;
    wire N__52455;
    wire N__52450;
    wire N__52447;
    wire N__52446;
    wire N__52445;
    wire N__52442;
    wire N__52441;
    wire N__52440;
    wire N__52439;
    wire N__52438;
    wire N__52437;
    wire N__52434;
    wire N__52431;
    wire N__52428;
    wire N__52425;
    wire N__52422;
    wire N__52419;
    wire N__52410;
    wire N__52407;
    wire N__52404;
    wire N__52399;
    wire N__52396;
    wire N__52391;
    wire N__52388;
    wire N__52385;
    wire N__52382;
    wire N__52381;
    wire N__52378;
    wire N__52375;
    wire N__52372;
    wire N__52371;
    wire N__52370;
    wire N__52367;
    wire N__52364;
    wire N__52357;
    wire N__52354;
    wire N__52349;
    wire N__52344;
    wire N__52333;
    wire N__52330;
    wire N__52327;
    wire N__52324;
    wire N__52319;
    wire N__52316;
    wire N__52311;
    wire N__52308;
    wire N__52303;
    wire N__52298;
    wire N__52293;
    wire N__52284;
    wire N__52279;
    wire N__52276;
    wire N__52271;
    wire N__52268;
    wire N__52263;
    wire N__52254;
    wire N__52251;
    wire N__52248;
    wire N__52245;
    wire N__52242;
    wire N__52239;
    wire N__52236;
    wire N__52235;
    wire N__52234;
    wire N__52233;
    wire N__52232;
    wire N__52231;
    wire N__52228;
    wire N__52227;
    wire N__52224;
    wire N__52223;
    wire N__52222;
    wire N__52221;
    wire N__52220;
    wire N__52217;
    wire N__52216;
    wire N__52215;
    wire N__52214;
    wire N__52213;
    wire N__52210;
    wire N__52207;
    wire N__52206;
    wire N__52205;
    wire N__52204;
    wire N__52203;
    wire N__52200;
    wire N__52199;
    wire N__52198;
    wire N__52195;
    wire N__52192;
    wire N__52191;
    wire N__52188;
    wire N__52187;
    wire N__52186;
    wire N__52183;
    wire N__52182;
    wire N__52179;
    wire N__52176;
    wire N__52173;
    wire N__52170;
    wire N__52167;
    wire N__52164;
    wire N__52161;
    wire N__52158;
    wire N__52153;
    wire N__52150;
    wire N__52147;
    wire N__52146;
    wire N__52145;
    wire N__52142;
    wire N__52139;
    wire N__52136;
    wire N__52133;
    wire N__52130;
    wire N__52125;
    wire N__52124;
    wire N__52123;
    wire N__52122;
    wire N__52119;
    wire N__52116;
    wire N__52113;
    wire N__52110;
    wire N__52107;
    wire N__52104;
    wire N__52099;
    wire N__52090;
    wire N__52087;
    wire N__52080;
    wire N__52077;
    wire N__52074;
    wire N__52071;
    wire N__52066;
    wire N__52061;
    wire N__52058;
    wire N__52055;
    wire N__52054;
    wire N__52051;
    wire N__52048;
    wire N__52045;
    wire N__52038;
    wire N__52027;
    wire N__52020;
    wire N__52017;
    wire N__52006;
    wire N__52003;
    wire N__51984;
    wire N__51981;
    wire N__51978;
    wire N__51975;
    wire N__51972;
    wire N__51969;
    wire N__51966;
    wire N__51963;
    wire N__51960;
    wire N__51957;
    wire N__51954;
    wire N__51951;
    wire N__51950;
    wire N__51947;
    wire N__51946;
    wire N__51943;
    wire N__51940;
    wire N__51937;
    wire N__51936;
    wire N__51931;
    wire N__51928;
    wire N__51927;
    wire N__51926;
    wire N__51925;
    wire N__51924;
    wire N__51923;
    wire N__51922;
    wire N__51921;
    wire N__51920;
    wire N__51919;
    wire N__51916;
    wire N__51915;
    wire N__51910;
    wire N__51907;
    wire N__51906;
    wire N__51905;
    wire N__51904;
    wire N__51903;
    wire N__51902;
    wire N__51899;
    wire N__51896;
    wire N__51893;
    wire N__51892;
    wire N__51891;
    wire N__51890;
    wire N__51887;
    wire N__51884;
    wire N__51881;
    wire N__51878;
    wire N__51875;
    wire N__51872;
    wire N__51871;
    wire N__51868;
    wire N__51867;
    wire N__51866;
    wire N__51861;
    wire N__51860;
    wire N__51859;
    wire N__51856;
    wire N__51853;
    wire N__51850;
    wire N__51847;
    wire N__51846;
    wire N__51843;
    wire N__51840;
    wire N__51837;
    wire N__51834;
    wire N__51831;
    wire N__51828;
    wire N__51825;
    wire N__51824;
    wire N__51821;
    wire N__51814;
    wire N__51809;
    wire N__51804;
    wire N__51801;
    wire N__51798;
    wire N__51795;
    wire N__51792;
    wire N__51791;
    wire N__51790;
    wire N__51787;
    wire N__51784;
    wire N__51781;
    wire N__51776;
    wire N__51773;
    wire N__51770;
    wire N__51765;
    wire N__51760;
    wire N__51755;
    wire N__51752;
    wire N__51743;
    wire N__51740;
    wire N__51733;
    wire N__51730;
    wire N__51727;
    wire N__51718;
    wire N__51707;
    wire N__51702;
    wire N__51697;
    wire N__51684;
    wire N__51681;
    wire N__51678;
    wire N__51675;
    wire N__51672;
    wire N__51669;
    wire N__51666;
    wire N__51663;
    wire N__51660;
    wire N__51657;
    wire N__51656;
    wire N__51653;
    wire N__51652;
    wire N__51649;
    wire N__51646;
    wire N__51643;
    wire N__51640;
    wire N__51637;
    wire N__51634;
    wire N__51631;
    wire N__51624;
    wire N__51621;
    wire N__51620;
    wire N__51617;
    wire N__51614;
    wire N__51611;
    wire N__51610;
    wire N__51607;
    wire N__51604;
    wire N__51601;
    wire N__51598;
    wire N__51591;
    wire N__51588;
    wire N__51587;
    wire N__51586;
    wire N__51583;
    wire N__51580;
    wire N__51577;
    wire N__51574;
    wire N__51571;
    wire N__51568;
    wire N__51565;
    wire N__51562;
    wire N__51555;
    wire N__51552;
    wire N__51549;
    wire N__51546;
    wire N__51543;
    wire N__51540;
    wire N__51537;
    wire N__51534;
    wire N__51531;
    wire N__51528;
    wire N__51525;
    wire N__51522;
    wire N__51519;
    wire N__51516;
    wire N__51513;
    wire N__51510;
    wire N__51507;
    wire N__51506;
    wire N__51505;
    wire N__51502;
    wire N__51499;
    wire N__51496;
    wire N__51493;
    wire N__51490;
    wire N__51487;
    wire N__51482;
    wire N__51477;
    wire N__51476;
    wire N__51473;
    wire N__51470;
    wire N__51467;
    wire N__51464;
    wire N__51463;
    wire N__51460;
    wire N__51457;
    wire N__51454;
    wire N__51447;
    wire N__51444;
    wire N__51441;
    wire N__51438;
    wire N__51435;
    wire N__51434;
    wire N__51431;
    wire N__51430;
    wire N__51427;
    wire N__51424;
    wire N__51421;
    wire N__51418;
    wire N__51415;
    wire N__51412;
    wire N__51409;
    wire N__51402;
    wire N__51399;
    wire N__51396;
    wire N__51395;
    wire N__51392;
    wire N__51389;
    wire N__51386;
    wire N__51383;
    wire N__51382;
    wire N__51377;
    wire N__51374;
    wire N__51369;
    wire N__51368;
    wire N__51365;
    wire N__51364;
    wire N__51361;
    wire N__51358;
    wire N__51355;
    wire N__51352;
    wire N__51347;
    wire N__51342;
    wire N__51339;
    wire N__51336;
    wire N__51333;
    wire N__51330;
    wire N__51327;
    wire N__51324;
    wire N__51321;
    wire N__51318;
    wire N__51315;
    wire N__51312;
    wire N__51309;
    wire N__51306;
    wire N__51303;
    wire N__51300;
    wire N__51299;
    wire N__51296;
    wire N__51293;
    wire N__51290;
    wire N__51285;
    wire N__51282;
    wire N__51279;
    wire N__51276;
    wire N__51273;
    wire N__51270;
    wire N__51267;
    wire N__51264;
    wire N__51261;
    wire N__51258;
    wire N__51255;
    wire N__51252;
    wire N__51251;
    wire N__51248;
    wire N__51245;
    wire N__51242;
    wire N__51241;
    wire N__51238;
    wire N__51235;
    wire N__51232;
    wire N__51229;
    wire N__51224;
    wire N__51221;
    wire N__51218;
    wire N__51213;
    wire N__51210;
    wire N__51207;
    wire N__51206;
    wire N__51203;
    wire N__51200;
    wire N__51197;
    wire N__51194;
    wire N__51191;
    wire N__51190;
    wire N__51187;
    wire N__51186;
    wire N__51183;
    wire N__51180;
    wire N__51177;
    wire N__51174;
    wire N__51171;
    wire N__51168;
    wire N__51163;
    wire N__51160;
    wire N__51157;
    wire N__51154;
    wire N__51151;
    wire N__51148;
    wire N__51145;
    wire N__51142;
    wire N__51139;
    wire N__51136;
    wire N__51129;
    wire N__51126;
    wire N__51123;
    wire N__51122;
    wire N__51121;
    wire N__51120;
    wire N__51119;
    wire N__51118;
    wire N__51113;
    wire N__51104;
    wire N__51101;
    wire N__51098;
    wire N__51095;
    wire N__51092;
    wire N__51089;
    wire N__51086;
    wire N__51081;
    wire N__51080;
    wire N__51079;
    wire N__51078;
    wire N__51077;
    wire N__51076;
    wire N__51075;
    wire N__51070;
    wire N__51059;
    wire N__51054;
    wire N__51053;
    wire N__51052;
    wire N__51049;
    wire N__51048;
    wire N__51045;
    wire N__51044;
    wire N__51037;
    wire N__51032;
    wire N__51029;
    wire N__51024;
    wire N__51023;
    wire N__51022;
    wire N__51019;
    wire N__51016;
    wire N__51015;
    wire N__51014;
    wire N__51013;
    wire N__51008;
    wire N__50999;
    wire N__50994;
    wire N__50993;
    wire N__50990;
    wire N__50987;
    wire N__50984;
    wire N__50983;
    wire N__50980;
    wire N__50979;
    wire N__50976;
    wire N__50973;
    wire N__50970;
    wire N__50967;
    wire N__50960;
    wire N__50955;
    wire N__50952;
    wire N__50949;
    wire N__50946;
    wire N__50943;
    wire N__50940;
    wire N__50937;
    wire N__50934;
    wire N__50933;
    wire N__50932;
    wire N__50931;
    wire N__50930;
    wire N__50927;
    wire N__50924;
    wire N__50923;
    wire N__50922;
    wire N__50921;
    wire N__50914;
    wire N__50909;
    wire N__50902;
    wire N__50899;
    wire N__50896;
    wire N__50893;
    wire N__50886;
    wire N__50885;
    wire N__50884;
    wire N__50883;
    wire N__50882;
    wire N__50881;
    wire N__50878;
    wire N__50875;
    wire N__50874;
    wire N__50873;
    wire N__50872;
    wire N__50871;
    wire N__50866;
    wire N__50865;
    wire N__50864;
    wire N__50861;
    wire N__50858;
    wire N__50855;
    wire N__50844;
    wire N__50841;
    wire N__50836;
    wire N__50833;
    wire N__50830;
    wire N__50821;
    wire N__50820;
    wire N__50817;
    wire N__50814;
    wire N__50811;
    wire N__50808;
    wire N__50805;
    wire N__50802;
    wire N__50797;
    wire N__50790;
    wire N__50787;
    wire N__50784;
    wire N__50781;
    wire N__50778;
    wire N__50775;
    wire N__50772;
    wire N__50769;
    wire N__50766;
    wire N__50763;
    wire N__50760;
    wire N__50757;
    wire N__50754;
    wire N__50751;
    wire N__50748;
    wire N__50747;
    wire N__50746;
    wire N__50743;
    wire N__50738;
    wire N__50735;
    wire N__50732;
    wire N__50727;
    wire N__50724;
    wire N__50721;
    wire N__50718;
    wire N__50717;
    wire N__50716;
    wire N__50715;
    wire N__50714;
    wire N__50711;
    wire N__50706;
    wire N__50701;
    wire N__50698;
    wire N__50693;
    wire N__50690;
    wire N__50687;
    wire N__50682;
    wire N__50681;
    wire N__50678;
    wire N__50675;
    wire N__50670;
    wire N__50667;
    wire N__50666;
    wire N__50663;
    wire N__50660;
    wire N__50655;
    wire N__50652;
    wire N__50649;
    wire N__50646;
    wire N__50643;
    wire N__50642;
    wire N__50637;
    wire N__50634;
    wire N__50631;
    wire N__50628;
    wire N__50625;
    wire N__50622;
    wire N__50621;
    wire N__50618;
    wire N__50615;
    wire N__50612;
    wire N__50611;
    wire N__50608;
    wire N__50605;
    wire N__50602;
    wire N__50597;
    wire N__50592;
    wire N__50589;
    wire N__50586;
    wire N__50585;
    wire N__50582;
    wire N__50581;
    wire N__50578;
    wire N__50575;
    wire N__50572;
    wire N__50565;
    wire N__50562;
    wire N__50559;
    wire N__50558;
    wire N__50555;
    wire N__50552;
    wire N__50551;
    wire N__50546;
    wire N__50545;
    wire N__50544;
    wire N__50543;
    wire N__50540;
    wire N__50539;
    wire N__50538;
    wire N__50537;
    wire N__50536;
    wire N__50533;
    wire N__50530;
    wire N__50525;
    wire N__50522;
    wire N__50517;
    wire N__50512;
    wire N__50509;
    wire N__50506;
    wire N__50493;
    wire N__50490;
    wire N__50487;
    wire N__50484;
    wire N__50481;
    wire N__50478;
    wire N__50475;
    wire N__50472;
    wire N__50469;
    wire N__50466;
    wire N__50463;
    wire N__50460;
    wire N__50457;
    wire N__50456;
    wire N__50453;
    wire N__50450;
    wire N__50449;
    wire N__50446;
    wire N__50443;
    wire N__50440;
    wire N__50437;
    wire N__50434;
    wire N__50427;
    wire N__50424;
    wire N__50421;
    wire N__50418;
    wire N__50415;
    wire N__50412;
    wire N__50409;
    wire N__50408;
    wire N__50407;
    wire N__50406;
    wire N__50405;
    wire N__50404;
    wire N__50403;
    wire N__50402;
    wire N__50401;
    wire N__50398;
    wire N__50397;
    wire N__50396;
    wire N__50395;
    wire N__50394;
    wire N__50393;
    wire N__50392;
    wire N__50391;
    wire N__50390;
    wire N__50389;
    wire N__50388;
    wire N__50387;
    wire N__50386;
    wire N__50381;
    wire N__50380;
    wire N__50379;
    wire N__50368;
    wire N__50359;
    wire N__50356;
    wire N__50355;
    wire N__50354;
    wire N__50353;
    wire N__50352;
    wire N__50351;
    wire N__50350;
    wire N__50349;
    wire N__50348;
    wire N__50347;
    wire N__50334;
    wire N__50329;
    wire N__50326;
    wire N__50323;
    wire N__50318;
    wire N__50313;
    wire N__50308;
    wire N__50301;
    wire N__50290;
    wire N__50285;
    wire N__50282;
    wire N__50277;
    wire N__50274;
    wire N__50265;
    wire N__50262;
    wire N__50257;
    wire N__50254;
    wire N__50251;
    wire N__50248;
    wire N__50245;
    wire N__50244;
    wire N__50239;
    wire N__50236;
    wire N__50233;
    wire N__50226;
    wire N__50223;
    wire N__50220;
    wire N__50219;
    wire N__50218;
    wire N__50215;
    wire N__50208;
    wire N__50205;
    wire N__50202;
    wire N__50199;
    wire N__50196;
    wire N__50193;
    wire N__50192;
    wire N__50191;
    wire N__50188;
    wire N__50185;
    wire N__50182;
    wire N__50175;
    wire N__50172;
    wire N__50169;
    wire N__50166;
    wire N__50163;
    wire N__50160;
    wire N__50157;
    wire N__50154;
    wire N__50151;
    wire N__50148;
    wire N__50145;
    wire N__50142;
    wire N__50141;
    wire N__50140;
    wire N__50139;
    wire N__50138;
    wire N__50137;
    wire N__50134;
    wire N__50131;
    wire N__50126;
    wire N__50121;
    wire N__50114;
    wire N__50113;
    wire N__50112;
    wire N__50109;
    wire N__50106;
    wire N__50103;
    wire N__50100;
    wire N__50091;
    wire N__50088;
    wire N__50087;
    wire N__50084;
    wire N__50081;
    wire N__50080;
    wire N__50077;
    wire N__50076;
    wire N__50073;
    wire N__50070;
    wire N__50067;
    wire N__50064;
    wire N__50061;
    wire N__50058;
    wire N__50053;
    wire N__50052;
    wire N__50051;
    wire N__50050;
    wire N__50049;
    wire N__50046;
    wire N__50043;
    wire N__50040;
    wire N__50037;
    wire N__50030;
    wire N__50019;
    wire N__50016;
    wire N__50015;
    wire N__50012;
    wire N__50009;
    wire N__50004;
    wire N__50001;
    wire N__49998;
    wire N__49997;
    wire N__49994;
    wire N__49991;
    wire N__49986;
    wire N__49983;
    wire N__49980;
    wire N__49977;
    wire N__49974;
    wire N__49971;
    wire N__49968;
    wire N__49965;
    wire N__49962;
    wire N__49961;
    wire N__49958;
    wire N__49955;
    wire N__49952;
    wire N__49949;
    wire N__49948;
    wire N__49943;
    wire N__49940;
    wire N__49935;
    wire N__49932;
    wire N__49929;
    wire N__49926;
    wire N__49923;
    wire N__49920;
    wire N__49917;
    wire N__49914;
    wire N__49911;
    wire N__49908;
    wire N__49905;
    wire N__49902;
    wire N__49899;
    wire N__49896;
    wire N__49893;
    wire N__49890;
    wire N__49887;
    wire N__49884;
    wire N__49881;
    wire N__49878;
    wire N__49875;
    wire N__49872;
    wire N__49869;
    wire N__49866;
    wire N__49863;
    wire N__49860;
    wire N__49857;
    wire N__49854;
    wire N__49851;
    wire N__49848;
    wire N__49845;
    wire N__49842;
    wire N__49839;
    wire N__49836;
    wire N__49833;
    wire N__49832;
    wire N__49829;
    wire N__49826;
    wire N__49823;
    wire N__49820;
    wire N__49819;
    wire N__49816;
    wire N__49813;
    wire N__49810;
    wire N__49803;
    wire N__49800;
    wire N__49797;
    wire N__49794;
    wire N__49791;
    wire N__49788;
    wire N__49785;
    wire N__49782;
    wire N__49779;
    wire N__49776;
    wire N__49773;
    wire N__49770;
    wire N__49767;
    wire N__49764;
    wire N__49761;
    wire N__49758;
    wire N__49755;
    wire N__49752;
    wire N__49751;
    wire N__49748;
    wire N__49747;
    wire N__49744;
    wire N__49741;
    wire N__49738;
    wire N__49735;
    wire N__49732;
    wire N__49729;
    wire N__49726;
    wire N__49719;
    wire N__49718;
    wire N__49715;
    wire N__49712;
    wire N__49709;
    wire N__49706;
    wire N__49703;
    wire N__49700;
    wire N__49697;
    wire N__49694;
    wire N__49693;
    wire N__49690;
    wire N__49687;
    wire N__49684;
    wire N__49677;
    wire N__49676;
    wire N__49673;
    wire N__49670;
    wire N__49669;
    wire N__49666;
    wire N__49663;
    wire N__49660;
    wire N__49657;
    wire N__49654;
    wire N__49651;
    wire N__49648;
    wire N__49641;
    wire N__49638;
    wire N__49637;
    wire N__49636;
    wire N__49633;
    wire N__49630;
    wire N__49627;
    wire N__49624;
    wire N__49621;
    wire N__49618;
    wire N__49615;
    wire N__49612;
    wire N__49609;
    wire N__49602;
    wire N__49599;
    wire N__49596;
    wire N__49593;
    wire N__49590;
    wire N__49587;
    wire N__49584;
    wire N__49581;
    wire N__49578;
    wire N__49575;
    wire N__49572;
    wire N__49569;
    wire N__49566;
    wire N__49563;
    wire N__49560;
    wire N__49557;
    wire N__49554;
    wire N__49551;
    wire N__49548;
    wire N__49545;
    wire N__49542;
    wire N__49539;
    wire N__49536;
    wire N__49533;
    wire N__49530;
    wire N__49527;
    wire N__49524;
    wire N__49521;
    wire N__49518;
    wire N__49515;
    wire N__49512;
    wire N__49509;
    wire N__49506;
    wire N__49503;
    wire N__49500;
    wire N__49497;
    wire N__49494;
    wire N__49493;
    wire N__49490;
    wire N__49487;
    wire N__49484;
    wire N__49481;
    wire N__49480;
    wire N__49477;
    wire N__49474;
    wire N__49471;
    wire N__49464;
    wire N__49461;
    wire N__49458;
    wire N__49455;
    wire N__49454;
    wire N__49453;
    wire N__49450;
    wire N__49447;
    wire N__49444;
    wire N__49437;
    wire N__49434;
    wire N__49431;
    wire N__49428;
    wire N__49427;
    wire N__49424;
    wire N__49423;
    wire N__49420;
    wire N__49417;
    wire N__49414;
    wire N__49411;
    wire N__49408;
    wire N__49405;
    wire N__49402;
    wire N__49399;
    wire N__49394;
    wire N__49391;
    wire N__49386;
    wire N__49383;
    wire N__49382;
    wire N__49379;
    wire N__49378;
    wire N__49375;
    wire N__49372;
    wire N__49369;
    wire N__49366;
    wire N__49363;
    wire N__49360;
    wire N__49357;
    wire N__49354;
    wire N__49349;
    wire N__49344;
    wire N__49341;
    wire N__49340;
    wire N__49339;
    wire N__49336;
    wire N__49333;
    wire N__49330;
    wire N__49327;
    wire N__49324;
    wire N__49321;
    wire N__49318;
    wire N__49313;
    wire N__49308;
    wire N__49307;
    wire N__49304;
    wire N__49301;
    wire N__49298;
    wire N__49295;
    wire N__49292;
    wire N__49289;
    wire N__49286;
    wire N__49285;
    wire N__49282;
    wire N__49279;
    wire N__49276;
    wire N__49269;
    wire N__49268;
    wire N__49265;
    wire N__49262;
    wire N__49259;
    wire N__49256;
    wire N__49255;
    wire N__49252;
    wire N__49249;
    wire N__49246;
    wire N__49241;
    wire N__49238;
    wire N__49233;
    wire N__49230;
    wire N__49227;
    wire N__49224;
    wire N__49221;
    wire N__49218;
    wire N__49215;
    wire N__49212;
    wire N__49209;
    wire N__49206;
    wire N__49203;
    wire N__49200;
    wire N__49197;
    wire N__49194;
    wire N__49191;
    wire N__49188;
    wire N__49185;
    wire N__49182;
    wire N__49179;
    wire N__49176;
    wire N__49173;
    wire N__49170;
    wire N__49167;
    wire N__49164;
    wire N__49163;
    wire N__49160;
    wire N__49157;
    wire N__49156;
    wire N__49153;
    wire N__49148;
    wire N__49143;
    wire N__49140;
    wire N__49137;
    wire N__49134;
    wire N__49131;
    wire N__49128;
    wire N__49125;
    wire N__49122;
    wire N__49119;
    wire N__49116;
    wire N__49113;
    wire N__49110;
    wire N__49107;
    wire N__49104;
    wire N__49101;
    wire N__49098;
    wire N__49095;
    wire N__49094;
    wire N__49093;
    wire N__49090;
    wire N__49087;
    wire N__49084;
    wire N__49083;
    wire N__49080;
    wire N__49075;
    wire N__49072;
    wire N__49071;
    wire N__49064;
    wire N__49063;
    wire N__49060;
    wire N__49059;
    wire N__49056;
    wire N__49053;
    wire N__49050;
    wire N__49047;
    wire N__49044;
    wire N__49041;
    wire N__49038;
    wire N__49035;
    wire N__49034;
    wire N__49033;
    wire N__49028;
    wire N__49023;
    wire N__49020;
    wire N__49017;
    wire N__49008;
    wire N__49005;
    wire N__49004;
    wire N__49003;
    wire N__49000;
    wire N__48997;
    wire N__48994;
    wire N__48991;
    wire N__48988;
    wire N__48985;
    wire N__48982;
    wire N__48975;
    wire N__48974;
    wire N__48971;
    wire N__48968;
    wire N__48965;
    wire N__48964;
    wire N__48961;
    wire N__48958;
    wire N__48955;
    wire N__48950;
    wire N__48945;
    wire N__48942;
    wire N__48939;
    wire N__48936;
    wire N__48935;
    wire N__48934;
    wire N__48931;
    wire N__48926;
    wire N__48921;
    wire N__48918;
    wire N__48915;
    wire N__48914;
    wire N__48911;
    wire N__48910;
    wire N__48907;
    wire N__48904;
    wire N__48901;
    wire N__48898;
    wire N__48891;
    wire N__48888;
    wire N__48885;
    wire N__48882;
    wire N__48879;
    wire N__48878;
    wire N__48875;
    wire N__48872;
    wire N__48867;
    wire N__48866;
    wire N__48863;
    wire N__48862;
    wire N__48859;
    wire N__48856;
    wire N__48853;
    wire N__48848;
    wire N__48845;
    wire N__48842;
    wire N__48837;
    wire N__48834;
    wire N__48831;
    wire N__48828;
    wire N__48825;
    wire N__48822;
    wire N__48819;
    wire N__48816;
    wire N__48813;
    wire N__48810;
    wire N__48807;
    wire N__48804;
    wire N__48801;
    wire N__48798;
    wire N__48795;
    wire N__48792;
    wire N__48789;
    wire N__48786;
    wire N__48783;
    wire N__48780;
    wire N__48777;
    wire N__48774;
    wire N__48771;
    wire N__48768;
    wire N__48765;
    wire N__48762;
    wire N__48759;
    wire N__48756;
    wire N__48753;
    wire N__48750;
    wire N__48749;
    wire N__48746;
    wire N__48745;
    wire N__48742;
    wire N__48739;
    wire N__48736;
    wire N__48733;
    wire N__48726;
    wire N__48725;
    wire N__48724;
    wire N__48723;
    wire N__48722;
    wire N__48711;
    wire N__48708;
    wire N__48705;
    wire N__48702;
    wire N__48701;
    wire N__48698;
    wire N__48695;
    wire N__48694;
    wire N__48691;
    wire N__48686;
    wire N__48681;
    wire N__48678;
    wire N__48677;
    wire N__48674;
    wire N__48671;
    wire N__48670;
    wire N__48667;
    wire N__48664;
    wire N__48661;
    wire N__48654;
    wire N__48653;
    wire N__48652;
    wire N__48651;
    wire N__48642;
    wire N__48641;
    wire N__48640;
    wire N__48639;
    wire N__48638;
    wire N__48635;
    wire N__48626;
    wire N__48621;
    wire N__48618;
    wire N__48617;
    wire N__48616;
    wire N__48613;
    wire N__48610;
    wire N__48607;
    wire N__48600;
    wire N__48597;
    wire N__48594;
    wire N__48591;
    wire N__48588;
    wire N__48585;
    wire N__48582;
    wire N__48581;
    wire N__48578;
    wire N__48575;
    wire N__48572;
    wire N__48569;
    wire N__48566;
    wire N__48565;
    wire N__48562;
    wire N__48559;
    wire N__48556;
    wire N__48551;
    wire N__48548;
    wire N__48545;
    wire N__48542;
    wire N__48537;
    wire N__48534;
    wire N__48531;
    wire N__48528;
    wire N__48525;
    wire N__48522;
    wire N__48519;
    wire N__48516;
    wire N__48513;
    wire N__48510;
    wire N__48507;
    wire N__48504;
    wire N__48501;
    wire N__48498;
    wire N__48495;
    wire N__48492;
    wire N__48489;
    wire N__48486;
    wire N__48483;
    wire N__48482;
    wire N__48479;
    wire N__48478;
    wire N__48475;
    wire N__48472;
    wire N__48469;
    wire N__48462;
    wire N__48459;
    wire N__48458;
    wire N__48457;
    wire N__48454;
    wire N__48451;
    wire N__48448;
    wire N__48445;
    wire N__48438;
    wire N__48435;
    wire N__48434;
    wire N__48431;
    wire N__48430;
    wire N__48427;
    wire N__48424;
    wire N__48421;
    wire N__48414;
    wire N__48411;
    wire N__48410;
    wire N__48409;
    wire N__48406;
    wire N__48401;
    wire N__48396;
    wire N__48393;
    wire N__48392;
    wire N__48391;
    wire N__48388;
    wire N__48383;
    wire N__48378;
    wire N__48375;
    wire N__48374;
    wire N__48373;
    wire N__48370;
    wire N__48365;
    wire N__48360;
    wire N__48357;
    wire N__48356;
    wire N__48355;
    wire N__48352;
    wire N__48349;
    wire N__48346;
    wire N__48343;
    wire N__48340;
    wire N__48333;
    wire N__48330;
    wire N__48329;
    wire N__48326;
    wire N__48325;
    wire N__48322;
    wire N__48317;
    wire N__48314;
    wire N__48311;
    wire N__48310;
    wire N__48307;
    wire N__48304;
    wire N__48301;
    wire N__48294;
    wire N__48293;
    wire N__48292;
    wire N__48291;
    wire N__48290;
    wire N__48287;
    wire N__48284;
    wire N__48281;
    wire N__48278;
    wire N__48275;
    wire N__48272;
    wire N__48263;
    wire N__48262;
    wire N__48259;
    wire N__48258;
    wire N__48257;
    wire N__48256;
    wire N__48253;
    wire N__48250;
    wire N__48247;
    wire N__48244;
    wire N__48241;
    wire N__48238;
    wire N__48235;
    wire N__48222;
    wire N__48221;
    wire N__48220;
    wire N__48219;
    wire N__48216;
    wire N__48213;
    wire N__48210;
    wire N__48209;
    wire N__48206;
    wire N__48205;
    wire N__48196;
    wire N__48195;
    wire N__48190;
    wire N__48187;
    wire N__48184;
    wire N__48183;
    wire N__48182;
    wire N__48181;
    wire N__48174;
    wire N__48167;
    wire N__48162;
    wire N__48159;
    wire N__48158;
    wire N__48157;
    wire N__48156;
    wire N__48153;
    wire N__48150;
    wire N__48147;
    wire N__48144;
    wire N__48141;
    wire N__48140;
    wire N__48133;
    wire N__48132;
    wire N__48129;
    wire N__48126;
    wire N__48123;
    wire N__48120;
    wire N__48111;
    wire N__48108;
    wire N__48107;
    wire N__48106;
    wire N__48105;
    wire N__48102;
    wire N__48099;
    wire N__48096;
    wire N__48093;
    wire N__48090;
    wire N__48085;
    wire N__48082;
    wire N__48081;
    wire N__48080;
    wire N__48077;
    wire N__48074;
    wire N__48071;
    wire N__48066;
    wire N__48057;
    wire N__48056;
    wire N__48053;
    wire N__48050;
    wire N__48049;
    wire N__48048;
    wire N__48045;
    wire N__48042;
    wire N__48039;
    wire N__48036;
    wire N__48033;
    wire N__48032;
    wire N__48029;
    wire N__48024;
    wire N__48021;
    wire N__48020;
    wire N__48017;
    wire N__48014;
    wire N__48009;
    wire N__48006;
    wire N__47997;
    wire N__47996;
    wire N__47995;
    wire N__47994;
    wire N__47993;
    wire N__47992;
    wire N__47991;
    wire N__47990;
    wire N__47989;
    wire N__47988;
    wire N__47987;
    wire N__47986;
    wire N__47985;
    wire N__47984;
    wire N__47983;
    wire N__47982;
    wire N__47981;
    wire N__47980;
    wire N__47979;
    wire N__47978;
    wire N__47937;
    wire N__47934;
    wire N__47931;
    wire N__47928;
    wire N__47925;
    wire N__47922;
    wire N__47921;
    wire N__47918;
    wire N__47915;
    wire N__47914;
    wire N__47913;
    wire N__47912;
    wire N__47907;
    wire N__47904;
    wire N__47899;
    wire N__47892;
    wire N__47889;
    wire N__47886;
    wire N__47883;
    wire N__47882;
    wire N__47881;
    wire N__47880;
    wire N__47879;
    wire N__47878;
    wire N__47877;
    wire N__47876;
    wire N__47875;
    wire N__47874;
    wire N__47873;
    wire N__47872;
    wire N__47871;
    wire N__47870;
    wire N__47869;
    wire N__47868;
    wire N__47867;
    wire N__47866;
    wire N__47865;
    wire N__47864;
    wire N__47863;
    wire N__47860;
    wire N__47859;
    wire N__47858;
    wire N__47857;
    wire N__47856;
    wire N__47855;
    wire N__47854;
    wire N__47853;
    wire N__47852;
    wire N__47851;
    wire N__47850;
    wire N__47849;
    wire N__47848;
    wire N__47847;
    wire N__47846;
    wire N__47845;
    wire N__47844;
    wire N__47843;
    wire N__47842;
    wire N__47833;
    wire N__47828;
    wire N__47823;
    wire N__47820;
    wire N__47815;
    wire N__47814;
    wire N__47813;
    wire N__47812;
    wire N__47811;
    wire N__47810;
    wire N__47803;
    wire N__47798;
    wire N__47795;
    wire N__47788;
    wire N__47785;
    wire N__47778;
    wire N__47771;
    wire N__47764;
    wire N__47759;
    wire N__47756;
    wire N__47743;
    wire N__47742;
    wire N__47741;
    wire N__47732;
    wire N__47731;
    wire N__47730;
    wire N__47729;
    wire N__47728;
    wire N__47727;
    wire N__47726;
    wire N__47725;
    wire N__47724;
    wire N__47721;
    wire N__47716;
    wire N__47711;
    wire N__47708;
    wire N__47707;
    wire N__47706;
    wire N__47703;
    wire N__47696;
    wire N__47681;
    wire N__47676;
    wire N__47673;
    wire N__47664;
    wire N__47655;
    wire N__47654;
    wire N__47653;
    wire N__47652;
    wire N__47651;
    wire N__47650;
    wire N__47649;
    wire N__47648;
    wire N__47647;
    wire N__47646;
    wire N__47645;
    wire N__47644;
    wire N__47639;
    wire N__47634;
    wire N__47629;
    wire N__47620;
    wire N__47613;
    wire N__47602;
    wire N__47591;
    wire N__47588;
    wire N__47571;
    wire N__47568;
    wire N__47565;
    wire N__47564;
    wire N__47563;
    wire N__47562;
    wire N__47557;
    wire N__47552;
    wire N__47547;
    wire N__47546;
    wire N__47545;
    wire N__47538;
    wire N__47535;
    wire N__47532;
    wire N__47529;
    wire N__47526;
    wire N__47523;
    wire N__47520;
    wire N__47517;
    wire N__47514;
    wire N__47511;
    wire N__47510;
    wire N__47507;
    wire N__47504;
    wire N__47501;
    wire N__47498;
    wire N__47493;
    wire N__47490;
    wire N__47487;
    wire N__47484;
    wire N__47481;
    wire N__47478;
    wire N__47475;
    wire N__47472;
    wire N__47469;
    wire N__47468;
    wire N__47463;
    wire N__47460;
    wire N__47457;
    wire N__47456;
    wire N__47453;
    wire N__47450;
    wire N__47445;
    wire N__47442;
    wire N__47439;
    wire N__47436;
    wire N__47433;
    wire N__47430;
    wire N__47427;
    wire N__47426;
    wire N__47423;
    wire N__47420;
    wire N__47415;
    wire N__47414;
    wire N__47413;
    wire N__47412;
    wire N__47411;
    wire N__47410;
    wire N__47409;
    wire N__47404;
    wire N__47403;
    wire N__47400;
    wire N__47391;
    wire N__47388;
    wire N__47385;
    wire N__47384;
    wire N__47383;
    wire N__47382;
    wire N__47381;
    wire N__47380;
    wire N__47379;
    wire N__47378;
    wire N__47375;
    wire N__47372;
    wire N__47369;
    wire N__47366;
    wire N__47357;
    wire N__47350;
    wire N__47347;
    wire N__47344;
    wire N__47341;
    wire N__47328;
    wire N__47325;
    wire N__47322;
    wire N__47319;
    wire N__47316;
    wire N__47313;
    wire N__47310;
    wire N__47307;
    wire N__47304;
    wire N__47301;
    wire N__47298;
    wire N__47295;
    wire N__47292;
    wire N__47289;
    wire N__47286;
    wire N__47283;
    wire N__47280;
    wire N__47277;
    wire N__47274;
    wire N__47271;
    wire N__47268;
    wire N__47265;
    wire N__47262;
    wire N__47259;
    wire N__47256;
    wire N__47253;
    wire N__47250;
    wire N__47247;
    wire N__47246;
    wire N__47245;
    wire N__47244;
    wire N__47243;
    wire N__47240;
    wire N__47237;
    wire N__47232;
    wire N__47229;
    wire N__47222;
    wire N__47219;
    wire N__47216;
    wire N__47213;
    wire N__47208;
    wire N__47207;
    wire N__47206;
    wire N__47201;
    wire N__47198;
    wire N__47197;
    wire N__47196;
    wire N__47193;
    wire N__47190;
    wire N__47187;
    wire N__47184;
    wire N__47179;
    wire N__47172;
    wire N__47171;
    wire N__47170;
    wire N__47169;
    wire N__47168;
    wire N__47165;
    wire N__47164;
    wire N__47161;
    wire N__47158;
    wire N__47153;
    wire N__47150;
    wire N__47147;
    wire N__47140;
    wire N__47137;
    wire N__47134;
    wire N__47129;
    wire N__47124;
    wire N__47123;
    wire N__47122;
    wire N__47119;
    wire N__47118;
    wire N__47115;
    wire N__47112;
    wire N__47111;
    wire N__47110;
    wire N__47107;
    wire N__47104;
    wire N__47099;
    wire N__47094;
    wire N__47093;
    wire N__47090;
    wire N__47085;
    wire N__47082;
    wire N__47079;
    wire N__47076;
    wire N__47073;
    wire N__47068;
    wire N__47061;
    wire N__47058;
    wire N__47055;
    wire N__47052;
    wire N__47049;
    wire N__47046;
    wire N__47043;
    wire N__47042;
    wire N__47041;
    wire N__47038;
    wire N__47037;
    wire N__47034;
    wire N__47031;
    wire N__47028;
    wire N__47025;
    wire N__47018;
    wire N__47013;
    wire N__47012;
    wire N__47009;
    wire N__47008;
    wire N__47007;
    wire N__47004;
    wire N__47001;
    wire N__46998;
    wire N__46995;
    wire N__46992;
    wire N__46989;
    wire N__46980;
    wire N__46977;
    wire N__46974;
    wire N__46971;
    wire N__46968;
    wire N__46965;
    wire N__46962;
    wire N__46959;
    wire N__46956;
    wire N__46953;
    wire N__46950;
    wire N__46947;
    wire N__46946;
    wire N__46943;
    wire N__46942;
    wire N__46939;
    wire N__46938;
    wire N__46935;
    wire N__46932;
    wire N__46929;
    wire N__46926;
    wire N__46923;
    wire N__46914;
    wire N__46911;
    wire N__46910;
    wire N__46909;
    wire N__46908;
    wire N__46907;
    wire N__46904;
    wire N__46901;
    wire N__46900;
    wire N__46897;
    wire N__46896;
    wire N__46893;
    wire N__46892;
    wire N__46891;
    wire N__46888;
    wire N__46885;
    wire N__46876;
    wire N__46869;
    wire N__46866;
    wire N__46863;
    wire N__46860;
    wire N__46857;
    wire N__46854;
    wire N__46849;
    wire N__46846;
    wire N__46843;
    wire N__46840;
    wire N__46837;
    wire N__46832;
    wire N__46829;
    wire N__46824;
    wire N__46821;
    wire N__46818;
    wire N__46817;
    wire N__46814;
    wire N__46813;
    wire N__46812;
    wire N__46811;
    wire N__46808;
    wire N__46807;
    wire N__46804;
    wire N__46799;
    wire N__46796;
    wire N__46793;
    wire N__46790;
    wire N__46787;
    wire N__46782;
    wire N__46779;
    wire N__46772;
    wire N__46769;
    wire N__46764;
    wire N__46763;
    wire N__46762;
    wire N__46761;
    wire N__46760;
    wire N__46757;
    wire N__46756;
    wire N__46753;
    wire N__46746;
    wire N__46743;
    wire N__46740;
    wire N__46737;
    wire N__46732;
    wire N__46725;
    wire N__46722;
    wire N__46719;
    wire N__46716;
    wire N__46713;
    wire N__46710;
    wire N__46707;
    wire N__46704;
    wire N__46701;
    wire N__46698;
    wire N__46695;
    wire N__46692;
    wire N__46689;
    wire N__46686;
    wire N__46683;
    wire N__46680;
    wire N__46677;
    wire N__46674;
    wire N__46671;
    wire N__46668;
    wire N__46667;
    wire N__46664;
    wire N__46661;
    wire N__46660;
    wire N__46657;
    wire N__46654;
    wire N__46651;
    wire N__46644;
    wire N__46641;
    wire N__46638;
    wire N__46635;
    wire N__46634;
    wire N__46631;
    wire N__46628;
    wire N__46627;
    wire N__46624;
    wire N__46619;
    wire N__46614;
    wire N__46611;
    wire N__46608;
    wire N__46605;
    wire N__46602;
    wire N__46599;
    wire N__46598;
    wire N__46597;
    wire N__46594;
    wire N__46589;
    wire N__46586;
    wire N__46583;
    wire N__46578;
    wire N__46575;
    wire N__46572;
    wire N__46569;
    wire N__46566;
    wire N__46563;
    wire N__46560;
    wire N__46557;
    wire N__46556;
    wire N__46553;
    wire N__46552;
    wire N__46549;
    wire N__46546;
    wire N__46541;
    wire N__46538;
    wire N__46535;
    wire N__46530;
    wire N__46527;
    wire N__46526;
    wire N__46525;
    wire N__46524;
    wire N__46523;
    wire N__46520;
    wire N__46517;
    wire N__46514;
    wire N__46511;
    wire N__46508;
    wire N__46507;
    wire N__46502;
    wire N__46501;
    wire N__46500;
    wire N__46497;
    wire N__46494;
    wire N__46491;
    wire N__46488;
    wire N__46485;
    wire N__46482;
    wire N__46479;
    wire N__46476;
    wire N__46471;
    wire N__46468;
    wire N__46465;
    wire N__46462;
    wire N__46461;
    wire N__46458;
    wire N__46453;
    wire N__46450;
    wire N__46447;
    wire N__46444;
    wire N__46441;
    wire N__46438;
    wire N__46435;
    wire N__46428;
    wire N__46419;
    wire N__46416;
    wire N__46413;
    wire N__46410;
    wire N__46407;
    wire N__46404;
    wire N__46401;
    wire N__46398;
    wire N__46395;
    wire N__46392;
    wire N__46389;
    wire N__46386;
    wire N__46383;
    wire N__46380;
    wire N__46377;
    wire N__46376;
    wire N__46373;
    wire N__46370;
    wire N__46369;
    wire N__46366;
    wire N__46363;
    wire N__46360;
    wire N__46355;
    wire N__46350;
    wire N__46347;
    wire N__46346;
    wire N__46343;
    wire N__46340;
    wire N__46339;
    wire N__46336;
    wire N__46333;
    wire N__46330;
    wire N__46327;
    wire N__46322;
    wire N__46317;
    wire N__46314;
    wire N__46311;
    wire N__46308;
    wire N__46307;
    wire N__46306;
    wire N__46303;
    wire N__46298;
    wire N__46293;
    wire N__46290;
    wire N__46287;
    wire N__46284;
    wire N__46281;
    wire N__46278;
    wire N__46275;
    wire N__46272;
    wire N__46271;
    wire N__46270;
    wire N__46267;
    wire N__46264;
    wire N__46261;
    wire N__46258;
    wire N__46255;
    wire N__46252;
    wire N__46249;
    wire N__46246;
    wire N__46243;
    wire N__46240;
    wire N__46237;
    wire N__46234;
    wire N__46227;
    wire N__46224;
    wire N__46221;
    wire N__46218;
    wire N__46215;
    wire N__46212;
    wire N__46211;
    wire N__46208;
    wire N__46205;
    wire N__46202;
    wire N__46199;
    wire N__46198;
    wire N__46195;
    wire N__46192;
    wire N__46189;
    wire N__46186;
    wire N__46183;
    wire N__46180;
    wire N__46173;
    wire N__46172;
    wire N__46169;
    wire N__46166;
    wire N__46163;
    wire N__46160;
    wire N__46159;
    wire N__46154;
    wire N__46151;
    wire N__46148;
    wire N__46145;
    wire N__46142;
    wire N__46137;
    wire N__46134;
    wire N__46131;
    wire N__46128;
    wire N__46125;
    wire N__46122;
    wire N__46119;
    wire N__46116;
    wire N__46115;
    wire N__46112;
    wire N__46109;
    wire N__46106;
    wire N__46101;
    wire N__46098;
    wire N__46095;
    wire N__46092;
    wire N__46089;
    wire N__46086;
    wire N__46083;
    wire N__46080;
    wire N__46077;
    wire N__46074;
    wire N__46071;
    wire N__46068;
    wire N__46065;
    wire N__46064;
    wire N__46061;
    wire N__46060;
    wire N__46059;
    wire N__46058;
    wire N__46057;
    wire N__46056;
    wire N__46055;
    wire N__46054;
    wire N__46053;
    wire N__46052;
    wire N__46051;
    wire N__46050;
    wire N__46047;
    wire N__46046;
    wire N__46045;
    wire N__46044;
    wire N__46043;
    wire N__46042;
    wire N__46041;
    wire N__46038;
    wire N__46035;
    wire N__46032;
    wire N__46027;
    wire N__46014;
    wire N__46013;
    wire N__46010;
    wire N__46007;
    wire N__45996;
    wire N__45993;
    wire N__45992;
    wire N__45991;
    wire N__45990;
    wire N__45989;
    wire N__45984;
    wire N__45977;
    wire N__45974;
    wire N__45967;
    wire N__45962;
    wire N__45959;
    wire N__45954;
    wire N__45949;
    wire N__45944;
    wire N__45941;
    wire N__45934;
    wire N__45931;
    wire N__45926;
    wire N__45921;
    wire N__45920;
    wire N__45919;
    wire N__45916;
    wire N__45915;
    wire N__45912;
    wire N__45909;
    wire N__45908;
    wire N__45907;
    wire N__45906;
    wire N__45905;
    wire N__45904;
    wire N__45903;
    wire N__45902;
    wire N__45899;
    wire N__45896;
    wire N__45879;
    wire N__45876;
    wire N__45875;
    wire N__45874;
    wire N__45873;
    wire N__45872;
    wire N__45871;
    wire N__45870;
    wire N__45869;
    wire N__45868;
    wire N__45867;
    wire N__45866;
    wire N__45863;
    wire N__45860;
    wire N__45857;
    wire N__45854;
    wire N__45843;
    wire N__45842;
    wire N__45839;
    wire N__45836;
    wire N__45833;
    wire N__45832;
    wire N__45831;
    wire N__45826;
    wire N__45819;
    wire N__45814;
    wire N__45811;
    wire N__45808;
    wire N__45805;
    wire N__45798;
    wire N__45795;
    wire N__45788;
    wire N__45781;
    wire N__45776;
    wire N__45773;
    wire N__45768;
    wire N__45765;
    wire N__45764;
    wire N__45763;
    wire N__45760;
    wire N__45755;
    wire N__45752;
    wire N__45749;
    wire N__45744;
    wire N__45743;
    wire N__45742;
    wire N__45739;
    wire N__45736;
    wire N__45733;
    wire N__45730;
    wire N__45727;
    wire N__45724;
    wire N__45719;
    wire N__45714;
    wire N__45711;
    wire N__45708;
    wire N__45705;
    wire N__45702;
    wire N__45699;
    wire N__45696;
    wire N__45693;
    wire N__45692;
    wire N__45691;
    wire N__45688;
    wire N__45683;
    wire N__45678;
    wire N__45675;
    wire N__45674;
    wire N__45671;
    wire N__45670;
    wire N__45667;
    wire N__45664;
    wire N__45661;
    wire N__45658;
    wire N__45651;
    wire N__45648;
    wire N__45645;
    wire N__45642;
    wire N__45639;
    wire N__45636;
    wire N__45633;
    wire N__45630;
    wire N__45627;
    wire N__45624;
    wire N__45621;
    wire N__45618;
    wire N__45617;
    wire N__45614;
    wire N__45613;
    wire N__45610;
    wire N__45605;
    wire N__45602;
    wire N__45599;
    wire N__45594;
    wire N__45591;
    wire N__45588;
    wire N__45585;
    wire N__45582;
    wire N__45579;
    wire N__45576;
    wire N__45573;
    wire N__45572;
    wire N__45571;
    wire N__45570;
    wire N__45569;
    wire N__45568;
    wire N__45567;
    wire N__45552;
    wire N__45549;
    wire N__45546;
    wire N__45543;
    wire N__45540;
    wire N__45537;
    wire N__45534;
    wire N__45531;
    wire N__45530;
    wire N__45529;
    wire N__45526;
    wire N__45523;
    wire N__45520;
    wire N__45513;
    wire N__45510;
    wire N__45507;
    wire N__45504;
    wire N__45501;
    wire N__45498;
    wire N__45495;
    wire N__45492;
    wire N__45489;
    wire N__45486;
    wire N__45485;
    wire N__45482;
    wire N__45479;
    wire N__45476;
    wire N__45473;
    wire N__45470;
    wire N__45469;
    wire N__45466;
    wire N__45465;
    wire N__45464;
    wire N__45463;
    wire N__45462;
    wire N__45461;
    wire N__45460;
    wire N__45459;
    wire N__45458;
    wire N__45457;
    wire N__45456;
    wire N__45455;
    wire N__45454;
    wire N__45453;
    wire N__45452;
    wire N__45451;
    wire N__45450;
    wire N__45449;
    wire N__45448;
    wire N__45447;
    wire N__45446;
    wire N__45445;
    wire N__45444;
    wire N__45443;
    wire N__45442;
    wire N__45441;
    wire N__45438;
    wire N__45435;
    wire N__45432;
    wire N__45429;
    wire N__45428;
    wire N__45427;
    wire N__45426;
    wire N__45423;
    wire N__45422;
    wire N__45419;
    wire N__45418;
    wire N__45417;
    wire N__45416;
    wire N__45415;
    wire N__45412;
    wire N__45411;
    wire N__45410;
    wire N__45409;
    wire N__45408;
    wire N__45407;
    wire N__45406;
    wire N__45405;
    wire N__45404;
    wire N__45403;
    wire N__45402;
    wire N__45397;
    wire N__45392;
    wire N__45391;
    wire N__45390;
    wire N__45389;
    wire N__45388;
    wire N__45385;
    wire N__45382;
    wire N__45373;
    wire N__45364;
    wire N__45361;
    wire N__45360;
    wire N__45359;
    wire N__45358;
    wire N__45357;
    wire N__45354;
    wire N__45349;
    wire N__45346;
    wire N__45341;
    wire N__45336;
    wire N__45333;
    wire N__45326;
    wire N__45319;
    wire N__45310;
    wire N__45303;
    wire N__45294;
    wire N__45285;
    wire N__45282;
    wire N__45277;
    wire N__45274;
    wire N__45271;
    wire N__45266;
    wire N__45263;
    wire N__45254;
    wire N__45251;
    wire N__45248;
    wire N__45247;
    wire N__45246;
    wire N__45245;
    wire N__45244;
    wire N__45243;
    wire N__45242;
    wire N__45241;
    wire N__45240;
    wire N__45239;
    wire N__45236;
    wire N__45233;
    wire N__45232;
    wire N__45229;
    wire N__45222;
    wire N__45205;
    wire N__45202;
    wire N__45201;
    wire N__45194;
    wire N__45191;
    wire N__45182;
    wire N__45179;
    wire N__45178;
    wire N__45177;
    wire N__45176;
    wire N__45175;
    wire N__45174;
    wire N__45169;
    wire N__45162;
    wire N__45155;
    wire N__45148;
    wire N__45139;
    wire N__45136;
    wire N__45127;
    wire N__45120;
    wire N__45117;
    wire N__45114;
    wire N__45101;
    wire N__45090;
    wire N__45089;
    wire N__45088;
    wire N__45087;
    wire N__45086;
    wire N__45085;
    wire N__45084;
    wire N__45083;
    wire N__45082;
    wire N__45081;
    wire N__45080;
    wire N__45079;
    wire N__45078;
    wire N__45077;
    wire N__45076;
    wire N__45075;
    wire N__45074;
    wire N__45073;
    wire N__45072;
    wire N__45071;
    wire N__45070;
    wire N__45069;
    wire N__45068;
    wire N__45067;
    wire N__45066;
    wire N__45065;
    wire N__45064;
    wire N__45061;
    wire N__45060;
    wire N__45059;
    wire N__45058;
    wire N__45057;
    wire N__45054;
    wire N__45053;
    wire N__45052;
    wire N__45051;
    wire N__45050;
    wire N__45049;
    wire N__45048;
    wire N__45047;
    wire N__45046;
    wire N__45045;
    wire N__45044;
    wire N__45043;
    wire N__45042;
    wire N__45041;
    wire N__45040;
    wire N__45039;
    wire N__45036;
    wire N__45035;
    wire N__45034;
    wire N__45033;
    wire N__45032;
    wire N__45031;
    wire N__45030;
    wire N__45029;
    wire N__45028;
    wire N__45027;
    wire N__45026;
    wire N__45023;
    wire N__45020;
    wire N__45013;
    wire N__45010;
    wire N__44999;
    wire N__44992;
    wire N__44983;
    wire N__44974;
    wire N__44971;
    wire N__44968;
    wire N__44965;
    wire N__44964;
    wire N__44961;
    wire N__44956;
    wire N__44953;
    wire N__44950;
    wire N__44949;
    wire N__44948;
    wire N__44943;
    wire N__44936;
    wire N__44931;
    wire N__44930;
    wire N__44929;
    wire N__44926;
    wire N__44923;
    wire N__44914;
    wire N__44909;
    wire N__44906;
    wire N__44903;
    wire N__44902;
    wire N__44901;
    wire N__44900;
    wire N__44899;
    wire N__44898;
    wire N__44897;
    wire N__44896;
    wire N__44895;
    wire N__44894;
    wire N__44889;
    wire N__44882;
    wire N__44873;
    wire N__44870;
    wire N__44853;
    wire N__44850;
    wire N__44847;
    wire N__44844;
    wire N__44835;
    wire N__44832;
    wire N__44829;
    wire N__44822;
    wire N__44817;
    wire N__44804;
    wire N__44801;
    wire N__44796;
    wire N__44793;
    wire N__44788;
    wire N__44781;
    wire N__44776;
    wire N__44771;
    wire N__44766;
    wire N__44763;
    wire N__44758;
    wire N__44751;
    wire N__44746;
    wire N__44721;
    wire N__44718;
    wire N__44715;
    wire N__44712;
    wire N__44709;
    wire N__44706;
    wire N__44703;
    wire N__44700;
    wire N__44697;
    wire N__44694;
    wire N__44691;
    wire N__44688;
    wire N__44685;
    wire N__44682;
    wire N__44679;
    wire N__44676;
    wire N__44675;
    wire N__44672;
    wire N__44669;
    wire N__44666;
    wire N__44665;
    wire N__44664;
    wire N__44663;
    wire N__44662;
    wire N__44661;
    wire N__44660;
    wire N__44659;
    wire N__44658;
    wire N__44657;
    wire N__44654;
    wire N__44651;
    wire N__44648;
    wire N__44647;
    wire N__44644;
    wire N__44641;
    wire N__44640;
    wire N__44639;
    wire N__44636;
    wire N__44635;
    wire N__44632;
    wire N__44629;
    wire N__44628;
    wire N__44625;
    wire N__44624;
    wire N__44621;
    wire N__44618;
    wire N__44617;
    wire N__44616;
    wire N__44615;
    wire N__44614;
    wire N__44609;
    wire N__44606;
    wire N__44603;
    wire N__44598;
    wire N__44593;
    wire N__44592;
    wire N__44591;
    wire N__44590;
    wire N__44585;
    wire N__44582;
    wire N__44577;
    wire N__44572;
    wire N__44567;
    wire N__44564;
    wire N__44557;
    wire N__44552;
    wire N__44549;
    wire N__44548;
    wire N__44547;
    wire N__44542;
    wire N__44541;
    wire N__44538;
    wire N__44535;
    wire N__44534;
    wire N__44533;
    wire N__44530;
    wire N__44527;
    wire N__44518;
    wire N__44515;
    wire N__44510;
    wire N__44509;
    wire N__44508;
    wire N__44505;
    wire N__44500;
    wire N__44497;
    wire N__44486;
    wire N__44479;
    wire N__44474;
    wire N__44469;
    wire N__44454;
    wire N__44451;
    wire N__44448;
    wire N__44445;
    wire N__44442;
    wire N__44439;
    wire N__44436;
    wire N__44433;
    wire N__44432;
    wire N__44431;
    wire N__44428;
    wire N__44427;
    wire N__44422;
    wire N__44419;
    wire N__44418;
    wire N__44415;
    wire N__44414;
    wire N__44413;
    wire N__44410;
    wire N__44409;
    wire N__44408;
    wire N__44407;
    wire N__44406;
    wire N__44403;
    wire N__44400;
    wire N__44397;
    wire N__44394;
    wire N__44391;
    wire N__44388;
    wire N__44383;
    wire N__44378;
    wire N__44373;
    wire N__44372;
    wire N__44371;
    wire N__44370;
    wire N__44369;
    wire N__44368;
    wire N__44367;
    wire N__44360;
    wire N__44355;
    wire N__44350;
    wire N__44343;
    wire N__44340;
    wire N__44335;
    wire N__44334;
    wire N__44333;
    wire N__44332;
    wire N__44331;
    wire N__44330;
    wire N__44329;
    wire N__44328;
    wire N__44327;
    wire N__44326;
    wire N__44323;
    wire N__44320;
    wire N__44315;
    wire N__44310;
    wire N__44305;
    wire N__44300;
    wire N__44289;
    wire N__44274;
    wire N__44271;
    wire N__44268;
    wire N__44265;
    wire N__44262;
    wire N__44259;
    wire N__44256;
    wire N__44253;
    wire N__44250;
    wire N__44247;
    wire N__44244;
    wire N__44241;
    wire N__44238;
    wire N__44235;
    wire N__44232;
    wire N__44229;
    wire N__44226;
    wire N__44223;
    wire N__44220;
    wire N__44217;
    wire N__44214;
    wire N__44211;
    wire N__44208;
    wire N__44205;
    wire N__44202;
    wire N__44199;
    wire N__44196;
    wire N__44193;
    wire N__44190;
    wire N__44187;
    wire N__44184;
    wire N__44181;
    wire N__44178;
    wire N__44175;
    wire N__44172;
    wire N__44169;
    wire N__44166;
    wire N__44163;
    wire N__44160;
    wire N__44157;
    wire N__44154;
    wire N__44151;
    wire N__44148;
    wire N__44145;
    wire N__44142;
    wire N__44141;
    wire N__44140;
    wire N__44135;
    wire N__44132;
    wire N__44127;
    wire N__44124;
    wire N__44121;
    wire N__44118;
    wire N__44115;
    wire N__44112;
    wire N__44109;
    wire N__44106;
    wire N__44105;
    wire N__44102;
    wire N__44099;
    wire N__44096;
    wire N__44093;
    wire N__44092;
    wire N__44089;
    wire N__44088;
    wire N__44085;
    wire N__44082;
    wire N__44079;
    wire N__44076;
    wire N__44071;
    wire N__44068;
    wire N__44065;
    wire N__44062;
    wire N__44061;
    wire N__44058;
    wire N__44055;
    wire N__44052;
    wire N__44049;
    wire N__44046;
    wire N__44043;
    wire N__44040;
    wire N__44035;
    wire N__44030;
    wire N__44025;
    wire N__44022;
    wire N__44019;
    wire N__44016;
    wire N__44013;
    wire N__44010;
    wire N__44007;
    wire N__44004;
    wire N__44003;
    wire N__44000;
    wire N__43997;
    wire N__43994;
    wire N__43991;
    wire N__43988;
    wire N__43985;
    wire N__43982;
    wire N__43979;
    wire N__43974;
    wire N__43971;
    wire N__43968;
    wire N__43965;
    wire N__43962;
    wire N__43959;
    wire N__43956;
    wire N__43955;
    wire N__43954;
    wire N__43951;
    wire N__43948;
    wire N__43945;
    wire N__43942;
    wire N__43939;
    wire N__43938;
    wire N__43933;
    wire N__43932;
    wire N__43931;
    wire N__43928;
    wire N__43925;
    wire N__43922;
    wire N__43917;
    wire N__43914;
    wire N__43905;
    wire N__43904;
    wire N__43903;
    wire N__43902;
    wire N__43901;
    wire N__43898;
    wire N__43891;
    wire N__43888;
    wire N__43887;
    wire N__43886;
    wire N__43885;
    wire N__43882;
    wire N__43879;
    wire N__43874;
    wire N__43869;
    wire N__43866;
    wire N__43857;
    wire N__43854;
    wire N__43853;
    wire N__43852;
    wire N__43849;
    wire N__43844;
    wire N__43841;
    wire N__43836;
    wire N__43833;
    wire N__43830;
    wire N__43829;
    wire N__43828;
    wire N__43825;
    wire N__43822;
    wire N__43819;
    wire N__43814;
    wire N__43813;
    wire N__43810;
    wire N__43807;
    wire N__43804;
    wire N__43799;
    wire N__43794;
    wire N__43791;
    wire N__43790;
    wire N__43789;
    wire N__43786;
    wire N__43781;
    wire N__43778;
    wire N__43773;
    wire N__43770;
    wire N__43767;
    wire N__43764;
    wire N__43761;
    wire N__43758;
    wire N__43755;
    wire N__43752;
    wire N__43749;
    wire N__43748;
    wire N__43747;
    wire N__43746;
    wire N__43743;
    wire N__43740;
    wire N__43739;
    wire N__43734;
    wire N__43733;
    wire N__43728;
    wire N__43725;
    wire N__43722;
    wire N__43721;
    wire N__43720;
    wire N__43717;
    wire N__43712;
    wire N__43709;
    wire N__43704;
    wire N__43701;
    wire N__43698;
    wire N__43695;
    wire N__43686;
    wire N__43683;
    wire N__43680;
    wire N__43677;
    wire N__43674;
    wire N__43671;
    wire N__43670;
    wire N__43669;
    wire N__43666;
    wire N__43665;
    wire N__43664;
    wire N__43659;
    wire N__43656;
    wire N__43651;
    wire N__43648;
    wire N__43645;
    wire N__43638;
    wire N__43635;
    wire N__43632;
    wire N__43629;
    wire N__43626;
    wire N__43623;
    wire N__43620;
    wire N__43619;
    wire N__43616;
    wire N__43613;
    wire N__43612;
    wire N__43609;
    wire N__43606;
    wire N__43603;
    wire N__43600;
    wire N__43597;
    wire N__43594;
    wire N__43587;
    wire N__43584;
    wire N__43583;
    wire N__43582;
    wire N__43581;
    wire N__43580;
    wire N__43579;
    wire N__43578;
    wire N__43577;
    wire N__43576;
    wire N__43575;
    wire N__43574;
    wire N__43573;
    wire N__43572;
    wire N__43571;
    wire N__43570;
    wire N__43569;
    wire N__43566;
    wire N__43563;
    wire N__43562;
    wire N__43561;
    wire N__43560;
    wire N__43559;
    wire N__43556;
    wire N__43553;
    wire N__43550;
    wire N__43549;
    wire N__43546;
    wire N__43545;
    wire N__43542;
    wire N__43541;
    wire N__43540;
    wire N__43537;
    wire N__43534;
    wire N__43533;
    wire N__43530;
    wire N__43529;
    wire N__43526;
    wire N__43523;
    wire N__43520;
    wire N__43519;
    wire N__43518;
    wire N__43515;
    wire N__43514;
    wire N__43513;
    wire N__43512;
    wire N__43511;
    wire N__43508;
    wire N__43505;
    wire N__43502;
    wire N__43499;
    wire N__43496;
    wire N__43493;
    wire N__43492;
    wire N__43491;
    wire N__43488;
    wire N__43487;
    wire N__43484;
    wire N__43481;
    wire N__43478;
    wire N__43463;
    wire N__43460;
    wire N__43455;
    wire N__43452;
    wire N__43437;
    wire N__43436;
    wire N__43435;
    wire N__43432;
    wire N__43431;
    wire N__43428;
    wire N__43423;
    wire N__43420;
    wire N__43417;
    wire N__43412;
    wire N__43397;
    wire N__43392;
    wire N__43389;
    wire N__43384;
    wire N__43381;
    wire N__43378;
    wire N__43371;
    wire N__43370;
    wire N__43367;
    wire N__43366;
    wire N__43365;
    wire N__43362;
    wire N__43359;
    wire N__43356;
    wire N__43351;
    wire N__43342;
    wire N__43335;
    wire N__43330;
    wire N__43325;
    wire N__43322;
    wire N__43315;
    wire N__43310;
    wire N__43299;
    wire N__43296;
    wire N__43293;
    wire N__43290;
    wire N__43287;
    wire N__43284;
    wire N__43281;
    wire N__43278;
    wire N__43275;
    wire N__43272;
    wire N__43269;
    wire N__43268;
    wire N__43265;
    wire N__43262;
    wire N__43257;
    wire N__43254;
    wire N__43251;
    wire N__43248;
    wire N__43245;
    wire N__43242;
    wire N__43239;
    wire N__43236;
    wire N__43235;
    wire N__43232;
    wire N__43229;
    wire N__43224;
    wire N__43221;
    wire N__43218;
    wire N__43215;
    wire N__43212;
    wire N__43209;
    wire N__43206;
    wire N__43205;
    wire N__43202;
    wire N__43199;
    wire N__43196;
    wire N__43193;
    wire N__43188;
    wire N__43185;
    wire N__43182;
    wire N__43179;
    wire N__43176;
    wire N__43173;
    wire N__43170;
    wire N__43167;
    wire N__43164;
    wire N__43161;
    wire N__43158;
    wire N__43155;
    wire N__43152;
    wire N__43149;
    wire N__43146;
    wire N__43143;
    wire N__43142;
    wire N__43139;
    wire N__43136;
    wire N__43135;
    wire N__43134;
    wire N__43131;
    wire N__43124;
    wire N__43119;
    wire N__43116;
    wire N__43113;
    wire N__43110;
    wire N__43107;
    wire N__43104;
    wire N__43101;
    wire N__43098;
    wire N__43095;
    wire N__43092;
    wire N__43089;
    wire N__43086;
    wire N__43083;
    wire N__43080;
    wire N__43077;
    wire N__43074;
    wire N__43071;
    wire N__43068;
    wire N__43065;
    wire N__43062;
    wire N__43059;
    wire N__43056;
    wire N__43053;
    wire N__43050;
    wire N__43047;
    wire N__43044;
    wire N__43041;
    wire N__43038;
    wire N__43035;
    wire N__43034;
    wire N__43031;
    wire N__43028;
    wire N__43023;
    wire N__43020;
    wire N__43017;
    wire N__43014;
    wire N__43011;
    wire N__43008;
    wire N__43005;
    wire N__43004;
    wire N__43003;
    wire N__43000;
    wire N__42997;
    wire N__42994;
    wire N__42991;
    wire N__42986;
    wire N__42983;
    wire N__42980;
    wire N__42975;
    wire N__42972;
    wire N__42969;
    wire N__42966;
    wire N__42965;
    wire N__42964;
    wire N__42961;
    wire N__42956;
    wire N__42951;
    wire N__42948;
    wire N__42945;
    wire N__42944;
    wire N__42941;
    wire N__42940;
    wire N__42937;
    wire N__42934;
    wire N__42931;
    wire N__42928;
    wire N__42921;
    wire N__42918;
    wire N__42915;
    wire N__42912;
    wire N__42909;
    wire N__42906;
    wire N__42905;
    wire N__42904;
    wire N__42901;
    wire N__42898;
    wire N__42895;
    wire N__42888;
    wire N__42885;
    wire N__42882;
    wire N__42879;
    wire N__42876;
    wire N__42873;
    wire N__42870;
    wire N__42867;
    wire N__42864;
    wire N__42861;
    wire N__42858;
    wire N__42855;
    wire N__42852;
    wire N__42849;
    wire N__42846;
    wire N__42843;
    wire N__42840;
    wire N__42837;
    wire N__42834;
    wire N__42831;
    wire N__42828;
    wire N__42825;
    wire N__42822;
    wire N__42819;
    wire N__42816;
    wire N__42813;
    wire N__42812;
    wire N__42809;
    wire N__42806;
    wire N__42803;
    wire N__42800;
    wire N__42797;
    wire N__42794;
    wire N__42793;
    wire N__42790;
    wire N__42787;
    wire N__42784;
    wire N__42777;
    wire N__42774;
    wire N__42771;
    wire N__42768;
    wire N__42765;
    wire N__42762;
    wire N__42759;
    wire N__42758;
    wire N__42755;
    wire N__42752;
    wire N__42751;
    wire N__42748;
    wire N__42743;
    wire N__42738;
    wire N__42735;
    wire N__42732;
    wire N__42729;
    wire N__42728;
    wire N__42725;
    wire N__42724;
    wire N__42721;
    wire N__42718;
    wire N__42715;
    wire N__42712;
    wire N__42705;
    wire N__42702;
    wire N__42701;
    wire N__42698;
    wire N__42697;
    wire N__42694;
    wire N__42691;
    wire N__42686;
    wire N__42681;
    wire N__42678;
    wire N__42675;
    wire N__42674;
    wire N__42671;
    wire N__42670;
    wire N__42667;
    wire N__42664;
    wire N__42661;
    wire N__42658;
    wire N__42655;
    wire N__42650;
    wire N__42645;
    wire N__42644;
    wire N__42643;
    wire N__42640;
    wire N__42637;
    wire N__42634;
    wire N__42629;
    wire N__42626;
    wire N__42623;
    wire N__42620;
    wire N__42617;
    wire N__42612;
    wire N__42609;
    wire N__42608;
    wire N__42605;
    wire N__42604;
    wire N__42601;
    wire N__42598;
    wire N__42593;
    wire N__42590;
    wire N__42587;
    wire N__42582;
    wire N__42579;
    wire N__42578;
    wire N__42577;
    wire N__42574;
    wire N__42569;
    wire N__42566;
    wire N__42563;
    wire N__42558;
    wire N__42555;
    wire N__42554;
    wire N__42551;
    wire N__42550;
    wire N__42547;
    wire N__42544;
    wire N__42541;
    wire N__42538;
    wire N__42531;
    wire N__42528;
    wire N__42527;
    wire N__42524;
    wire N__42521;
    wire N__42518;
    wire N__42515;
    wire N__42514;
    wire N__42511;
    wire N__42508;
    wire N__42505;
    wire N__42502;
    wire N__42497;
    wire N__42494;
    wire N__42489;
    wire N__42486;
    wire N__42483;
    wire N__42482;
    wire N__42481;
    wire N__42478;
    wire N__42475;
    wire N__42472;
    wire N__42467;
    wire N__42464;
    wire N__42461;
    wire N__42458;
    wire N__42455;
    wire N__42452;
    wire N__42447;
    wire N__42446;
    wire N__42445;
    wire N__42440;
    wire N__42437;
    wire N__42434;
    wire N__42431;
    wire N__42428;
    wire N__42423;
    wire N__42420;
    wire N__42419;
    wire N__42416;
    wire N__42413;
    wire N__42412;
    wire N__42409;
    wire N__42404;
    wire N__42399;
    wire N__42396;
    wire N__42393;
    wire N__42390;
    wire N__42387;
    wire N__42384;
    wire N__42381;
    wire N__42378;
    wire N__42375;
    wire N__42372;
    wire N__42369;
    wire N__42366;
    wire N__42363;
    wire N__42360;
    wire N__42357;
    wire N__42354;
    wire N__42351;
    wire N__42348;
    wire N__42345;
    wire N__42342;
    wire N__42339;
    wire N__42336;
    wire N__42333;
    wire N__42330;
    wire N__42327;
    wire N__42324;
    wire N__42321;
    wire N__42318;
    wire N__42315;
    wire N__42312;
    wire N__42309;
    wire N__42306;
    wire N__42303;
    wire N__42300;
    wire N__42297;
    wire N__42294;
    wire N__42291;
    wire N__42288;
    wire N__42285;
    wire N__42282;
    wire N__42279;
    wire N__42278;
    wire N__42277;
    wire N__42274;
    wire N__42269;
    wire N__42266;
    wire N__42263;
    wire N__42260;
    wire N__42257;
    wire N__42252;
    wire N__42249;
    wire N__42248;
    wire N__42247;
    wire N__42244;
    wire N__42239;
    wire N__42236;
    wire N__42233;
    wire N__42230;
    wire N__42227;
    wire N__42224;
    wire N__42221;
    wire N__42216;
    wire N__42213;
    wire N__42212;
    wire N__42209;
    wire N__42208;
    wire N__42205;
    wire N__42202;
    wire N__42199;
    wire N__42196;
    wire N__42191;
    wire N__42188;
    wire N__42185;
    wire N__42182;
    wire N__42177;
    wire N__42176;
    wire N__42175;
    wire N__42172;
    wire N__42169;
    wire N__42166;
    wire N__42163;
    wire N__42160;
    wire N__42153;
    wire N__42150;
    wire N__42147;
    wire N__42144;
    wire N__42141;
    wire N__42138;
    wire N__42135;
    wire N__42132;
    wire N__42129;
    wire N__42126;
    wire N__42123;
    wire N__42120;
    wire N__42117;
    wire N__42114;
    wire N__42111;
    wire N__42108;
    wire N__42105;
    wire N__42102;
    wire N__42099;
    wire N__42096;
    wire N__42093;
    wire N__42090;
    wire N__42087;
    wire N__42084;
    wire N__42081;
    wire N__42078;
    wire N__42075;
    wire N__42072;
    wire N__42069;
    wire N__42066;
    wire N__42063;
    wire N__42060;
    wire N__42057;
    wire N__42054;
    wire N__42051;
    wire N__42048;
    wire N__42045;
    wire N__42042;
    wire N__42039;
    wire N__42036;
    wire N__42033;
    wire N__42030;
    wire N__42027;
    wire N__42024;
    wire N__42021;
    wire N__42018;
    wire N__42015;
    wire N__42012;
    wire N__42011;
    wire N__42010;
    wire N__42007;
    wire N__42004;
    wire N__42001;
    wire N__41998;
    wire N__41993;
    wire N__41988;
    wire N__41985;
    wire N__41982;
    wire N__41979;
    wire N__41976;
    wire N__41973;
    wire N__41970;
    wire N__41967;
    wire N__41964;
    wire N__41961;
    wire N__41958;
    wire N__41955;
    wire N__41952;
    wire N__41949;
    wire N__41946;
    wire N__41943;
    wire N__41940;
    wire N__41937;
    wire N__41934;
    wire N__41931;
    wire N__41928;
    wire N__41925;
    wire N__41922;
    wire N__41919;
    wire N__41916;
    wire N__41913;
    wire N__41910;
    wire N__41907;
    wire N__41904;
    wire N__41901;
    wire N__41898;
    wire N__41895;
    wire N__41892;
    wire N__41889;
    wire N__41886;
    wire N__41883;
    wire N__41880;
    wire N__41877;
    wire N__41874;
    wire N__41871;
    wire N__41868;
    wire N__41865;
    wire N__41862;
    wire N__41859;
    wire N__41856;
    wire N__41853;
    wire N__41850;
    wire N__41847;
    wire N__41844;
    wire N__41841;
    wire N__41838;
    wire N__41835;
    wire N__41832;
    wire N__41829;
    wire N__41826;
    wire N__41823;
    wire N__41820;
    wire N__41817;
    wire N__41814;
    wire N__41811;
    wire N__41808;
    wire N__41807;
    wire N__41806;
    wire N__41803;
    wire N__41800;
    wire N__41797;
    wire N__41796;
    wire N__41791;
    wire N__41788;
    wire N__41787;
    wire N__41786;
    wire N__41783;
    wire N__41778;
    wire N__41773;
    wire N__41766;
    wire N__41763;
    wire N__41760;
    wire N__41757;
    wire N__41754;
    wire N__41753;
    wire N__41752;
    wire N__41749;
    wire N__41746;
    wire N__41743;
    wire N__41740;
    wire N__41735;
    wire N__41734;
    wire N__41733;
    wire N__41730;
    wire N__41729;
    wire N__41726;
    wire N__41723;
    wire N__41720;
    wire N__41717;
    wire N__41714;
    wire N__41703;
    wire N__41700;
    wire N__41697;
    wire N__41694;
    wire N__41691;
    wire N__41690;
    wire N__41689;
    wire N__41688;
    wire N__41685;
    wire N__41682;
    wire N__41679;
    wire N__41676;
    wire N__41671;
    wire N__41668;
    wire N__41665;
    wire N__41662;
    wire N__41659;
    wire N__41658;
    wire N__41655;
    wire N__41652;
    wire N__41649;
    wire N__41646;
    wire N__41643;
    wire N__41638;
    wire N__41635;
    wire N__41628;
    wire N__41625;
    wire N__41622;
    wire N__41619;
    wire N__41616;
    wire N__41613;
    wire N__41610;
    wire N__41609;
    wire N__41606;
    wire N__41603;
    wire N__41598;
    wire N__41595;
    wire N__41592;
    wire N__41589;
    wire N__41586;
    wire N__41583;
    wire N__41580;
    wire N__41577;
    wire N__41576;
    wire N__41575;
    wire N__41574;
    wire N__41571;
    wire N__41564;
    wire N__41563;
    wire N__41560;
    wire N__41557;
    wire N__41554;
    wire N__41551;
    wire N__41548;
    wire N__41541;
    wire N__41538;
    wire N__41535;
    wire N__41532;
    wire N__41529;
    wire N__41526;
    wire N__41523;
    wire N__41522;
    wire N__41521;
    wire N__41518;
    wire N__41517;
    wire N__41512;
    wire N__41509;
    wire N__41506;
    wire N__41503;
    wire N__41500;
    wire N__41497;
    wire N__41494;
    wire N__41487;
    wire N__41484;
    wire N__41481;
    wire N__41478;
    wire N__41475;
    wire N__41472;
    wire N__41469;
    wire N__41466;
    wire N__41463;
    wire N__41460;
    wire N__41457;
    wire N__41454;
    wire N__41451;
    wire N__41448;
    wire N__41445;
    wire N__41442;
    wire N__41439;
    wire N__41436;
    wire N__41433;
    wire N__41430;
    wire N__41427;
    wire N__41424;
    wire N__41421;
    wire N__41420;
    wire N__41417;
    wire N__41414;
    wire N__41413;
    wire N__41410;
    wire N__41407;
    wire N__41406;
    wire N__41403;
    wire N__41400;
    wire N__41397;
    wire N__41394;
    wire N__41385;
    wire N__41382;
    wire N__41379;
    wire N__41378;
    wire N__41377;
    wire N__41376;
    wire N__41375;
    wire N__41372;
    wire N__41369;
    wire N__41366;
    wire N__41363;
    wire N__41360;
    wire N__41355;
    wire N__41352;
    wire N__41349;
    wire N__41348;
    wire N__41343;
    wire N__41338;
    wire N__41335;
    wire N__41328;
    wire N__41325;
    wire N__41322;
    wire N__41319;
    wire N__41316;
    wire N__41313;
    wire N__41310;
    wire N__41307;
    wire N__41304;
    wire N__41301;
    wire N__41298;
    wire N__41295;
    wire N__41292;
    wire N__41289;
    wire N__41286;
    wire N__41283;
    wire N__41280;
    wire N__41277;
    wire N__41274;
    wire N__41271;
    wire N__41268;
    wire N__41265;
    wire N__41262;
    wire N__41259;
    wire N__41256;
    wire N__41253;
    wire N__41250;
    wire N__41247;
    wire N__41244;
    wire N__41241;
    wire N__41238;
    wire N__41235;
    wire N__41234;
    wire N__41231;
    wire N__41228;
    wire N__41225;
    wire N__41222;
    wire N__41221;
    wire N__41218;
    wire N__41215;
    wire N__41212;
    wire N__41209;
    wire N__41202;
    wire N__41201;
    wire N__41198;
    wire N__41197;
    wire N__41194;
    wire N__41191;
    wire N__41188;
    wire N__41185;
    wire N__41182;
    wire N__41179;
    wire N__41176;
    wire N__41169;
    wire N__41166;
    wire N__41163;
    wire N__41160;
    wire N__41157;
    wire N__41154;
    wire N__41151;
    wire N__41148;
    wire N__41145;
    wire N__41142;
    wire N__41139;
    wire N__41136;
    wire N__41133;
    wire N__41130;
    wire N__41127;
    wire N__41126;
    wire N__41125;
    wire N__41122;
    wire N__41119;
    wire N__41116;
    wire N__41113;
    wire N__41110;
    wire N__41107;
    wire N__41104;
    wire N__41101;
    wire N__41098;
    wire N__41093;
    wire N__41088;
    wire N__41087;
    wire N__41084;
    wire N__41083;
    wire N__41078;
    wire N__41075;
    wire N__41072;
    wire N__41067;
    wire N__41064;
    wire N__41061;
    wire N__41058;
    wire N__41055;
    wire N__41054;
    wire N__41053;
    wire N__41050;
    wire N__41047;
    wire N__41044;
    wire N__41041;
    wire N__41038;
    wire N__41035;
    wire N__41028;
    wire N__41025;
    wire N__41022;
    wire N__41021;
    wire N__41020;
    wire N__41017;
    wire N__41014;
    wire N__41011;
    wire N__41008;
    wire N__41005;
    wire N__41002;
    wire N__40997;
    wire N__40994;
    wire N__40991;
    wire N__40986;
    wire N__40985;
    wire N__40982;
    wire N__40979;
    wire N__40974;
    wire N__40973;
    wire N__40970;
    wire N__40967;
    wire N__40962;
    wire N__40961;
    wire N__40958;
    wire N__40957;
    wire N__40954;
    wire N__40949;
    wire N__40946;
    wire N__40943;
    wire N__40938;
    wire N__40935;
    wire N__40932;
    wire N__40929;
    wire N__40926;
    wire N__40923;
    wire N__40920;
    wire N__40917;
    wire N__40914;
    wire N__40911;
    wire N__40908;
    wire N__40905;
    wire N__40902;
    wire N__40899;
    wire N__40896;
    wire N__40893;
    wire N__40892;
    wire N__40889;
    wire N__40888;
    wire N__40885;
    wire N__40882;
    wire N__40879;
    wire N__40876;
    wire N__40871;
    wire N__40868;
    wire N__40865;
    wire N__40860;
    wire N__40857;
    wire N__40854;
    wire N__40851;
    wire N__40848;
    wire N__40845;
    wire N__40842;
    wire N__40839;
    wire N__40836;
    wire N__40833;
    wire N__40830;
    wire N__40827;
    wire N__40824;
    wire N__40823;
    wire N__40822;
    wire N__40819;
    wire N__40816;
    wire N__40813;
    wire N__40806;
    wire N__40803;
    wire N__40800;
    wire N__40797;
    wire N__40794;
    wire N__40791;
    wire N__40788;
    wire N__40785;
    wire N__40782;
    wire N__40779;
    wire N__40776;
    wire N__40773;
    wire N__40770;
    wire N__40767;
    wire N__40766;
    wire N__40763;
    wire N__40760;
    wire N__40759;
    wire N__40754;
    wire N__40751;
    wire N__40748;
    wire N__40745;
    wire N__40742;
    wire N__40739;
    wire N__40736;
    wire N__40731;
    wire N__40728;
    wire N__40725;
    wire N__40722;
    wire N__40721;
    wire N__40718;
    wire N__40717;
    wire N__40714;
    wire N__40711;
    wire N__40708;
    wire N__40705;
    wire N__40698;
    wire N__40697;
    wire N__40696;
    wire N__40693;
    wire N__40690;
    wire N__40687;
    wire N__40684;
    wire N__40681;
    wire N__40678;
    wire N__40675;
    wire N__40672;
    wire N__40669;
    wire N__40666;
    wire N__40663;
    wire N__40660;
    wire N__40653;
    wire N__40650;
    wire N__40647;
    wire N__40644;
    wire N__40641;
    wire N__40638;
    wire N__40635;
    wire N__40632;
    wire N__40629;
    wire N__40626;
    wire N__40623;
    wire N__40620;
    wire N__40617;
    wire N__40614;
    wire N__40611;
    wire N__40608;
    wire N__40605;
    wire N__40602;
    wire N__40599;
    wire N__40596;
    wire N__40593;
    wire N__40590;
    wire N__40587;
    wire N__40584;
    wire N__40581;
    wire N__40578;
    wire N__40575;
    wire N__40572;
    wire N__40569;
    wire N__40566;
    wire N__40563;
    wire N__40560;
    wire N__40557;
    wire N__40554;
    wire N__40551;
    wire N__40548;
    wire N__40545;
    wire N__40544;
    wire N__40543;
    wire N__40540;
    wire N__40535;
    wire N__40530;
    wire N__40529;
    wire N__40526;
    wire N__40523;
    wire N__40520;
    wire N__40517;
    wire N__40514;
    wire N__40511;
    wire N__40510;
    wire N__40507;
    wire N__40504;
    wire N__40501;
    wire N__40498;
    wire N__40491;
    wire N__40488;
    wire N__40485;
    wire N__40482;
    wire N__40479;
    wire N__40476;
    wire N__40473;
    wire N__40470;
    wire N__40467;
    wire N__40464;
    wire N__40461;
    wire N__40458;
    wire N__40455;
    wire N__40452;
    wire N__40449;
    wire N__40446;
    wire N__40443;
    wire N__40440;
    wire N__40437;
    wire N__40434;
    wire N__40431;
    wire N__40428;
    wire N__40425;
    wire N__40422;
    wire N__40419;
    wire N__40416;
    wire N__40413;
    wire N__40410;
    wire N__40407;
    wire N__40404;
    wire N__40401;
    wire N__40398;
    wire N__40395;
    wire N__40392;
    wire N__40389;
    wire N__40386;
    wire N__40383;
    wire N__40380;
    wire N__40377;
    wire N__40374;
    wire N__40371;
    wire N__40368;
    wire N__40365;
    wire N__40362;
    wire N__40359;
    wire N__40356;
    wire N__40353;
    wire N__40350;
    wire N__40347;
    wire N__40344;
    wire N__40341;
    wire N__40338;
    wire N__40335;
    wire N__40332;
    wire N__40329;
    wire N__40326;
    wire N__40323;
    wire N__40320;
    wire N__40317;
    wire N__40314;
    wire N__40311;
    wire N__40308;
    wire N__40305;
    wire N__40302;
    wire N__40299;
    wire N__40296;
    wire N__40293;
    wire N__40290;
    wire N__40287;
    wire N__40284;
    wire N__40281;
    wire N__40278;
    wire N__40275;
    wire N__40272;
    wire N__40269;
    wire N__40266;
    wire N__40263;
    wire N__40260;
    wire N__40257;
    wire N__40254;
    wire N__40251;
    wire N__40248;
    wire N__40245;
    wire N__40242;
    wire N__40239;
    wire N__40236;
    wire N__40233;
    wire N__40230;
    wire N__40227;
    wire N__40224;
    wire N__40221;
    wire N__40218;
    wire N__40215;
    wire N__40212;
    wire N__40209;
    wire N__40206;
    wire N__40203;
    wire N__40200;
    wire N__40197;
    wire N__40194;
    wire N__40191;
    wire N__40188;
    wire N__40185;
    wire N__40182;
    wire N__40179;
    wire N__40176;
    wire N__40173;
    wire N__40170;
    wire N__40167;
    wire N__40164;
    wire N__40161;
    wire N__40158;
    wire N__40155;
    wire N__40152;
    wire N__40149;
    wire N__40146;
    wire N__40143;
    wire N__40140;
    wire N__40137;
    wire N__40134;
    wire N__40131;
    wire N__40128;
    wire N__40125;
    wire N__40122;
    wire N__40119;
    wire N__40116;
    wire N__40113;
    wire N__40112;
    wire N__40111;
    wire N__40108;
    wire N__40105;
    wire N__40102;
    wire N__40099;
    wire N__40098;
    wire N__40097;
    wire N__40096;
    wire N__40093;
    wire N__40090;
    wire N__40087;
    wire N__40080;
    wire N__40077;
    wire N__40074;
    wire N__40069;
    wire N__40064;
    wire N__40061;
    wire N__40060;
    wire N__40059;
    wire N__40056;
    wire N__40053;
    wire N__40048;
    wire N__40041;
    wire N__40038;
    wire N__40037;
    wire N__40034;
    wire N__40033;
    wire N__40030;
    wire N__40027;
    wire N__40024;
    wire N__40021;
    wire N__40018;
    wire N__40015;
    wire N__40012;
    wire N__40009;
    wire N__40002;
    wire N__40001;
    wire N__40000;
    wire N__39997;
    wire N__39994;
    wire N__39991;
    wire N__39988;
    wire N__39985;
    wire N__39982;
    wire N__39979;
    wire N__39976;
    wire N__39971;
    wire N__39966;
    wire N__39963;
    wire N__39960;
    wire N__39957;
    wire N__39954;
    wire N__39951;
    wire N__39948;
    wire N__39945;
    wire N__39942;
    wire N__39939;
    wire N__39936;
    wire N__39933;
    wire N__39930;
    wire N__39927;
    wire N__39924;
    wire N__39921;
    wire N__39918;
    wire N__39915;
    wire N__39912;
    wire N__39909;
    wire N__39908;
    wire N__39905;
    wire N__39902;
    wire N__39897;
    wire N__39894;
    wire N__39893;
    wire N__39890;
    wire N__39887;
    wire N__39882;
    wire N__39879;
    wire N__39878;
    wire N__39875;
    wire N__39872;
    wire N__39867;
    wire N__39864;
    wire N__39863;
    wire N__39860;
    wire N__39857;
    wire N__39852;
    wire N__39849;
    wire N__39848;
    wire N__39845;
    wire N__39842;
    wire N__39837;
    wire N__39834;
    wire N__39833;
    wire N__39830;
    wire N__39827;
    wire N__39824;
    wire N__39819;
    wire N__39816;
    wire N__39815;
    wire N__39814;
    wire N__39813;
    wire N__39812;
    wire N__39811;
    wire N__39810;
    wire N__39809;
    wire N__39800;
    wire N__39799;
    wire N__39798;
    wire N__39797;
    wire N__39796;
    wire N__39795;
    wire N__39794;
    wire N__39793;
    wire N__39792;
    wire N__39791;
    wire N__39782;
    wire N__39779;
    wire N__39770;
    wire N__39761;
    wire N__39758;
    wire N__39757;
    wire N__39754;
    wire N__39747;
    wire N__39744;
    wire N__39743;
    wire N__39742;
    wire N__39739;
    wire N__39736;
    wire N__39733;
    wire N__39730;
    wire N__39725;
    wire N__39714;
    wire N__39711;
    wire N__39710;
    wire N__39707;
    wire N__39704;
    wire N__39701;
    wire N__39696;
    wire N__39695;
    wire N__39692;
    wire N__39689;
    wire N__39686;
    wire N__39683;
    wire N__39680;
    wire N__39677;
    wire N__39674;
    wire N__39671;
    wire N__39666;
    wire N__39663;
    wire N__39660;
    wire N__39657;
    wire N__39654;
    wire N__39653;
    wire N__39650;
    wire N__39647;
    wire N__39646;
    wire N__39643;
    wire N__39640;
    wire N__39637;
    wire N__39634;
    wire N__39631;
    wire N__39624;
    wire N__39621;
    wire N__39618;
    wire N__39617;
    wire N__39614;
    wire N__39613;
    wire N__39612;
    wire N__39611;
    wire N__39608;
    wire N__39605;
    wire N__39596;
    wire N__39595;
    wire N__39590;
    wire N__39587;
    wire N__39584;
    wire N__39579;
    wire N__39576;
    wire N__39573;
    wire N__39570;
    wire N__39567;
    wire N__39566;
    wire N__39565;
    wire N__39564;
    wire N__39561;
    wire N__39558;
    wire N__39555;
    wire N__39552;
    wire N__39547;
    wire N__39540;
    wire N__39537;
    wire N__39536;
    wire N__39535;
    wire N__39532;
    wire N__39529;
    wire N__39526;
    wire N__39521;
    wire N__39516;
    wire N__39513;
    wire N__39512;
    wire N__39509;
    wire N__39506;
    wire N__39505;
    wire N__39500;
    wire N__39497;
    wire N__39494;
    wire N__39489;
    wire N__39486;
    wire N__39485;
    wire N__39482;
    wire N__39479;
    wire N__39476;
    wire N__39475;
    wire N__39470;
    wire N__39467;
    wire N__39464;
    wire N__39459;
    wire N__39456;
    wire N__39455;
    wire N__39452;
    wire N__39449;
    wire N__39448;
    wire N__39445;
    wire N__39442;
    wire N__39439;
    wire N__39434;
    wire N__39429;
    wire N__39426;
    wire N__39425;
    wire N__39422;
    wire N__39421;
    wire N__39418;
    wire N__39415;
    wire N__39412;
    wire N__39405;
    wire N__39402;
    wire N__39401;
    wire N__39400;
    wire N__39397;
    wire N__39396;
    wire N__39393;
    wire N__39392;
    wire N__39389;
    wire N__39386;
    wire N__39383;
    wire N__39382;
    wire N__39381;
    wire N__39378;
    wire N__39375;
    wire N__39374;
    wire N__39373;
    wire N__39366;
    wire N__39363;
    wire N__39362;
    wire N__39359;
    wire N__39354;
    wire N__39351;
    wire N__39350;
    wire N__39347;
    wire N__39346;
    wire N__39345;
    wire N__39340;
    wire N__39337;
    wire N__39336;
    wire N__39329;
    wire N__39326;
    wire N__39325;
    wire N__39322;
    wire N__39319;
    wire N__39316;
    wire N__39315;
    wire N__39314;
    wire N__39309;
    wire N__39306;
    wire N__39305;
    wire N__39300;
    wire N__39297;
    wire N__39296;
    wire N__39293;
    wire N__39290;
    wire N__39287;
    wire N__39286;
    wire N__39283;
    wire N__39282;
    wire N__39281;
    wire N__39278;
    wire N__39273;
    wire N__39270;
    wire N__39265;
    wire N__39262;
    wire N__39259;
    wire N__39254;
    wire N__39253;
    wire N__39244;
    wire N__39241;
    wire N__39236;
    wire N__39231;
    wire N__39226;
    wire N__39223;
    wire N__39220;
    wire N__39217;
    wire N__39212;
    wire N__39207;
    wire N__39204;
    wire N__39199;
    wire N__39196;
    wire N__39193;
    wire N__39186;
    wire N__39183;
    wire N__39180;
    wire N__39177;
    wire N__39174;
    wire N__39171;
    wire N__39168;
    wire N__39165;
    wire N__39162;
    wire N__39159;
    wire N__39156;
    wire N__39153;
    wire N__39150;
    wire N__39147;
    wire N__39146;
    wire N__39145;
    wire N__39144;
    wire N__39143;
    wire N__39142;
    wire N__39141;
    wire N__39140;
    wire N__39137;
    wire N__39134;
    wire N__39133;
    wire N__39132;
    wire N__39125;
    wire N__39120;
    wire N__39117;
    wire N__39116;
    wire N__39115;
    wire N__39114;
    wire N__39113;
    wire N__39110;
    wire N__39109;
    wire N__39108;
    wire N__39107;
    wire N__39106;
    wire N__39105;
    wire N__39102;
    wire N__39099;
    wire N__39096;
    wire N__39093;
    wire N__39088;
    wire N__39079;
    wire N__39076;
    wire N__39073;
    wire N__39064;
    wire N__39059;
    wire N__39042;
    wire N__39039;
    wire N__39036;
    wire N__39033;
    wire N__39032;
    wire N__39029;
    wire N__39026;
    wire N__39023;
    wire N__39018;
    wire N__39015;
    wire N__39012;
    wire N__39011;
    wire N__39008;
    wire N__39005;
    wire N__39002;
    wire N__38999;
    wire N__38994;
    wire N__38991;
    wire N__38988;
    wire N__38985;
    wire N__38982;
    wire N__38979;
    wire N__38976;
    wire N__38973;
    wire N__38970;
    wire N__38967;
    wire N__38964;
    wire N__38961;
    wire N__38960;
    wire N__38957;
    wire N__38954;
    wire N__38949;
    wire N__38946;
    wire N__38943;
    wire N__38940;
    wire N__38937;
    wire N__38934;
    wire N__38931;
    wire N__38928;
    wire N__38925;
    wire N__38922;
    wire N__38919;
    wire N__38916;
    wire N__38913;
    wire N__38912;
    wire N__38909;
    wire N__38906;
    wire N__38905;
    wire N__38904;
    wire N__38903;
    wire N__38900;
    wire N__38897;
    wire N__38894;
    wire N__38893;
    wire N__38892;
    wire N__38891;
    wire N__38886;
    wire N__38881;
    wire N__38878;
    wire N__38873;
    wire N__38870;
    wire N__38867;
    wire N__38862;
    wire N__38859;
    wire N__38856;
    wire N__38851;
    wire N__38848;
    wire N__38845;
    wire N__38842;
    wire N__38835;
    wire N__38832;
    wire N__38829;
    wire N__38826;
    wire N__38823;
    wire N__38822;
    wire N__38821;
    wire N__38820;
    wire N__38817;
    wire N__38814;
    wire N__38809;
    wire N__38808;
    wire N__38807;
    wire N__38806;
    wire N__38803;
    wire N__38802;
    wire N__38799;
    wire N__38796;
    wire N__38791;
    wire N__38788;
    wire N__38785;
    wire N__38782;
    wire N__38779;
    wire N__38774;
    wire N__38771;
    wire N__38766;
    wire N__38763;
    wire N__38760;
    wire N__38757;
    wire N__38754;
    wire N__38751;
    wire N__38742;
    wire N__38739;
    wire N__38736;
    wire N__38733;
    wire N__38730;
    wire N__38727;
    wire N__38726;
    wire N__38723;
    wire N__38720;
    wire N__38715;
    wire N__38712;
    wire N__38709;
    wire N__38706;
    wire N__38703;
    wire N__38700;
    wire N__38699;
    wire N__38696;
    wire N__38693;
    wire N__38690;
    wire N__38687;
    wire N__38682;
    wire N__38679;
    wire N__38676;
    wire N__38675;
    wire N__38674;
    wire N__38673;
    wire N__38670;
    wire N__38667;
    wire N__38666;
    wire N__38665;
    wire N__38664;
    wire N__38661;
    wire N__38658;
    wire N__38657;
    wire N__38656;
    wire N__38653;
    wire N__38650;
    wire N__38643;
    wire N__38638;
    wire N__38637;
    wire N__38634;
    wire N__38631;
    wire N__38626;
    wire N__38621;
    wire N__38618;
    wire N__38607;
    wire N__38604;
    wire N__38601;
    wire N__38598;
    wire N__38597;
    wire N__38596;
    wire N__38593;
    wire N__38588;
    wire N__38583;
    wire N__38580;
    wire N__38577;
    wire N__38576;
    wire N__38573;
    wire N__38570;
    wire N__38567;
    wire N__38566;
    wire N__38561;
    wire N__38558;
    wire N__38555;
    wire N__38550;
    wire N__38547;
    wire N__38544;
    wire N__38541;
    wire N__38538;
    wire N__38535;
    wire N__38532;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38520;
    wire N__38519;
    wire N__38518;
    wire N__38515;
    wire N__38510;
    wire N__38505;
    wire N__38502;
    wire N__38499;
    wire N__38496;
    wire N__38493;
    wire N__38490;
    wire N__38487;
    wire N__38484;
    wire N__38481;
    wire N__38480;
    wire N__38479;
    wire N__38476;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38461;
    wire N__38458;
    wire N__38455;
    wire N__38452;
    wire N__38445;
    wire N__38442;
    wire N__38439;
    wire N__38436;
    wire N__38433;
    wire N__38430;
    wire N__38429;
    wire N__38426;
    wire N__38425;
    wire N__38422;
    wire N__38419;
    wire N__38416;
    wire N__38413;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38394;
    wire N__38391;
    wire N__38388;
    wire N__38385;
    wire N__38382;
    wire N__38379;
    wire N__38376;
    wire N__38375;
    wire N__38374;
    wire N__38373;
    wire N__38372;
    wire N__38369;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38357;
    wire N__38352;
    wire N__38347;
    wire N__38344;
    wire N__38339;
    wire N__38336;
    wire N__38333;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38319;
    wire N__38318;
    wire N__38317;
    wire N__38316;
    wire N__38315;
    wire N__38312;
    wire N__38311;
    wire N__38308;
    wire N__38305;
    wire N__38304;
    wire N__38303;
    wire N__38302;
    wire N__38301;
    wire N__38298;
    wire N__38295;
    wire N__38292;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38278;
    wire N__38277;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38269;
    wire N__38268;
    wire N__38263;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38243;
    wire N__38240;
    wire N__38239;
    wire N__38238;
    wire N__38237;
    wire N__38234;
    wire N__38231;
    wire N__38228;
    wire N__38223;
    wire N__38222;
    wire N__38221;
    wire N__38220;
    wire N__38219;
    wire N__38218;
    wire N__38217;
    wire N__38216;
    wire N__38215;
    wire N__38214;
    wire N__38213;
    wire N__38212;
    wire N__38211;
    wire N__38208;
    wire N__38203;
    wire N__38196;
    wire N__38189;
    wire N__38184;
    wire N__38179;
    wire N__38176;
    wire N__38161;
    wire N__38152;
    wire N__38147;
    wire N__38138;
    wire N__38127;
    wire N__38124;
    wire N__38121;
    wire N__38118;
    wire N__38115;
    wire N__38112;
    wire N__38109;
    wire N__38106;
    wire N__38103;
    wire N__38100;
    wire N__38097;
    wire N__38094;
    wire N__38091;
    wire N__38088;
    wire N__38085;
    wire N__38082;
    wire N__38079;
    wire N__38078;
    wire N__38077;
    wire N__38074;
    wire N__38071;
    wire N__38068;
    wire N__38065;
    wire N__38062;
    wire N__38059;
    wire N__38056;
    wire N__38053;
    wire N__38050;
    wire N__38047;
    wire N__38044;
    wire N__38041;
    wire N__38034;
    wire N__38031;
    wire N__38028;
    wire N__38025;
    wire N__38022;
    wire N__38019;
    wire N__38016;
    wire N__38013;
    wire N__38010;
    wire N__38007;
    wire N__38004;
    wire N__38001;
    wire N__37998;
    wire N__37995;
    wire N__37992;
    wire N__37989;
    wire N__37986;
    wire N__37983;
    wire N__37980;
    wire N__37977;
    wire N__37974;
    wire N__37971;
    wire N__37968;
    wire N__37965;
    wire N__37962;
    wire N__37959;
    wire N__37956;
    wire N__37953;
    wire N__37950;
    wire N__37947;
    wire N__37944;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37934;
    wire N__37931;
    wire N__37928;
    wire N__37925;
    wire N__37922;
    wire N__37919;
    wire N__37914;
    wire N__37911;
    wire N__37908;
    wire N__37905;
    wire N__37904;
    wire N__37901;
    wire N__37898;
    wire N__37895;
    wire N__37890;
    wire N__37887;
    wire N__37884;
    wire N__37881;
    wire N__37880;
    wire N__37879;
    wire N__37878;
    wire N__37877;
    wire N__37876;
    wire N__37875;
    wire N__37874;
    wire N__37873;
    wire N__37870;
    wire N__37869;
    wire N__37868;
    wire N__37867;
    wire N__37866;
    wire N__37865;
    wire N__37864;
    wire N__37863;
    wire N__37848;
    wire N__37845;
    wire N__37844;
    wire N__37843;
    wire N__37840;
    wire N__37825;
    wire N__37824;
    wire N__37823;
    wire N__37820;
    wire N__37817;
    wire N__37814;
    wire N__37811;
    wire N__37810;
    wire N__37809;
    wire N__37808;
    wire N__37807;
    wire N__37806;
    wire N__37805;
    wire N__37804;
    wire N__37803;
    wire N__37798;
    wire N__37795;
    wire N__37792;
    wire N__37789;
    wire N__37784;
    wire N__37781;
    wire N__37768;
    wire N__37765;
    wire N__37762;
    wire N__37759;
    wire N__37754;
    wire N__37749;
    wire N__37742;
    wire N__37731;
    wire N__37728;
    wire N__37725;
    wire N__37722;
    wire N__37719;
    wire N__37716;
    wire N__37713;
    wire N__37710;
    wire N__37707;
    wire N__37706;
    wire N__37705;
    wire N__37702;
    wire N__37701;
    wire N__37700;
    wire N__37699;
    wire N__37698;
    wire N__37695;
    wire N__37694;
    wire N__37691;
    wire N__37690;
    wire N__37689;
    wire N__37688;
    wire N__37685;
    wire N__37682;
    wire N__37675;
    wire N__37672;
    wire N__37669;
    wire N__37666;
    wire N__37659;
    wire N__37658;
    wire N__37657;
    wire N__37656;
    wire N__37655;
    wire N__37654;
    wire N__37653;
    wire N__37652;
    wire N__37651;
    wire N__37650;
    wire N__37649;
    wire N__37648;
    wire N__37647;
    wire N__37646;
    wire N__37645;
    wire N__37644;
    wire N__37643;
    wire N__37642;
    wire N__37641;
    wire N__37640;
    wire N__37635;
    wire N__37632;
    wire N__37627;
    wire N__37622;
    wire N__37613;
    wire N__37604;
    wire N__37589;
    wire N__37580;
    wire N__37575;
    wire N__37570;
    wire N__37557;
    wire N__37554;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37530;
    wire N__37527;
    wire N__37524;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37485;
    wire N__37482;
    wire N__37479;
    wire N__37476;
    wire N__37473;
    wire N__37470;
    wire N__37467;
    wire N__37464;
    wire N__37461;
    wire N__37458;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37437;
    wire N__37434;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37407;
    wire N__37404;
    wire N__37401;
    wire N__37398;
    wire N__37395;
    wire N__37392;
    wire N__37389;
    wire N__37386;
    wire N__37383;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37365;
    wire N__37362;
    wire N__37359;
    wire N__37356;
    wire N__37353;
    wire N__37350;
    wire N__37347;
    wire N__37344;
    wire N__37341;
    wire N__37338;
    wire N__37335;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37302;
    wire N__37299;
    wire N__37296;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37281;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37269;
    wire N__37266;
    wire N__37263;
    wire N__37260;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37248;
    wire N__37245;
    wire N__37242;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37209;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37185;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37169;
    wire N__37168;
    wire N__37165;
    wire N__37162;
    wire N__37161;
    wire N__37160;
    wire N__37159;
    wire N__37156;
    wire N__37153;
    wire N__37150;
    wire N__37149;
    wire N__37148;
    wire N__37145;
    wire N__37140;
    wire N__37137;
    wire N__37132;
    wire N__37127;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37109;
    wire N__37108;
    wire N__37107;
    wire N__37106;
    wire N__37103;
    wire N__37100;
    wire N__37097;
    wire N__37092;
    wire N__37083;
    wire N__37082;
    wire N__37077;
    wire N__37074;
    wire N__37071;
    wire N__37068;
    wire N__37065;
    wire N__37064;
    wire N__37061;
    wire N__37058;
    wire N__37053;
    wire N__37050;
    wire N__37049;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37037;
    wire N__37032;
    wire N__37031;
    wire N__37028;
    wire N__37025;
    wire N__37020;
    wire N__37019;
    wire N__37016;
    wire N__37013;
    wire N__37008;
    wire N__37005;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36981;
    wire N__36978;
    wire N__36975;
    wire N__36972;
    wire N__36969;
    wire N__36968;
    wire N__36967;
    wire N__36964;
    wire N__36961;
    wire N__36960;
    wire N__36959;
    wire N__36958;
    wire N__36957;
    wire N__36956;
    wire N__36955;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36939;
    wire N__36934;
    wire N__36929;
    wire N__36926;
    wire N__36923;
    wire N__36918;
    wire N__36909;
    wire N__36908;
    wire N__36905;
    wire N__36904;
    wire N__36901;
    wire N__36900;
    wire N__36897;
    wire N__36894;
    wire N__36891;
    wire N__36888;
    wire N__36883;
    wire N__36880;
    wire N__36873;
    wire N__36870;
    wire N__36869;
    wire N__36868;
    wire N__36865;
    wire N__36862;
    wire N__36859;
    wire N__36856;
    wire N__36851;
    wire N__36846;
    wire N__36843;
    wire N__36840;
    wire N__36839;
    wire N__36838;
    wire N__36837;
    wire N__36836;
    wire N__36831;
    wire N__36828;
    wire N__36825;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36807;
    wire N__36804;
    wire N__36801;
    wire N__36798;
    wire N__36795;
    wire N__36792;
    wire N__36789;
    wire N__36786;
    wire N__36785;
    wire N__36780;
    wire N__36777;
    wire N__36774;
    wire N__36771;
    wire N__36770;
    wire N__36767;
    wire N__36764;
    wire N__36759;
    wire N__36756;
    wire N__36753;
    wire N__36750;
    wire N__36747;
    wire N__36744;
    wire N__36741;
    wire N__36738;
    wire N__36737;
    wire N__36736;
    wire N__36735;
    wire N__36734;
    wire N__36731;
    wire N__36722;
    wire N__36717;
    wire N__36716;
    wire N__36715;
    wire N__36714;
    wire N__36711;
    wire N__36708;
    wire N__36703;
    wire N__36696;
    wire N__36695;
    wire N__36690;
    wire N__36689;
    wire N__36686;
    wire N__36683;
    wire N__36678;
    wire N__36677;
    wire N__36676;
    wire N__36675;
    wire N__36672;
    wire N__36665;
    wire N__36662;
    wire N__36657;
    wire N__36654;
    wire N__36651;
    wire N__36648;
    wire N__36647;
    wire N__36644;
    wire N__36643;
    wire N__36642;
    wire N__36641;
    wire N__36640;
    wire N__36639;
    wire N__36638;
    wire N__36635;
    wire N__36634;
    wire N__36631;
    wire N__36626;
    wire N__36623;
    wire N__36616;
    wire N__36611;
    wire N__36600;
    wire N__36599;
    wire N__36596;
    wire N__36595;
    wire N__36592;
    wire N__36589;
    wire N__36586;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36567;
    wire N__36564;
    wire N__36561;
    wire N__36558;
    wire N__36555;
    wire N__36552;
    wire N__36549;
    wire N__36546;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36519;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36503;
    wire N__36500;
    wire N__36497;
    wire N__36494;
    wire N__36491;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36474;
    wire N__36473;
    wire N__36472;
    wire N__36469;
    wire N__36466;
    wire N__36463;
    wire N__36460;
    wire N__36453;
    wire N__36450;
    wire N__36449;
    wire N__36444;
    wire N__36441;
    wire N__36438;
    wire N__36435;
    wire N__36432;
    wire N__36431;
    wire N__36428;
    wire N__36425;
    wire N__36422;
    wire N__36417;
    wire N__36414;
    wire N__36411;
    wire N__36408;
    wire N__36405;
    wire N__36402;
    wire N__36399;
    wire N__36396;
    wire N__36393;
    wire N__36390;
    wire N__36387;
    wire N__36384;
    wire N__36381;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36369;
    wire N__36366;
    wire N__36363;
    wire N__36362;
    wire N__36359;
    wire N__36356;
    wire N__36355;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36317;
    wire N__36314;
    wire N__36311;
    wire N__36306;
    wire N__36305;
    wire N__36302;
    wire N__36299;
    wire N__36296;
    wire N__36295;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36283;
    wire N__36280;
    wire N__36273;
    wire N__36272;
    wire N__36269;
    wire N__36268;
    wire N__36265;
    wire N__36260;
    wire N__36259;
    wire N__36256;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36237;
    wire N__36236;
    wire N__36235;
    wire N__36228;
    wire N__36225;
    wire N__36222;
    wire N__36221;
    wire N__36220;
    wire N__36219;
    wire N__36218;
    wire N__36215;
    wire N__36206;
    wire N__36201;
    wire N__36198;
    wire N__36195;
    wire N__36192;
    wire N__36189;
    wire N__36186;
    wire N__36183;
    wire N__36182;
    wire N__36179;
    wire N__36176;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36159;
    wire N__36158;
    wire N__36155;
    wire N__36152;
    wire N__36147;
    wire N__36144;
    wire N__36141;
    wire N__36140;
    wire N__36137;
    wire N__36134;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36113;
    wire N__36110;
    wire N__36107;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36095;
    wire N__36092;
    wire N__36089;
    wire N__36086;
    wire N__36083;
    wire N__36080;
    wire N__36077;
    wire N__36074;
    wire N__36071;
    wire N__36068;
    wire N__36065;
    wire N__36062;
    wire N__36059;
    wire N__36056;
    wire N__36053;
    wire N__36050;
    wire N__36047;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36029;
    wire N__36026;
    wire N__36023;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36006;
    wire N__36003;
    wire N__36000;
    wire N__35997;
    wire N__35996;
    wire N__35993;
    wire N__35992;
    wire N__35991;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35987;
    wire N__35986;
    wire N__35983;
    wire N__35974;
    wire N__35973;
    wire N__35968;
    wire N__35963;
    wire N__35960;
    wire N__35957;
    wire N__35954;
    wire N__35949;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35935;
    wire N__35930;
    wire N__35925;
    wire N__35922;
    wire N__35919;
    wire N__35916;
    wire N__35915;
    wire N__35912;
    wire N__35909;
    wire N__35906;
    wire N__35903;
    wire N__35900;
    wire N__35897;
    wire N__35892;
    wire N__35889;
    wire N__35888;
    wire N__35885;
    wire N__35882;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35862;
    wire N__35861;
    wire N__35860;
    wire N__35857;
    wire N__35856;
    wire N__35855;
    wire N__35854;
    wire N__35853;
    wire N__35848;
    wire N__35845;
    wire N__35838;
    wire N__35835;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35813;
    wire N__35808;
    wire N__35803;
    wire N__35796;
    wire N__35795;
    wire N__35792;
    wire N__35789;
    wire N__35786;
    wire N__35783;
    wire N__35780;
    wire N__35777;
    wire N__35774;
    wire N__35771;
    wire N__35768;
    wire N__35763;
    wire N__35762;
    wire N__35761;
    wire N__35758;
    wire N__35757;
    wire N__35756;
    wire N__35755;
    wire N__35752;
    wire N__35749;
    wire N__35748;
    wire N__35743;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35726;
    wire N__35725;
    wire N__35724;
    wire N__35719;
    wire N__35716;
    wire N__35711;
    wire N__35708;
    wire N__35705;
    wire N__35700;
    wire N__35691;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35681;
    wire N__35680;
    wire N__35677;
    wire N__35672;
    wire N__35667;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35642;
    wire N__35639;
    wire N__35636;
    wire N__35631;
    wire N__35628;
    wire N__35625;
    wire N__35622;
    wire N__35619;
    wire N__35616;
    wire N__35613;
    wire N__35610;
    wire N__35607;
    wire N__35604;
    wire N__35603;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35580;
    wire N__35577;
    wire N__35574;
    wire N__35573;
    wire N__35570;
    wire N__35567;
    wire N__35564;
    wire N__35561;
    wire N__35558;
    wire N__35553;
    wire N__35550;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35537;
    wire N__35534;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35519;
    wire N__35516;
    wire N__35513;
    wire N__35508;
    wire N__35505;
    wire N__35502;
    wire N__35499;
    wire N__35496;
    wire N__35493;
    wire N__35490;
    wire N__35487;
    wire N__35484;
    wire N__35483;
    wire N__35482;
    wire N__35481;
    wire N__35474;
    wire N__35471;
    wire N__35468;
    wire N__35465;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35457;
    wire N__35454;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35439;
    wire N__35436;
    wire N__35433;
    wire N__35430;
    wire N__35427;
    wire N__35424;
    wire N__35421;
    wire N__35418;
    wire N__35415;
    wire N__35410;
    wire N__35407;
    wire N__35400;
    wire N__35397;
    wire N__35396;
    wire N__35395;
    wire N__35394;
    wire N__35391;
    wire N__35388;
    wire N__35383;
    wire N__35380;
    wire N__35375;
    wire N__35370;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35360;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35348;
    wire N__35343;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35331;
    wire N__35330;
    wire N__35327;
    wire N__35324;
    wire N__35321;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35307;
    wire N__35304;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35294;
    wire N__35291;
    wire N__35288;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35274;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35264;
    wire N__35261;
    wire N__35258;
    wire N__35255;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35241;
    wire N__35238;
    wire N__35235;
    wire N__35234;
    wire N__35231;
    wire N__35228;
    wire N__35225;
    wire N__35220;
    wire N__35217;
    wire N__35214;
    wire N__35211;
    wire N__35208;
    wire N__35205;
    wire N__35202;
    wire N__35199;
    wire N__35198;
    wire N__35195;
    wire N__35192;
    wire N__35189;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35177;
    wire N__35174;
    wire N__35171;
    wire N__35168;
    wire N__35163;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35130;
    wire N__35127;
    wire N__35124;
    wire N__35121;
    wire N__35118;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35106;
    wire N__35103;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35090;
    wire N__35087;
    wire N__35084;
    wire N__35079;
    wire N__35076;
    wire N__35073;
    wire N__35070;
    wire N__35067;
    wire N__35064;
    wire N__35061;
    wire N__35060;
    wire N__35057;
    wire N__35054;
    wire N__35051;
    wire N__35048;
    wire N__35045;
    wire N__35040;
    wire N__35037;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35022;
    wire N__35019;
    wire N__35018;
    wire N__35015;
    wire N__35012;
    wire N__35009;
    wire N__35004;
    wire N__35001;
    wire N__34998;
    wire N__34995;
    wire N__34992;
    wire N__34989;
    wire N__34988;
    wire N__34985;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34968;
    wire N__34965;
    wire N__34962;
    wire N__34959;
    wire N__34956;
    wire N__34953;
    wire N__34950;
    wire N__34947;
    wire N__34944;
    wire N__34943;
    wire N__34940;
    wire N__34937;
    wire N__34934;
    wire N__34931;
    wire N__34928;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34910;
    wire N__34907;
    wire N__34904;
    wire N__34901;
    wire N__34898;
    wire N__34895;
    wire N__34890;
    wire N__34887;
    wire N__34884;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34872;
    wire N__34869;
    wire N__34866;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34856;
    wire N__34853;
    wire N__34852;
    wire N__34851;
    wire N__34848;
    wire N__34845;
    wire N__34844;
    wire N__34843;
    wire N__34840;
    wire N__34837;
    wire N__34832;
    wire N__34827;
    wire N__34818;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34791;
    wire N__34788;
    wire N__34785;
    wire N__34782;
    wire N__34779;
    wire N__34776;
    wire N__34773;
    wire N__34770;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34758;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34731;
    wire N__34728;
    wire N__34725;
    wire N__34722;
    wire N__34719;
    wire N__34716;
    wire N__34713;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34701;
    wire N__34698;
    wire N__34695;
    wire N__34692;
    wire N__34689;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34677;
    wire N__34674;
    wire N__34671;
    wire N__34670;
    wire N__34667;
    wire N__34662;
    wire N__34659;
    wire N__34656;
    wire N__34655;
    wire N__34654;
    wire N__34651;
    wire N__34646;
    wire N__34641;
    wire N__34640;
    wire N__34639;
    wire N__34636;
    wire N__34633;
    wire N__34630;
    wire N__34629;
    wire N__34626;
    wire N__34621;
    wire N__34618;
    wire N__34615;
    wire N__34612;
    wire N__34609;
    wire N__34604;
    wire N__34599;
    wire N__34598;
    wire N__34597;
    wire N__34594;
    wire N__34589;
    wire N__34584;
    wire N__34581;
    wire N__34578;
    wire N__34575;
    wire N__34572;
    wire N__34569;
    wire N__34566;
    wire N__34563;
    wire N__34560;
    wire N__34557;
    wire N__34556;
    wire N__34555;
    wire N__34552;
    wire N__34551;
    wire N__34544;
    wire N__34543;
    wire N__34540;
    wire N__34537;
    wire N__34532;
    wire N__34529;
    wire N__34526;
    wire N__34521;
    wire N__34518;
    wire N__34515;
    wire N__34512;
    wire N__34511;
    wire N__34508;
    wire N__34505;
    wire N__34502;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34485;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34470;
    wire N__34467;
    wire N__34464;
    wire N__34461;
    wire N__34458;
    wire N__34457;
    wire N__34456;
    wire N__34455;
    wire N__34454;
    wire N__34453;
    wire N__34450;
    wire N__34449;
    wire N__34442;
    wire N__34433;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34421;
    wire N__34420;
    wire N__34417;
    wire N__34414;
    wire N__34411;
    wire N__34404;
    wire N__34403;
    wire N__34400;
    wire N__34397;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34382;
    wire N__34381;
    wire N__34376;
    wire N__34375;
    wire N__34372;
    wire N__34369;
    wire N__34366;
    wire N__34359;
    wire N__34358;
    wire N__34355;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34343;
    wire N__34340;
    wire N__34335;
    wire N__34334;
    wire N__34333;
    wire N__34332;
    wire N__34331;
    wire N__34330;
    wire N__34317;
    wire N__34314;
    wire N__34313;
    wire N__34310;
    wire N__34307;
    wire N__34302;
    wire N__34299;
    wire N__34296;
    wire N__34295;
    wire N__34292;
    wire N__34289;
    wire N__34286;
    wire N__34281;
    wire N__34280;
    wire N__34277;
    wire N__34276;
    wire N__34273;
    wire N__34272;
    wire N__34269;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34248;
    wire N__34245;
    wire N__34244;
    wire N__34241;
    wire N__34240;
    wire N__34237;
    wire N__34234;
    wire N__34231;
    wire N__34224;
    wire N__34221;
    wire N__34218;
    wire N__34217;
    wire N__34216;
    wire N__34213;
    wire N__34210;
    wire N__34207;
    wire N__34204;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34190;
    wire N__34189;
    wire N__34186;
    wire N__34183;
    wire N__34180;
    wire N__34173;
    wire N__34170;
    wire N__34169;
    wire N__34168;
    wire N__34167;
    wire N__34166;
    wire N__34163;
    wire N__34154;
    wire N__34149;
    wire N__34148;
    wire N__34147;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34137;
    wire N__34132;
    wire N__34129;
    wire N__34126;
    wire N__34125;
    wire N__34122;
    wire N__34117;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34102;
    wire N__34099;
    wire N__34092;
    wire N__34091;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34077;
    wire N__34074;
    wire N__34071;
    wire N__34068;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34049;
    wire N__34046;
    wire N__34043;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__34001;
    wire N__33998;
    wire N__33995;
    wire N__33994;
    wire N__33991;
    wire N__33988;
    wire N__33985;
    wire N__33980;
    wire N__33977;
    wire N__33976;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33962;
    wire N__33959;
    wire N__33956;
    wire N__33951;
    wire N__33950;
    wire N__33949;
    wire N__33948;
    wire N__33947;
    wire N__33946;
    wire N__33945;
    wire N__33944;
    wire N__33943;
    wire N__33942;
    wire N__33941;
    wire N__33940;
    wire N__33939;
    wire N__33938;
    wire N__33937;
    wire N__33936;
    wire N__33935;
    wire N__33934;
    wire N__33933;
    wire N__33932;
    wire N__33931;
    wire N__33930;
    wire N__33929;
    wire N__33926;
    wire N__33923;
    wire N__33922;
    wire N__33921;
    wire N__33920;
    wire N__33919;
    wire N__33918;
    wire N__33917;
    wire N__33916;
    wire N__33901;
    wire N__33886;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33862;
    wire N__33849;
    wire N__33846;
    wire N__33841;
    wire N__33838;
    wire N__33825;
    wire N__33822;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33783;
    wire N__33780;
    wire N__33779;
    wire N__33776;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33761;
    wire N__33758;
    wire N__33755;
    wire N__33752;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33737;
    wire N__33734;
    wire N__33731;
    wire N__33730;
    wire N__33727;
    wire N__33722;
    wire N__33717;
    wire N__33714;
    wire N__33711;
    wire N__33710;
    wire N__33707;
    wire N__33704;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33694;
    wire N__33691;
    wire N__33688;
    wire N__33683;
    wire N__33678;
    wire N__33675;
    wire N__33674;
    wire N__33673;
    wire N__33670;
    wire N__33665;
    wire N__33662;
    wire N__33659;
    wire N__33654;
    wire N__33651;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33635;
    wire N__33630;
    wire N__33627;
    wire N__33624;
    wire N__33621;
    wire N__33618;
    wire N__33615;
    wire N__33612;
    wire N__33609;
    wire N__33606;
    wire N__33603;
    wire N__33600;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33558;
    wire N__33557;
    wire N__33556;
    wire N__33553;
    wire N__33550;
    wire N__33547;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33521;
    wire N__33518;
    wire N__33515;
    wire N__33512;
    wire N__33509;
    wire N__33506;
    wire N__33501;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33489;
    wire N__33486;
    wire N__33483;
    wire N__33480;
    wire N__33479;
    wire N__33476;
    wire N__33473;
    wire N__33470;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33453;
    wire N__33450;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33431;
    wire N__33428;
    wire N__33425;
    wire N__33422;
    wire N__33419;
    wire N__33416;
    wire N__33413;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33387;
    wire N__33384;
    wire N__33381;
    wire N__33378;
    wire N__33375;
    wire N__33372;
    wire N__33369;
    wire N__33366;
    wire N__33365;
    wire N__33362;
    wire N__33359;
    wire N__33356;
    wire N__33353;
    wire N__33350;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33336;
    wire N__33333;
    wire N__33330;
    wire N__33327;
    wire N__33324;
    wire N__33321;
    wire N__33318;
    wire N__33315;
    wire N__33312;
    wire N__33309;
    wire N__33306;
    wire N__33303;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33291;
    wire N__33288;
    wire N__33285;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33270;
    wire N__33267;
    wire N__33264;
    wire N__33261;
    wire N__33258;
    wire N__33255;
    wire N__33252;
    wire N__33249;
    wire N__33246;
    wire N__33243;
    wire N__33240;
    wire N__33237;
    wire N__33234;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33207;
    wire N__33204;
    wire N__33201;
    wire N__33198;
    wire N__33195;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33183;
    wire N__33180;
    wire N__33177;
    wire N__33174;
    wire N__33171;
    wire N__33168;
    wire N__33165;
    wire N__33162;
    wire N__33159;
    wire N__33156;
    wire N__33153;
    wire N__33150;
    wire N__33147;
    wire N__33144;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33132;
    wire N__33129;
    wire N__33126;
    wire N__33123;
    wire N__33120;
    wire N__33117;
    wire N__33114;
    wire N__33111;
    wire N__33108;
    wire N__33105;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33087;
    wire N__33084;
    wire N__33081;
    wire N__33078;
    wire N__33075;
    wire N__33072;
    wire N__33069;
    wire N__33066;
    wire N__33063;
    wire N__33060;
    wire N__33057;
    wire N__33054;
    wire N__33051;
    wire N__33048;
    wire N__33045;
    wire N__33042;
    wire N__33039;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33021;
    wire N__33018;
    wire N__33015;
    wire N__33012;
    wire N__33009;
    wire N__33006;
    wire N__33003;
    wire N__33000;
    wire N__32997;
    wire N__32994;
    wire N__32993;
    wire N__32992;
    wire N__32989;
    wire N__32986;
    wire N__32983;
    wire N__32982;
    wire N__32977;
    wire N__32974;
    wire N__32973;
    wire N__32970;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32952;
    wire N__32951;
    wire N__32950;
    wire N__32949;
    wire N__32946;
    wire N__32943;
    wire N__32938;
    wire N__32931;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32907;
    wire N__32904;
    wire N__32903;
    wire N__32902;
    wire N__32901;
    wire N__32900;
    wire N__32899;
    wire N__32896;
    wire N__32885;
    wire N__32884;
    wire N__32883;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32865;
    wire N__32862;
    wire N__32859;
    wire N__32858;
    wire N__32857;
    wire N__32856;
    wire N__32855;
    wire N__32852;
    wire N__32843;
    wire N__32838;
    wire N__32835;
    wire N__32832;
    wire N__32829;
    wire N__32826;
    wire N__32825;
    wire N__32822;
    wire N__32819;
    wire N__32818;
    wire N__32817;
    wire N__32814;
    wire N__32811;
    wire N__32806;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32783;
    wire N__32782;
    wire N__32777;
    wire N__32774;
    wire N__32771;
    wire N__32770;
    wire N__32767;
    wire N__32764;
    wire N__32761;
    wire N__32758;
    wire N__32751;
    wire N__32750;
    wire N__32745;
    wire N__32744;
    wire N__32743;
    wire N__32740;
    wire N__32733;
    wire N__32730;
    wire N__32727;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32715;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32702;
    wire N__32699;
    wire N__32698;
    wire N__32697;
    wire N__32696;
    wire N__32693;
    wire N__32688;
    wire N__32685;
    wire N__32682;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32668;
    wire N__32667;
    wire N__32666;
    wire N__32661;
    wire N__32658;
    wire N__32653;
    wire N__32646;
    wire N__32643;
    wire N__32640;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32634;
    wire N__32633;
    wire N__32632;
    wire N__32631;
    wire N__32626;
    wire N__32621;
    wire N__32618;
    wire N__32613;
    wire N__32606;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32593;
    wire N__32592;
    wire N__32591;
    wire N__32588;
    wire N__32585;
    wire N__32582;
    wire N__32577;
    wire N__32568;
    wire N__32567;
    wire N__32566;
    wire N__32561;
    wire N__32558;
    wire N__32557;
    wire N__32552;
    wire N__32549;
    wire N__32546;
    wire N__32541;
    wire N__32540;
    wire N__32539;
    wire N__32538;
    wire N__32529;
    wire N__32526;
    wire N__32523;
    wire N__32520;
    wire N__32517;
    wire N__32516;
    wire N__32513;
    wire N__32512;
    wire N__32509;
    wire N__32506;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32490;
    wire N__32489;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32470;
    wire N__32465;
    wire N__32462;
    wire N__32451;
    wire N__32448;
    wire N__32445;
    wire N__32442;
    wire N__32439;
    wire N__32436;
    wire N__32433;
    wire N__32430;
    wire N__32427;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32412;
    wire N__32409;
    wire N__32406;
    wire N__32403;
    wire N__32400;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32388;
    wire N__32385;
    wire N__32382;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32363;
    wire N__32362;
    wire N__32361;
    wire N__32360;
    wire N__32357;
    wire N__32350;
    wire N__32347;
    wire N__32344;
    wire N__32341;
    wire N__32338;
    wire N__32337;
    wire N__32336;
    wire N__32331;
    wire N__32328;
    wire N__32323;
    wire N__32320;
    wire N__32313;
    wire N__32312;
    wire N__32311;
    wire N__32306;
    wire N__32303;
    wire N__32298;
    wire N__32297;
    wire N__32294;
    wire N__32291;
    wire N__32288;
    wire N__32285;
    wire N__32280;
    wire N__32277;
    wire N__32276;
    wire N__32273;
    wire N__32272;
    wire N__32271;
    wire N__32268;
    wire N__32265;
    wire N__32260;
    wire N__32257;
    wire N__32250;
    wire N__32247;
    wire N__32244;
    wire N__32241;
    wire N__32238;
    wire N__32235;
    wire N__32232;
    wire N__32229;
    wire N__32226;
    wire N__32223;
    wire N__32222;
    wire N__32219;
    wire N__32216;
    wire N__32213;
    wire N__32208;
    wire N__32207;
    wire N__32204;
    wire N__32201;
    wire N__32198;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32177;
    wire N__32172;
    wire N__32171;
    wire N__32170;
    wire N__32167;
    wire N__32164;
    wire N__32161;
    wire N__32158;
    wire N__32155;
    wire N__32152;
    wire N__32149;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32123;
    wire N__32120;
    wire N__32117;
    wire N__32114;
    wire N__32111;
    wire N__32110;
    wire N__32105;
    wire N__32102;
    wire N__32097;
    wire N__32094;
    wire N__32091;
    wire N__32088;
    wire N__32085;
    wire N__32082;
    wire N__32081;
    wire N__32080;
    wire N__32077;
    wire N__32072;
    wire N__32067;
    wire N__32064;
    wire N__32061;
    wire N__32058;
    wire N__32057;
    wire N__32052;
    wire N__32049;
    wire N__32046;
    wire N__32043;
    wire N__32040;
    wire N__32039;
    wire N__32036;
    wire N__32031;
    wire N__32028;
    wire N__32025;
    wire N__32022;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32001;
    wire N__31998;
    wire N__31995;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31985;
    wire N__31982;
    wire N__31981;
    wire N__31978;
    wire N__31975;
    wire N__31972;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31953;
    wire N__31950;
    wire N__31947;
    wire N__31944;
    wire N__31941;
    wire N__31938;
    wire N__31935;
    wire N__31932;
    wire N__31929;
    wire N__31926;
    wire N__31923;
    wire N__31920;
    wire N__31917;
    wire N__31914;
    wire N__31911;
    wire N__31908;
    wire N__31905;
    wire N__31902;
    wire N__31899;
    wire N__31896;
    wire N__31893;
    wire N__31890;
    wire N__31887;
    wire N__31884;
    wire N__31881;
    wire N__31878;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31857;
    wire N__31854;
    wire N__31851;
    wire N__31848;
    wire N__31845;
    wire N__31842;
    wire N__31839;
    wire N__31836;
    wire N__31833;
    wire N__31830;
    wire N__31827;
    wire N__31824;
    wire N__31821;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31782;
    wire N__31779;
    wire N__31776;
    wire N__31773;
    wire N__31770;
    wire N__31767;
    wire N__31764;
    wire N__31761;
    wire N__31758;
    wire N__31755;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31716;
    wire N__31713;
    wire N__31710;
    wire N__31707;
    wire N__31704;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31692;
    wire N__31689;
    wire N__31686;
    wire N__31683;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31656;
    wire N__31653;
    wire N__31650;
    wire N__31647;
    wire N__31644;
    wire N__31641;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31626;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31608;
    wire N__31605;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31589;
    wire N__31586;
    wire N__31583;
    wire N__31580;
    wire N__31575;
    wire N__31572;
    wire N__31569;
    wire N__31566;
    wire N__31563;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31548;
    wire N__31545;
    wire N__31542;
    wire N__31539;
    wire N__31536;
    wire N__31533;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31500;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31487;
    wire N__31482;
    wire N__31479;
    wire N__31478;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31458;
    wire N__31457;
    wire N__31456;
    wire N__31455;
    wire N__31452;
    wire N__31451;
    wire N__31448;
    wire N__31445;
    wire N__31442;
    wire N__31439;
    wire N__31436;
    wire N__31433;
    wire N__31430;
    wire N__31427;
    wire N__31418;
    wire N__31413;
    wire N__31410;
    wire N__31407;
    wire N__31404;
    wire N__31401;
    wire N__31398;
    wire N__31395;
    wire N__31392;
    wire N__31389;
    wire N__31386;
    wire N__31385;
    wire N__31384;
    wire N__31383;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31365;
    wire N__31364;
    wire N__31361;
    wire N__31358;
    wire N__31355;
    wire N__31350;
    wire N__31347;
    wire N__31344;
    wire N__31343;
    wire N__31340;
    wire N__31337;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31311;
    wire N__31308;
    wire N__31305;
    wire N__31302;
    wire N__31301;
    wire N__31298;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31283;
    wire N__31282;
    wire N__31281;
    wire N__31280;
    wire N__31275;
    wire N__31268;
    wire N__31263;
    wire N__31262;
    wire N__31261;
    wire N__31260;
    wire N__31259;
    wire N__31258;
    wire N__31257;
    wire N__31256;
    wire N__31255;
    wire N__31248;
    wire N__31241;
    wire N__31234;
    wire N__31227;
    wire N__31226;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31218;
    wire N__31215;
    wire N__31208;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31184;
    wire N__31181;
    wire N__31176;
    wire N__31173;
    wire N__31172;
    wire N__31171;
    wire N__31168;
    wire N__31163;
    wire N__31162;
    wire N__31161;
    wire N__31160;
    wire N__31157;
    wire N__31154;
    wire N__31147;
    wire N__31140;
    wire N__31139;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31120;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31108;
    wire N__31101;
    wire N__31098;
    wire N__31095;
    wire N__31092;
    wire N__31091;
    wire N__31090;
    wire N__31089;
    wire N__31088;
    wire N__31087;
    wire N__31086;
    wire N__31083;
    wire N__31078;
    wire N__31071;
    wire N__31068;
    wire N__31061;
    wire N__31056;
    wire N__31053;
    wire N__31052;
    wire N__31051;
    wire N__31044;
    wire N__31041;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31028;
    wire N__31027;
    wire N__31026;
    wire N__31023;
    wire N__31020;
    wire N__31017;
    wire N__31014;
    wire N__31005;
    wire N__31002;
    wire N__30999;
    wire N__30996;
    wire N__30993;
    wire N__30990;
    wire N__30989;
    wire N__30986;
    wire N__30983;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30966;
    wire N__30963;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30948;
    wire N__30945;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30909;
    wire N__30906;
    wire N__30905;
    wire N__30902;
    wire N__30899;
    wire N__30896;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30882;
    wire N__30879;
    wire N__30878;
    wire N__30875;
    wire N__30870;
    wire N__30867;
    wire N__30866;
    wire N__30863;
    wire N__30860;
    wire N__30857;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30825;
    wire N__30822;
    wire N__30819;
    wire N__30816;
    wire N__30813;
    wire N__30810;
    wire N__30807;
    wire N__30804;
    wire N__30801;
    wire N__30798;
    wire N__30795;
    wire N__30792;
    wire N__30789;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30735;
    wire N__30732;
    wire N__30729;
    wire N__30726;
    wire N__30723;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30711;
    wire N__30708;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30615;
    wire N__30612;
    wire N__30609;
    wire N__30608;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30596;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30584;
    wire N__30581;
    wire N__30576;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30561;
    wire N__30558;
    wire N__30557;
    wire N__30556;
    wire N__30555;
    wire N__30554;
    wire N__30549;
    wire N__30542;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30528;
    wire N__30525;
    wire N__30522;
    wire N__30519;
    wire N__30516;
    wire N__30515;
    wire N__30514;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30501;
    wire N__30498;
    wire N__30495;
    wire N__30492;
    wire N__30489;
    wire N__30484;
    wire N__30477;
    wire N__30476;
    wire N__30475;
    wire N__30474;
    wire N__30473;
    wire N__30472;
    wire N__30471;
    wire N__30464;
    wire N__30463;
    wire N__30462;
    wire N__30461;
    wire N__30460;
    wire N__30459;
    wire N__30458;
    wire N__30455;
    wire N__30452;
    wire N__30449;
    wire N__30446;
    wire N__30443;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30413;
    wire N__30410;
    wire N__30405;
    wire N__30402;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30381;
    wire N__30380;
    wire N__30379;
    wire N__30374;
    wire N__30371;
    wire N__30368;
    wire N__30363;
    wire N__30360;
    wire N__30357;
    wire N__30354;
    wire N__30351;
    wire N__30350;
    wire N__30349;
    wire N__30346;
    wire N__30341;
    wire N__30336;
    wire N__30335;
    wire N__30332;
    wire N__30329;
    wire N__30324;
    wire N__30323;
    wire N__30320;
    wire N__30317;
    wire N__30312;
    wire N__30311;
    wire N__30308;
    wire N__30305;
    wire N__30300;
    wire N__30299;
    wire N__30296;
    wire N__30293;
    wire N__30288;
    wire N__30285;
    wire N__30284;
    wire N__30281;
    wire N__30278;
    wire N__30273;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30259;
    wire N__30256;
    wire N__30251;
    wire N__30246;
    wire N__30243;
    wire N__30242;
    wire N__30239;
    wire N__30238;
    wire N__30235;
    wire N__30232;
    wire N__30229;
    wire N__30226;
    wire N__30219;
    wire N__30216;
    wire N__30213;
    wire N__30210;
    wire N__30207;
    wire N__30204;
    wire N__30203;
    wire N__30202;
    wire N__30195;
    wire N__30192;
    wire N__30189;
    wire N__30186;
    wire N__30183;
    wire N__30180;
    wire N__30177;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30137;
    wire N__30134;
    wire N__30131;
    wire N__30128;
    wire N__30123;
    wire N__30122;
    wire N__30121;
    wire N__30118;
    wire N__30115;
    wire N__30112;
    wire N__30109;
    wire N__30106;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30083;
    wire N__30082;
    wire N__30081;
    wire N__30078;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30068;
    wire N__30063;
    wire N__30054;
    wire N__30053;
    wire N__30052;
    wire N__30049;
    wire N__30046;
    wire N__30041;
    wire N__30036;
    wire N__30035;
    wire N__30034;
    wire N__30033;
    wire N__30030;
    wire N__30027;
    wire N__30026;
    wire N__30023;
    wire N__30020;
    wire N__30017;
    wire N__30012;
    wire N__30003;
    wire N__30000;
    wire N__29999;
    wire N__29996;
    wire N__29993;
    wire N__29988;
    wire N__29987;
    wire N__29986;
    wire N__29983;
    wire N__29976;
    wire N__29973;
    wire N__29970;
    wire N__29969;
    wire N__29968;
    wire N__29965;
    wire N__29962;
    wire N__29959;
    wire N__29958;
    wire N__29957;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29943;
    wire N__29942;
    wire N__29941;
    wire N__29940;
    wire N__29937;
    wire N__29932;
    wire N__29929;
    wire N__29924;
    wire N__29921;
    wire N__29920;
    wire N__29913;
    wire N__29910;
    wire N__29905;
    wire N__29900;
    wire N__29895;
    wire N__29892;
    wire N__29889;
    wire N__29888;
    wire N__29885;
    wire N__29882;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29868;
    wire N__29865;
    wire N__29862;
    wire N__29859;
    wire N__29856;
    wire N__29855;
    wire N__29852;
    wire N__29849;
    wire N__29846;
    wire N__29841;
    wire N__29838;
    wire N__29835;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29820;
    wire N__29817;
    wire N__29814;
    wire N__29811;
    wire N__29808;
    wire N__29805;
    wire N__29802;
    wire N__29799;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29787;
    wire N__29784;
    wire N__29781;
    wire N__29778;
    wire N__29775;
    wire N__29772;
    wire N__29769;
    wire N__29766;
    wire N__29763;
    wire N__29760;
    wire N__29757;
    wire N__29754;
    wire N__29751;
    wire N__29748;
    wire N__29745;
    wire N__29742;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29730;
    wire N__29727;
    wire N__29724;
    wire N__29721;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29694;
    wire N__29691;
    wire N__29690;
    wire N__29689;
    wire N__29686;
    wire N__29681;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29658;
    wire N__29655;
    wire N__29652;
    wire N__29649;
    wire N__29646;
    wire N__29643;
    wire N__29640;
    wire N__29637;
    wire N__29634;
    wire N__29631;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29619;
    wire N__29616;
    wire N__29613;
    wire N__29610;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29598;
    wire N__29595;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29514;
    wire N__29511;
    wire N__29508;
    wire N__29505;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29469;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29454;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29442;
    wire N__29439;
    wire N__29436;
    wire N__29433;
    wire N__29430;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29405;
    wire N__29402;
    wire N__29399;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29390;
    wire N__29389;
    wire N__29382;
    wire N__29377;
    wire N__29374;
    wire N__29367;
    wire N__29366;
    wire N__29365;
    wire N__29364;
    wire N__29363;
    wire N__29360;
    wire N__29353;
    wire N__29350;
    wire N__29347;
    wire N__29340;
    wire N__29337;
    wire N__29334;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29313;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29301;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29280;
    wire N__29277;
    wire N__29274;
    wire N__29271;
    wire N__29268;
    wire N__29265;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29250;
    wire N__29247;
    wire N__29244;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29234;
    wire N__29229;
    wire N__29226;
    wire N__29225;
    wire N__29224;
    wire N__29223;
    wire N__29222;
    wire N__29221;
    wire N__29220;
    wire N__29219;
    wire N__29216;
    wire N__29209;
    wire N__29204;
    wire N__29199;
    wire N__29190;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29178;
    wire N__29177;
    wire N__29172;
    wire N__29169;
    wire N__29168;
    wire N__29167;
    wire N__29166;
    wire N__29157;
    wire N__29154;
    wire N__29151;
    wire N__29148;
    wire N__29147;
    wire N__29146;
    wire N__29145;
    wire N__29142;
    wire N__29135;
    wire N__29130;
    wire N__29129;
    wire N__29126;
    wire N__29123;
    wire N__29118;
    wire N__29117;
    wire N__29114;
    wire N__29111;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29099;
    wire N__29096;
    wire N__29095;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29079;
    wire N__29076;
    wire N__29075;
    wire N__29074;
    wire N__29071;
    wire N__29066;
    wire N__29061;
    wire N__29060;
    wire N__29057;
    wire N__29054;
    wire N__29049;
    wire N__29048;
    wire N__29045;
    wire N__29042;
    wire N__29041;
    wire N__29038;
    wire N__29037;
    wire N__29034;
    wire N__29033;
    wire N__29030;
    wire N__29027;
    wire N__29024;
    wire N__29021;
    wire N__29016;
    wire N__29007;
    wire N__29006;
    wire N__29003;
    wire N__29000;
    wire N__28999;
    wire N__28996;
    wire N__28995;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28965;
    wire N__28962;
    wire N__28959;
    wire N__28958;
    wire N__28957;
    wire N__28956;
    wire N__28953;
    wire N__28946;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28932;
    wire N__28929;
    wire N__28926;
    wire N__28923;
    wire N__28920;
    wire N__28917;
    wire N__28914;
    wire N__28911;
    wire N__28910;
    wire N__28909;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28897;
    wire N__28890;
    wire N__28887;
    wire N__28886;
    wire N__28883;
    wire N__28880;
    wire N__28875;
    wire N__28874;
    wire N__28871;
    wire N__28868;
    wire N__28863;
    wire N__28862;
    wire N__28861;
    wire N__28858;
    wire N__28853;
    wire N__28850;
    wire N__28849;
    wire N__28848;
    wire N__28847;
    wire N__28844;
    wire N__28841;
    wire N__28834;
    wire N__28831;
    wire N__28826;
    wire N__28821;
    wire N__28820;
    wire N__28819;
    wire N__28812;
    wire N__28809;
    wire N__28806;
    wire N__28803;
    wire N__28800;
    wire N__28797;
    wire N__28796;
    wire N__28793;
    wire N__28790;
    wire N__28787;
    wire N__28782;
    wire N__28779;
    wire N__28776;
    wire N__28773;
    wire N__28770;
    wire N__28767;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28755;
    wire N__28752;
    wire N__28749;
    wire N__28746;
    wire N__28743;
    wire N__28740;
    wire N__28737;
    wire N__28734;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28722;
    wire N__28719;
    wire N__28716;
    wire N__28713;
    wire N__28710;
    wire N__28707;
    wire N__28704;
    wire N__28701;
    wire N__28698;
    wire N__28695;
    wire N__28692;
    wire N__28689;
    wire N__28686;
    wire N__28683;
    wire N__28680;
    wire N__28677;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28665;
    wire N__28662;
    wire N__28659;
    wire N__28656;
    wire N__28653;
    wire N__28650;
    wire N__28647;
    wire N__28644;
    wire N__28641;
    wire N__28638;
    wire N__28635;
    wire N__28632;
    wire N__28629;
    wire N__28626;
    wire N__28623;
    wire N__28620;
    wire N__28617;
    wire N__28614;
    wire N__28611;
    wire N__28608;
    wire N__28605;
    wire N__28602;
    wire N__28599;
    wire N__28596;
    wire N__28593;
    wire N__28590;
    wire N__28587;
    wire N__28584;
    wire N__28583;
    wire N__28580;
    wire N__28577;
    wire N__28574;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28562;
    wire N__28559;
    wire N__28556;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28542;
    wire N__28539;
    wire N__28536;
    wire N__28533;
    wire N__28530;
    wire N__28527;
    wire N__28524;
    wire N__28521;
    wire N__28518;
    wire N__28515;
    wire N__28512;
    wire N__28509;
    wire N__28506;
    wire N__28503;
    wire N__28500;
    wire N__28497;
    wire N__28494;
    wire N__28491;
    wire N__28488;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28476;
    wire N__28473;
    wire N__28470;
    wire N__28467;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28404;
    wire N__28401;
    wire N__28398;
    wire N__28395;
    wire N__28392;
    wire N__28389;
    wire N__28386;
    wire N__28383;
    wire N__28380;
    wire N__28377;
    wire N__28374;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28362;
    wire N__28359;
    wire N__28356;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28326;
    wire N__28325;
    wire N__28322;
    wire N__28321;
    wire N__28314;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28290;
    wire N__28287;
    wire N__28284;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28248;
    wire N__28245;
    wire N__28242;
    wire N__28239;
    wire N__28236;
    wire N__28233;
    wire N__28230;
    wire N__28227;
    wire N__28224;
    wire N__28221;
    wire N__28218;
    wire N__28215;
    wire N__28212;
    wire N__28209;
    wire N__28206;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28181;
    wire N__28178;
    wire N__28175;
    wire N__28174;
    wire N__28171;
    wire N__28168;
    wire N__28165;
    wire N__28162;
    wire N__28159;
    wire N__28152;
    wire N__28149;
    wire N__28146;
    wire N__28143;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28128;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28104;
    wire N__28101;
    wire N__28098;
    wire N__28095;
    wire N__28092;
    wire N__28089;
    wire N__28086;
    wire N__28083;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28047;
    wire N__28044;
    wire N__28041;
    wire N__28038;
    wire N__28035;
    wire N__28032;
    wire N__28029;
    wire N__28026;
    wire N__28023;
    wire N__28020;
    wire N__28017;
    wire N__28014;
    wire N__28011;
    wire N__28008;
    wire N__28005;
    wire N__28002;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27990;
    wire N__27987;
    wire N__27984;
    wire N__27981;
    wire N__27978;
    wire N__27977;
    wire N__27974;
    wire N__27971;
    wire N__27966;
    wire N__27965;
    wire N__27962;
    wire N__27959;
    wire N__27954;
    wire N__27951;
    wire N__27948;
    wire N__27945;
    wire N__27942;
    wire N__27939;
    wire N__27936;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27912;
    wire N__27911;
    wire N__27908;
    wire N__27905;
    wire N__27900;
    wire N__27897;
    wire N__27894;
    wire N__27891;
    wire N__27888;
    wire N__27885;
    wire N__27884;
    wire N__27881;
    wire N__27878;
    wire N__27873;
    wire N__27870;
    wire N__27869;
    wire N__27866;
    wire N__27863;
    wire N__27858;
    wire N__27855;
    wire N__27854;
    wire N__27851;
    wire N__27848;
    wire N__27845;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27827;
    wire N__27824;
    wire N__27823;
    wire N__27822;
    wire N__27821;
    wire N__27818;
    wire N__27817;
    wire N__27814;
    wire N__27803;
    wire N__27798;
    wire N__27795;
    wire N__27792;
    wire N__27789;
    wire N__27788;
    wire N__27787;
    wire N__27786;
    wire N__27785;
    wire N__27784;
    wire N__27783;
    wire N__27782;
    wire N__27781;
    wire N__27780;
    wire N__27779;
    wire N__27778;
    wire N__27777;
    wire N__27776;
    wire N__27775;
    wire N__27774;
    wire N__27773;
    wire N__27772;
    wire N__27771;
    wire N__27770;
    wire N__27769;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27745;
    wire N__27728;
    wire N__27719;
    wire N__27708;
    wire N__27707;
    wire N__27704;
    wire N__27701;
    wire N__27698;
    wire N__27695;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27665;
    wire N__27662;
    wire N__27659;
    wire N__27654;
    wire N__27653;
    wire N__27650;
    wire N__27647;
    wire N__27642;
    wire N__27639;
    wire N__27638;
    wire N__27635;
    wire N__27632;
    wire N__27627;
    wire N__27626;
    wire N__27623;
    wire N__27620;
    wire N__27615;
    wire N__27612;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27600;
    wire N__27599;
    wire N__27598;
    wire N__27597;
    wire N__27596;
    wire N__27591;
    wire N__27584;
    wire N__27579;
    wire N__27578;
    wire N__27573;
    wire N__27572;
    wire N__27569;
    wire N__27568;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27556;
    wire N__27553;
    wire N__27548;
    wire N__27545;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27504;
    wire N__27501;
    wire N__27498;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27486;
    wire N__27483;
    wire N__27480;
    wire N__27477;
    wire N__27474;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27345;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27321;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27285;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27273;
    wire N__27270;
    wire N__27267;
    wire N__27264;
    wire N__27261;
    wire N__27258;
    wire N__27255;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27240;
    wire N__27237;
    wire N__27236;
    wire N__27235;
    wire N__27232;
    wire N__27229;
    wire N__27226;
    wire N__27223;
    wire N__27220;
    wire N__27217;
    wire N__27210;
    wire N__27209;
    wire N__27208;
    wire N__27207;
    wire N__27204;
    wire N__27199;
    wire N__27196;
    wire N__27195;
    wire N__27194;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27184;
    wire N__27183;
    wire N__27182;
    wire N__27177;
    wire N__27174;
    wire N__27169;
    wire N__27166;
    wire N__27161;
    wire N__27150;
    wire N__27149;
    wire N__27148;
    wire N__27147;
    wire N__27146;
    wire N__27145;
    wire N__27144;
    wire N__27143;
    wire N__27142;
    wire N__27141;
    wire N__27140;
    wire N__27139;
    wire N__27138;
    wire N__27137;
    wire N__27136;
    wire N__27135;
    wire N__27134;
    wire N__27133;
    wire N__27132;
    wire N__27131;
    wire N__27128;
    wire N__27125;
    wire N__27114;
    wire N__27111;
    wire N__27108;
    wire N__27107;
    wire N__27098;
    wire N__27083;
    wire N__27080;
    wire N__27073;
    wire N__27070;
    wire N__27069;
    wire N__27068;
    wire N__27065;
    wire N__27060;
    wire N__27055;
    wire N__27052;
    wire N__27047;
    wire N__27036;
    wire N__27035;
    wire N__27032;
    wire N__27027;
    wire N__27024;
    wire N__27021;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27003;
    wire N__27000;
    wire N__26999;
    wire N__26998;
    wire N__26997;
    wire N__26996;
    wire N__26995;
    wire N__26994;
    wire N__26991;
    wire N__26990;
    wire N__26983;
    wire N__26982;
    wire N__26977;
    wire N__26976;
    wire N__26973;
    wire N__26970;
    wire N__26967;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26948;
    wire N__26937;
    wire N__26934;
    wire N__26933;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26924;
    wire N__26923;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26906;
    wire N__26895;
    wire N__26894;
    wire N__26893;
    wire N__26890;
    wire N__26889;
    wire N__26888;
    wire N__26883;
    wire N__26878;
    wire N__26875;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26847;
    wire N__26844;
    wire N__26841;
    wire N__26838;
    wire N__26835;
    wire N__26832;
    wire N__26829;
    wire N__26826;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26808;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26790;
    wire N__26787;
    wire N__26784;
    wire N__26781;
    wire N__26778;
    wire N__26775;
    wire N__26772;
    wire N__26769;
    wire N__26766;
    wire N__26763;
    wire N__26760;
    wire N__26757;
    wire N__26754;
    wire N__26751;
    wire N__26748;
    wire N__26745;
    wire N__26742;
    wire N__26739;
    wire N__26736;
    wire N__26733;
    wire N__26730;
    wire N__26727;
    wire N__26724;
    wire N__26721;
    wire N__26718;
    wire N__26715;
    wire N__26712;
    wire N__26709;
    wire N__26706;
    wire N__26703;
    wire N__26700;
    wire N__26697;
    wire N__26694;
    wire N__26691;
    wire N__26688;
    wire N__26685;
    wire N__26682;
    wire N__26679;
    wire N__26676;
    wire N__26673;
    wire N__26672;
    wire N__26669;
    wire N__26666;
    wire N__26665;
    wire N__26662;
    wire N__26659;
    wire N__26656;
    wire N__26655;
    wire N__26652;
    wire N__26647;
    wire N__26644;
    wire N__26637;
    wire N__26636;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26618;
    wire N__26613;
    wire N__26610;
    wire N__26607;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26595;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26580;
    wire N__26577;
    wire N__26574;
    wire N__26571;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26556;
    wire N__26553;
    wire N__26552;
    wire N__26549;
    wire N__26548;
    wire N__26545;
    wire N__26542;
    wire N__26539;
    wire N__26538;
    wire N__26535;
    wire N__26530;
    wire N__26527;
    wire N__26524;
    wire N__26519;
    wire N__26514;
    wire N__26511;
    wire N__26510;
    wire N__26509;
    wire N__26506;
    wire N__26503;
    wire N__26502;
    wire N__26499;
    wire N__26496;
    wire N__26493;
    wire N__26490;
    wire N__26487;
    wire N__26482;
    wire N__26479;
    wire N__26472;
    wire N__26469;
    wire N__26466;
    wire N__26465;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26457;
    wire N__26454;
    wire N__26451;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26437;
    wire N__26434;
    wire N__26427;
    wire N__26424;
    wire N__26421;
    wire N__26420;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26412;
    wire N__26409;
    wire N__26404;
    wire N__26401;
    wire N__26398;
    wire N__26393;
    wire N__26388;
    wire N__26385;
    wire N__26384;
    wire N__26381;
    wire N__26380;
    wire N__26377;
    wire N__26376;
    wire N__26373;
    wire N__26370;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26355;
    wire N__26352;
    wire N__26343;
    wire N__26340;
    wire N__26339;
    wire N__26338;
    wire N__26337;
    wire N__26336;
    wire N__26335;
    wire N__26334;
    wire N__26333;
    wire N__26332;
    wire N__26331;
    wire N__26330;
    wire N__26329;
    wire N__26328;
    wire N__26327;
    wire N__26326;
    wire N__26325;
    wire N__26324;
    wire N__26321;
    wire N__26320;
    wire N__26317;
    wire N__26316;
    wire N__26313;
    wire N__26312;
    wire N__26307;
    wire N__26302;
    wire N__26297;
    wire N__26296;
    wire N__26293;
    wire N__26292;
    wire N__26289;
    wire N__26288;
    wire N__26285;
    wire N__26284;
    wire N__26281;
    wire N__26278;
    wire N__26277;
    wire N__26276;
    wire N__26273;
    wire N__26272;
    wire N__26271;
    wire N__26268;
    wire N__26265;
    wire N__26264;
    wire N__26263;
    wire N__26258;
    wire N__26249;
    wire N__26246;
    wire N__26241;
    wire N__26230;
    wire N__26213;
    wire N__26202;
    wire N__26187;
    wire N__26186;
    wire N__26183;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26169;
    wire N__26166;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26152;
    wire N__26147;
    wire N__26142;
    wire N__26139;
    wire N__26136;
    wire N__26133;
    wire N__26130;
    wire N__26127;
    wire N__26124;
    wire N__26121;
    wire N__26118;
    wire N__26115;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26100;
    wire N__26097;
    wire N__26096;
    wire N__26093;
    wire N__26090;
    wire N__26087;
    wire N__26082;
    wire N__26079;
    wire N__26078;
    wire N__26075;
    wire N__26072;
    wire N__26069;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26057;
    wire N__26054;
    wire N__26051;
    wire N__26048;
    wire N__26043;
    wire N__26040;
    wire N__26039;
    wire N__26038;
    wire N__26037;
    wire N__26036;
    wire N__26029;
    wire N__26024;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26009;
    wire N__26006;
    wire N__26003;
    wire N__26000;
    wire N__25995;
    wire N__25992;
    wire N__25991;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25981;
    wire N__25978;
    wire N__25971;
    wire N__25968;
    wire N__25965;
    wire N__25962;
    wire N__25959;
    wire N__25958;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25938;
    wire N__25935;
    wire N__25932;
    wire N__25929;
    wire N__25926;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25918;
    wire N__25915;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25899;
    wire N__25896;
    wire N__25893;
    wire N__25890;
    wire N__25887;
    wire N__25884;
    wire N__25883;
    wire N__25880;
    wire N__25877;
    wire N__25874;
    wire N__25869;
    wire N__25866;
    wire N__25863;
    wire N__25860;
    wire N__25857;
    wire N__25854;
    wire N__25851;
    wire N__25848;
    wire N__25845;
    wire N__25844;
    wire N__25841;
    wire N__25840;
    wire N__25839;
    wire N__25838;
    wire N__25835;
    wire N__25832;
    wire N__25829;
    wire N__25824;
    wire N__25821;
    wire N__25812;
    wire N__25809;
    wire N__25808;
    wire N__25805;
    wire N__25804;
    wire N__25803;
    wire N__25802;
    wire N__25799;
    wire N__25796;
    wire N__25789;
    wire N__25782;
    wire N__25781;
    wire N__25780;
    wire N__25779;
    wire N__25778;
    wire N__25775;
    wire N__25766;
    wire N__25763;
    wire N__25760;
    wire N__25755;
    wire N__25752;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25743;
    wire N__25742;
    wire N__25741;
    wire N__25740;
    wire N__25737;
    wire N__25736;
    wire N__25733;
    wire N__25716;
    wire N__25711;
    wire N__25704;
    wire N__25701;
    wire N__25698;
    wire N__25697;
    wire N__25696;
    wire N__25695;
    wire N__25690;
    wire N__25687;
    wire N__25686;
    wire N__25683;
    wire N__25682;
    wire N__25681;
    wire N__25678;
    wire N__25673;
    wire N__25670;
    wire N__25665;
    wire N__25660;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25644;
    wire N__25641;
    wire N__25638;
    wire N__25635;
    wire N__25632;
    wire N__25629;
    wire N__25628;
    wire N__25627;
    wire N__25626;
    wire N__25623;
    wire N__25618;
    wire N__25617;
    wire N__25616;
    wire N__25613;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25595;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25578;
    wire N__25577;
    wire N__25574;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25554;
    wire N__25545;
    wire N__25542;
    wire N__25539;
    wire N__25536;
    wire N__25535;
    wire N__25534;
    wire N__25531;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25523;
    wire N__25520;
    wire N__25517;
    wire N__25514;
    wire N__25509;
    wire N__25506;
    wire N__25503;
    wire N__25496;
    wire N__25491;
    wire N__25488;
    wire N__25487;
    wire N__25484;
    wire N__25483;
    wire N__25480;
    wire N__25477;
    wire N__25474;
    wire N__25471;
    wire N__25468;
    wire N__25461;
    wire N__25460;
    wire N__25459;
    wire N__25458;
    wire N__25453;
    wire N__25448;
    wire N__25447;
    wire N__25444;
    wire N__25441;
    wire N__25440;
    wire N__25437;
    wire N__25432;
    wire N__25429;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25410;
    wire N__25407;
    wire N__25404;
    wire N__25401;
    wire N__25398;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25386;
    wire N__25385;
    wire N__25382;
    wire N__25379;
    wire N__25376;
    wire N__25373;
    wire N__25370;
    wire N__25367;
    wire N__25364;
    wire N__25361;
    wire N__25358;
    wire N__25355;
    wire N__25352;
    wire N__25349;
    wire N__25346;
    wire N__25343;
    wire N__25340;
    wire N__25337;
    wire N__25334;
    wire N__25331;
    wire N__25328;
    wire N__25325;
    wire N__25322;
    wire N__25319;
    wire N__25316;
    wire N__25313;
    wire N__25310;
    wire N__25307;
    wire N__25304;
    wire N__25301;
    wire N__25298;
    wire N__25295;
    wire N__25292;
    wire N__25289;
    wire N__25284;
    wire N__25283;
    wire N__25280;
    wire N__25277;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25265;
    wire N__25262;
    wire N__25259;
    wire N__25256;
    wire N__25253;
    wire N__25250;
    wire N__25247;
    wire N__25244;
    wire N__25241;
    wire N__25238;
    wire N__25235;
    wire N__25232;
    wire N__25229;
    wire N__25226;
    wire N__25223;
    wire N__25220;
    wire N__25217;
    wire N__25214;
    wire N__25211;
    wire N__25208;
    wire N__25205;
    wire N__25202;
    wire N__25199;
    wire N__25196;
    wire N__25193;
    wire N__25190;
    wire N__25187;
    wire N__25182;
    wire N__25181;
    wire N__25178;
    wire N__25175;
    wire N__25172;
    wire N__25169;
    wire N__25166;
    wire N__25163;
    wire N__25160;
    wire N__25157;
    wire N__25154;
    wire N__25151;
    wire N__25148;
    wire N__25145;
    wire N__25142;
    wire N__25139;
    wire N__25136;
    wire N__25133;
    wire N__25130;
    wire N__25127;
    wire N__25124;
    wire N__25121;
    wire N__25118;
    wire N__25115;
    wire N__25112;
    wire N__25109;
    wire N__25106;
    wire N__25103;
    wire N__25100;
    wire N__25097;
    wire N__25094;
    wire N__25091;
    wire N__25088;
    wire N__25085;
    wire N__25080;
    wire N__25077;
    wire N__25076;
    wire N__25075;
    wire N__25074;
    wire N__25071;
    wire N__25064;
    wire N__25059;
    wire N__25056;
    wire N__25053;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25041;
    wire N__25038;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25026;
    wire N__25023;
    wire N__25020;
    wire N__25017;
    wire N__25014;
    wire N__25011;
    wire N__25008;
    wire N__25005;
    wire N__25004;
    wire N__25001;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24986;
    wire N__24983;
    wire N__24980;
    wire N__24977;
    wire N__24974;
    wire N__24971;
    wire N__24968;
    wire N__24965;
    wire N__24962;
    wire N__24959;
    wire N__24956;
    wire N__24953;
    wire N__24950;
    wire N__24947;
    wire N__24944;
    wire N__24941;
    wire N__24938;
    wire N__24935;
    wire N__24932;
    wire N__24929;
    wire N__24926;
    wire N__24923;
    wire N__24920;
    wire N__24917;
    wire N__24914;
    wire N__24911;
    wire N__24908;
    wire N__24905;
    wire N__24902;
    wire N__24899;
    wire N__24896;
    wire N__24891;
    wire N__24888;
    wire N__24887;
    wire N__24884;
    wire N__24881;
    wire N__24876;
    wire N__24873;
    wire N__24870;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24858;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24836;
    wire N__24833;
    wire N__24830;
    wire N__24825;
    wire N__24822;
    wire N__24819;
    wire N__24818;
    wire N__24815;
    wire N__24812;
    wire N__24807;
    wire N__24804;
    wire N__24803;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24788;
    wire N__24785;
    wire N__24782;
    wire N__24779;
    wire N__24776;
    wire N__24773;
    wire N__24770;
    wire N__24767;
    wire N__24764;
    wire N__24761;
    wire N__24758;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24743;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24731;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24719;
    wire N__24716;
    wire N__24713;
    wire N__24710;
    wire N__24707;
    wire N__24702;
    wire N__24699;
    wire N__24698;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24683;
    wire N__24680;
    wire N__24679;
    wire N__24674;
    wire N__24671;
    wire N__24666;
    wire N__24665;
    wire N__24662;
    wire N__24661;
    wire N__24658;
    wire N__24657;
    wire N__24654;
    wire N__24651;
    wire N__24648;
    wire N__24645;
    wire N__24642;
    wire N__24639;
    wire N__24634;
    wire N__24629;
    wire N__24624;
    wire N__24621;
    wire N__24620;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24605;
    wire N__24602;
    wire N__24601;
    wire N__24596;
    wire N__24593;
    wire N__24588;
    wire N__24585;
    wire N__24584;
    wire N__24583;
    wire N__24580;
    wire N__24577;
    wire N__24574;
    wire N__24571;
    wire N__24568;
    wire N__24565;
    wire N__24564;
    wire N__24557;
    wire N__24554;
    wire N__24549;
    wire N__24548;
    wire N__24545;
    wire N__24542;
    wire N__24537;
    wire N__24534;
    wire N__24533;
    wire N__24532;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24513;
    wire N__24510;
    wire N__24505;
    wire N__24502;
    wire N__24495;
    wire N__24492;
    wire N__24491;
    wire N__24488;
    wire N__24485;
    wire N__24484;
    wire N__24483;
    wire N__24478;
    wire N__24475;
    wire N__24472;
    wire N__24467;
    wire N__24464;
    wire N__24459;
    wire N__24456;
    wire N__24453;
    wire N__24452;
    wire N__24449;
    wire N__24446;
    wire N__24445;
    wire N__24440;
    wire N__24437;
    wire N__24434;
    wire N__24431;
    wire N__24430;
    wire N__24425;
    wire N__24422;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24396;
    wire N__24393;
    wire N__24392;
    wire N__24391;
    wire N__24388;
    wire N__24387;
    wire N__24384;
    wire N__24381;
    wire N__24378;
    wire N__24375;
    wire N__24372;
    wire N__24369;
    wire N__24364;
    wire N__24359;
    wire N__24354;
    wire N__24353;
    wire N__24350;
    wire N__24349;
    wire N__24346;
    wire N__24345;
    wire N__24342;
    wire N__24339;
    wire N__24336;
    wire N__24333;
    wire N__24328;
    wire N__24323;
    wire N__24318;
    wire N__24317;
    wire N__24314;
    wire N__24311;
    wire N__24310;
    wire N__24307;
    wire N__24304;
    wire N__24301;
    wire N__24298;
    wire N__24293;
    wire N__24292;
    wire N__24287;
    wire N__24284;
    wire N__24279;
    wire N__24276;
    wire N__24275;
    wire N__24274;
    wire N__24271;
    wire N__24268;
    wire N__24265;
    wire N__24262;
    wire N__24259;
    wire N__24256;
    wire N__24255;
    wire N__24248;
    wire N__24245;
    wire N__24240;
    wire N__24239;
    wire N__24236;
    wire N__24235;
    wire N__24232;
    wire N__24231;
    wire N__24228;
    wire N__24225;
    wire N__24222;
    wire N__24219;
    wire N__24216;
    wire N__24213;
    wire N__24208;
    wire N__24203;
    wire N__24198;
    wire N__24197;
    wire N__24194;
    wire N__24193;
    wire N__24190;
    wire N__24189;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24172;
    wire N__24167;
    wire N__24164;
    wire N__24159;
    wire N__24158;
    wire N__24155;
    wire N__24154;
    wire N__24151;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24133;
    wire N__24128;
    wire N__24123;
    wire N__24120;
    wire N__24119;
    wire N__24118;
    wire N__24117;
    wire N__24114;
    wire N__24111;
    wire N__24108;
    wire N__24105;
    wire N__24102;
    wire N__24099;
    wire N__24096;
    wire N__24093;
    wire N__24090;
    wire N__24083;
    wire N__24078;
    wire N__24077;
    wire N__24074;
    wire N__24073;
    wire N__24070;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24052;
    wire N__24047;
    wire N__24042;
    wire N__24041;
    wire N__24038;
    wire N__24037;
    wire N__24034;
    wire N__24033;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24016;
    wire N__24011;
    wire N__24006;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23976;
    wire N__23967;
    wire N__23964;
    wire N__23963;
    wire N__23962;
    wire N__23961;
    wire N__23958;
    wire N__23955;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23937;
    wire N__23934;
    wire N__23927;
    wire N__23922;
    wire N__23921;
    wire N__23920;
    wire N__23917;
    wire N__23914;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23904;
    wire N__23901;
    wire N__23898;
    wire N__23895;
    wire N__23888;
    wire N__23883;
    wire N__23882;
    wire N__23879;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23861;
    wire N__23860;
    wire N__23855;
    wire N__23852;
    wire N__23847;
    wire N__23844;
    wire N__23841;
    wire N__23840;
    wire N__23837;
    wire N__23836;
    wire N__23833;
    wire N__23830;
    wire N__23827;
    wire N__23824;
    wire N__23819;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23802;
    wire N__23799;
    wire N__23798;
    wire N__23795;
    wire N__23794;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23781;
    wire N__23778;
    wire N__23773;
    wire N__23768;
    wire N__23763;
    wire N__23760;
    wire N__23757;
    wire N__23754;
    wire N__23751;
    wire N__23748;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23732;
    wire N__23729;
    wire N__23726;
    wire N__23721;
    wire N__23720;
    wire N__23717;
    wire N__23716;
    wire N__23713;
    wire N__23710;
    wire N__23707;
    wire N__23704;
    wire N__23699;
    wire N__23698;
    wire N__23693;
    wire N__23690;
    wire N__23685;
    wire N__23684;
    wire N__23681;
    wire N__23678;
    wire N__23677;
    wire N__23674;
    wire N__23671;
    wire N__23668;
    wire N__23665;
    wire N__23660;
    wire N__23659;
    wire N__23654;
    wire N__23651;
    wire N__23646;
    wire N__23643;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23631;
    wire N__23628;
    wire N__23625;
    wire N__23622;
    wire N__23621;
    wire N__23618;
    wire N__23615;
    wire N__23610;
    wire N__23607;
    wire N__23606;
    wire N__23603;
    wire N__23600;
    wire N__23597;
    wire N__23592;
    wire N__23591;
    wire N__23588;
    wire N__23587;
    wire N__23582;
    wire N__23579;
    wire N__23574;
    wire N__23573;
    wire N__23568;
    wire N__23565;
    wire N__23564;
    wire N__23563;
    wire N__23560;
    wire N__23557;
    wire N__23554;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23542;
    wire N__23539;
    wire N__23536;
    wire N__23529;
    wire N__23528;
    wire N__23527;
    wire N__23524;
    wire N__23521;
    wire N__23518;
    wire N__23515;
    wire N__23508;
    wire N__23507;
    wire N__23506;
    wire N__23503;
    wire N__23500;
    wire N__23497;
    wire N__23490;
    wire N__23487;
    wire N__23486;
    wire N__23485;
    wire N__23480;
    wire N__23477;
    wire N__23472;
    wire N__23471;
    wire N__23468;
    wire N__23463;
    wire N__23460;
    wire N__23457;
    wire N__23454;
    wire N__23451;
    wire N__23450;
    wire N__23449;
    wire N__23448;
    wire N__23447;
    wire N__23446;
    wire N__23443;
    wire N__23442;
    wire N__23441;
    wire N__23438;
    wire N__23433;
    wire N__23428;
    wire N__23425;
    wire N__23422;
    wire N__23419;
    wire N__23406;
    wire N__23405;
    wire N__23404;
    wire N__23403;
    wire N__23402;
    wire N__23395;
    wire N__23390;
    wire N__23385;
    wire N__23384;
    wire N__23383;
    wire N__23378;
    wire N__23375;
    wire N__23370;
    wire N__23367;
    wire N__23366;
    wire N__23363;
    wire N__23360;
    wire N__23357;
    wire N__23354;
    wire N__23349;
    wire N__23348;
    wire N__23347;
    wire N__23344;
    wire N__23341;
    wire N__23338;
    wire N__23331;
    wire N__23328;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23313;
    wire N__23310;
    wire N__23309;
    wire N__23304;
    wire N__23301;
    wire N__23298;
    wire N__23297;
    wire N__23292;
    wire N__23289;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23279;
    wire N__23276;
    wire N__23273;
    wire N__23268;
    wire N__23265;
    wire N__23262;
    wire N__23259;
    wire N__23256;
    wire N__23253;
    wire N__23250;
    wire N__23247;
    wire N__23244;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23229;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23211;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23196;
    wire N__23193;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23181;
    wire N__23178;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23166;
    wire N__23163;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23151;
    wire N__23148;
    wire N__23145;
    wire N__23142;
    wire N__23139;
    wire N__23136;
    wire N__23133;
    wire N__23130;
    wire N__23127;
    wire N__23124;
    wire N__23121;
    wire N__23118;
    wire N__23115;
    wire N__23112;
    wire N__23109;
    wire N__23106;
    wire N__23103;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23087;
    wire N__23084;
    wire N__23081;
    wire N__23078;
    wire N__23075;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23046;
    wire N__23043;
    wire N__23040;
    wire N__23037;
    wire N__23034;
    wire N__23031;
    wire N__23028;
    wire N__23025;
    wire N__23022;
    wire N__23019;
    wire N__23016;
    wire N__23015;
    wire N__23012;
    wire N__23009;
    wire N__23004;
    wire N__23001;
    wire N__22998;
    wire N__22995;
    wire N__22992;
    wire N__22989;
    wire N__22988;
    wire N__22987;
    wire N__22986;
    wire N__22985;
    wire N__22978;
    wire N__22973;
    wire N__22968;
    wire N__22965;
    wire N__22962;
    wire N__22961;
    wire N__22958;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22941;
    wire N__22938;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22923;
    wire N__22922;
    wire N__22919;
    wire N__22916;
    wire N__22911;
    wire N__22908;
    wire N__22905;
    wire N__22902;
    wire N__22899;
    wire N__22896;
    wire N__22893;
    wire N__22890;
    wire N__22887;
    wire N__22884;
    wire N__22883;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22866;
    wire N__22863;
    wire N__22860;
    wire N__22859;
    wire N__22858;
    wire N__22857;
    wire N__22856;
    wire N__22855;
    wire N__22852;
    wire N__22847;
    wire N__22840;
    wire N__22833;
    wire N__22830;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22822;
    wire N__22819;
    wire N__22816;
    wire N__22813;
    wire N__22806;
    wire N__22805;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22788;
    wire N__22787;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22770;
    wire N__22767;
    wire N__22764;
    wire N__22763;
    wire N__22762;
    wire N__22759;
    wire N__22756;
    wire N__22755;
    wire N__22752;
    wire N__22751;
    wire N__22746;
    wire N__22745;
    wire N__22744;
    wire N__22743;
    wire N__22740;
    wire N__22737;
    wire N__22734;
    wire N__22731;
    wire N__22724;
    wire N__22713;
    wire N__22712;
    wire N__22707;
    wire N__22706;
    wire N__22705;
    wire N__22704;
    wire N__22703;
    wire N__22700;
    wire N__22697;
    wire N__22690;
    wire N__22683;
    wire N__22682;
    wire N__22681;
    wire N__22678;
    wire N__22673;
    wire N__22668;
    wire N__22665;
    wire N__22662;
    wire N__22659;
    wire N__22658;
    wire N__22653;
    wire N__22650;
    wire N__22649;
    wire N__22646;
    wire N__22643;
    wire N__22638;
    wire N__22637;
    wire N__22632;
    wire N__22629;
    wire N__22626;
    wire N__22623;
    wire N__22620;
    wire N__22617;
    wire N__22614;
    wire N__22611;
    wire N__22608;
    wire N__22605;
    wire N__22602;
    wire N__22599;
    wire N__22596;
    wire N__22593;
    wire N__22590;
    wire N__22587;
    wire N__22584;
    wire N__22581;
    wire N__22578;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22563;
    wire N__22560;
    wire N__22557;
    wire N__22554;
    wire N__22551;
    wire N__22548;
    wire N__22545;
    wire N__22542;
    wire N__22539;
    wire N__22536;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22518;
    wire N__22517;
    wire N__22516;
    wire N__22513;
    wire N__22510;
    wire N__22507;
    wire N__22500;
    wire N__22499;
    wire N__22496;
    wire N__22493;
    wire N__22488;
    wire N__22487;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22475;
    wire N__22474;
    wire N__22471;
    wire N__22466;
    wire N__22461;
    wire N__22458;
    wire N__22455;
    wire N__22452;
    wire N__22449;
    wire N__22446;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22434;
    wire N__22433;
    wire N__22430;
    wire N__22427;
    wire N__22424;
    wire N__22421;
    wire N__22416;
    wire N__22415;
    wire N__22414;
    wire N__22413;
    wire N__22412;
    wire N__22405;
    wire N__22400;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22374;
    wire N__22371;
    wire N__22368;
    wire N__22365;
    wire N__22362;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22329;
    wire N__22326;
    wire clock_ibuf_gb_io_gb_input;
    wire VCCG0;
    wire GNDG0;
    wire mcu_sclk_c;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net ;
    wire bfn_5_16_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_17_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_375 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_i ;
    wire N_1821_0;
    wire sdin1_c;
    wire sdin0_c;
    wire mcu_data_c;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93Z0Z_0_cascade_ ;
    wire sclk1_c;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32Z0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.un2_count_bits_1_0_a2_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_8 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ;
    wire bfn_6_18_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4 ;
    wire bfn_6_19_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_333 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_376 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.dout_read ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_237_cascade_ ;
    wire N_85_0;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_3 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_370_i ;
    wire N_1820_0;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_u_i_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.sclk_u_i_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_7;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_7;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_7_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_7 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_7_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_7 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1Z0Z_23_cascade_ ;
    wire N_29;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_read ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01Z0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_reti_0_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_8 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_369_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.csb_u_i_a2_0_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_331_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.m7_0_a2_3 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_459_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_8;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_466_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_448_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1826_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_5;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_5 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_6;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_6 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_7;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_7 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_7 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1827_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_7;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_863 ;
    wire s1_c;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_iZ0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_596_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_597 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_oZ0Z_26 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1615_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.csb_u_i_a2_0_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0 ;
    wire N_1822_0;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.csb_u_i_a2_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0 ;
    wire bfn_9_19_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_a2_1_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_21 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_22 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_op ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0 ;
    wire bfn_9_22_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_391_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_455_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_454_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_453_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_463_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_1;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_1;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_1_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_1;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_1_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_1_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_5_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_5 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_5;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_5;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_5_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_6 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_21 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_22 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.dout_op ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_12 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_15 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_10 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_391 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_8 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_1 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_10;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_3_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_3 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_3;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_3;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_3_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_3 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_31;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_31;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_31_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_31 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_31_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_31 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_28;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_29;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_30;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_31;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_31 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_3 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_3;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_4;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_4 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_4_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_4 ;
    wire bfn_11_15_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m7_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996_cascade_ ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0 ;
    wire bfn_11_19_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_3 ;
    wire sync_50hz_c;
    wire \cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config ;
    wire \cemf_module_64ch_ctrl_inst1.N_410_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.N_68_0_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_8;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_8;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_8_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_8 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_8 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_8_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_8 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_14;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_14;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_14_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_14;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_14_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_14_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_14 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_22;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_30;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_30;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_30_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_30 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_30_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_30 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_30 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_30 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_30;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_31;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_31 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_31;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_4 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_4;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_26;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_26;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_26;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_0_26 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_1_26_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_26;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_21;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_9;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_29;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_3;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_907 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_30;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_621 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_31;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_610 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_1;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_316 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_5;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_885 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_6;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_874 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_9;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_9;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_4;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_4;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_4 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_9;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_30;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_4;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_8;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_0;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_11;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_12;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_13;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_14;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_786 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_15;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_20;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15Z0Z_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_19 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_i_a2_1_1_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9 ;
    wire bfn_12_20_0_;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.en_ch_cnt_0_a2_0_a2_1 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1867_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un40_0_a2_4_a2_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16 ;
    wire sda_o;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_22_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_22 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_22;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_22;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_22 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_22 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_22 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_28;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_28;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_28_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_28 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_28_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_28 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_28 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_15;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_15;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_15_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_15;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_775 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_15_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_15_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_15 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_23;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_17;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_17;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_17_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_17;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_17_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_17_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_17 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_25;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_4_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_4_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_data_config_4;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRLZ0Z7_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_6_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_6 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_6 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_6;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_6;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_6 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_841 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_9_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_6_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3QZ0Z5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_5 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net ;
    wire \cemf_module_64ch_ctrl_inst1.N_1615 ;
    wire N_1614_cascade_;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_28;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_643 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_5 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_4;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_896 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_291_reti_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_276i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_retZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_4_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_2_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_0_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_o3_i_a2_1_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_5 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ns_i_a2_1_1_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_2 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_2_cascade_ ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_10 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net ;
    wire \cemf_module_64ch_ctrl_inst1.N_68_0 ;
    wire \cemf_module_64ch_ctrl_inst1.N_410_0 ;
    wire \cemf_module_64ch_ctrl_inst1.c_state_7 ;
    wire bfn_13_23_0_;
    wire \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_2 ;
    wire \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetterZ0 ;
    wire \INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC_net ;
    wire \I2C_top_level_inst1.I2C_Control_StartUp_inst.rst_neg_i ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_22 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_2;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_13;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_13;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_13_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_13;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_797 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_13_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_13 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_13_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_18;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_18;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_18_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_18_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_18 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_18 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_13 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_15 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_13_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3QZ0Z5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_4 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_4 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_9 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_9;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_22;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3Z0Z_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1959_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0_cascade_ ;
    wire \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net ;
    wire \I2C_top_level_inst1.I2C_Control_StartUp_inst.N_8_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.en_count_bits_0_i_a2_0_a2_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_277_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_18 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967i_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_276_reti ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_8_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_4 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_2_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1945 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1844 ;
    wire N_528_0;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.n_state41 ;
    wire \cemf_module_64ch_ctrl_inst1.c_state_19 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_3 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_2 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_275_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_275_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_2_cascade_ ;
    wire \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_59 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_2 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_2;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_2;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_2_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_2_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_2 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_10;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_10;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_10_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_10;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_830 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_10_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_10 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_10_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_10 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_18;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_18 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_11;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_11;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_11_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_11;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_819 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_11_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_11_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_19;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_20;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_20;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_20_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_20;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_283 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_20_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_20_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_6 ;
    wire cemf_module_64ch_ctrl_inst1_data_config_6;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_6_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRLZ0Z7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_7 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_6 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_6;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_5;
    wire cemf_module_64ch_ctrl_inst1_data_config_5;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRLZ0Z7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_5 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_5;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_14;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_242_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_5;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_16;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_18;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1911 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_8;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1920 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m20_0_a2_4_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_11_0_i_0_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1394_cascade_ ;
    wire s_sda_i_g;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1392 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1381_0_cascade_ ;
    wire \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392 ;
    wire \cemf_module_64ch_ctrl_inst1.c_state_i_2_2 ;
    wire \cemf_module_64ch_ctrl_inst1.end_conf_a ;
    wire \cemf_module_64ch_ctrl_inst1.N_1817_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2_8 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_0_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1873_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1874_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_2_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1950 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1949_cascade_ ;
    wire stop_fpga2_c;
    wire \cemf_module_64ch_ctrl_inst1.end_conf_b ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847 ;
    wire \serializer_mod_inst.shift_regZ0Z_112 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_4 ;
    wire \serializer_mod_inst.shift_regZ0Z_111 ;
    wire \serializer_mod_inst.shift_regZ0Z_119 ;
    wire \serializer_mod_inst.shift_regZ0Z_120 ;
    wire \serializer_mod_inst.shift_regZ0Z_36 ;
    wire \serializer_mod_inst.shift_regZ0Z_118 ;
    wire \serializer_mod_inst.shift_regZ0Z_37 ;
    wire \serializer_mod_inst.shift_regZ0Z_38 ;
    wire \serializer_mod_inst.shift_regZ0Z_33 ;
    wire \serializer_mod_inst.shift_regZ0Z_34 ;
    wire \serializer_mod_inst.shift_regZ0Z_35 ;
    wire \serializer_mod_inst.shift_regZ0Z_76 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_17;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_753 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_19;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_2;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_918 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_22;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_698 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_23;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_2 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_25;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_19;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_19;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_731 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_19 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_19_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_19 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_19 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_19 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_0;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_0;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_0_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_21;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_1 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_18;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_18 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_20;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_20 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_15_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_14 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_14_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGHZ0Z5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_14_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_14 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_14;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_23_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDDZ0Z7_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_6;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_6 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_3;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_4;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_6;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_0Z0Z_26 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_30;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1654_cascade_ ;
    wire N_12_0_cascade_;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_7;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0_cascade_ ;
    wire N_12_0;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_0_7 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_1786_2 ;
    wire N_979;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_id_prdata_1_4_u_i_0;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2_cascade_;
    wire N_1838_0_cascade_;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1379_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1400_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1374_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6 ;
    wire \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1399_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1395_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_0_10 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_14 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1409_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1372_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14 ;
    wire \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1880 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1848_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1884_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392_reti ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0_a2_6_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_2 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_li_0_1 ;
    wire c_state_ret_12_RNIDMPS1_0;
    wire c_state_ret_12_RNIDMPS1_0_cascade_;
    wire \cemf_module_64ch_ctrl_inst1.clr_sys_reg ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_1;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_349 ;
    wire \serializer_mod_inst.shift_regZ0Z_7 ;
    wire \serializer_mod_inst.shift_regZ0Z_31 ;
    wire \serializer_mod_inst.shift_regZ0Z_32 ;
    wire \serializer_mod_inst.shift_regZ0Z_113 ;
    wire \serializer_mod_inst.shift_regZ0Z_114 ;
    wire \serializer_mod_inst.shift_regZ0Z_110 ;
    wire \serializer_mod_inst.shift_regZ0Z_39 ;
    wire \serializer_mod_inst.shift_regZ0Z_77 ;
    wire \serializer_mod_inst.shift_regZ0Z_78 ;
    wire \serializer_mod_inst.shift_regZ0Z_40 ;
    wire \serializer_mod_inst.shift_regZ0Z_67 ;
    wire \serializer_mod_inst.shift_regZ0Z_68 ;
    wire \serializer_mod_inst.shift_regZ0Z_115 ;
    wire \serializer_mod_inst.shift_regZ0Z_116 ;
    wire \serializer_mod_inst.shift_regZ0Z_117 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa ;
    wire rst_n_c_i;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_12;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_12;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_12_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_12;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_808 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_12_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_12 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_12_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_12 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_11;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_11 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_12;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_12 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_13;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_13 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_14;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_14 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_15;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_15 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_16;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_17;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_17 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_2;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_2 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_24;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_24;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_19;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_19 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_25;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_27;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_28;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_28 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_28;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_29;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_29;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_3;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_3 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_3;
    wire serial_out_testing_c;
    wire rst_n_c;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1965 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_522_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4 ;
    wire \cemf_module_64ch_ctrl_inst1.start_conf_b ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_20;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_20_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DDZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_21 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_22 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_conf ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1831_0 ;
    wire N_1614;
    wire N_1841_0_cascade_;
    wire N_1613_cascade_;
    wire N_1860_0;
    wire N_202_0;
    wire N_1859_0;
    wire N_1861_0;
    wire N_1613;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_604 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0_cascade_ ;
    wire \I2C_top_level_inst1.s_command_4 ;
    wire \I2C_top_level_inst1.s_command_5 ;
    wire \I2C_top_level_inst1.s_command_6 ;
    wire N_1803;
    wire N_1803_cascade_;
    wire \I2C_top_level_inst1.s_command_7 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6Z0Z_26 ;
    wire \I2C_top_level_inst1.N_327_i ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_113_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_6 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4 ;
    wire \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_3_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_5_1 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_2_1 ;
    wire \I2C_top_level_inst1.N_4_0_cascade_ ;
    wire \I2C_top_level_inst1.N_259 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1848_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7Z0Z_26 ;
    wire \I2C_top_level_inst1.s_sda_o_qZ0Z_1 ;
    wire \I2C_top_level_inst1.s_sda_o_txZ0 ;
    wire \I2C_top_level_inst1.s_sda_o_qZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.start_conf_a ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1855_0 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1855_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1857_0 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1857_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_384 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1854_0 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1840_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0 ;
    wire \cemf_module_64ch_ctrl_inst1.N_383 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8Z0Z_26 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ;
    wire \cemf_module_64ch_ctrl_inst1.c_state_12 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1862 ;
    wire \cemf_module_64ch_ctrl_inst1.N_1816_0 ;
    wire \cemf_module_64ch_ctrl_inst1.c_state_8 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_reti_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_6 ;
    wire \serializer_mod_inst.shift_regZ0Z_11 ;
    wire \serializer_mod_inst.shift_regZ0Z_48 ;
    wire \serializer_mod_inst.shift_regZ0Z_51 ;
    wire \serializer_mod_inst.shift_regZ0Z_10 ;
    wire \serializer_mod_inst.shift_regZ0Z_55 ;
    wire \serializer_mod_inst.shift_regZ0Z_121 ;
    wire \serializer_mod_inst.shift_regZ0Z_14 ;
    wire \serializer_mod_inst.shift_regZ0Z_12 ;
    wire \serializer_mod_inst.shift_regZ0Z_13 ;
    wire \serializer_mod_inst.shift_regZ0Z_8 ;
    wire \serializer_mod_inst.shift_regZ0Z_9 ;
    wire \serializer_mod_inst.shift_regZ0Z_15 ;
    wire \serializer_mod_inst.shift_regZ0Z_79 ;
    wire \serializer_mod_inst.shift_regZ0Z_16 ;
    wire \serializer_mod_inst.shift_regZ0Z_17 ;
    wire \serializer_mod_inst.shift_regZ0Z_18 ;
    wire \serializer_mod_inst.shift_regZ0Z_107 ;
    wire \serializer_mod_inst.shift_regZ0Z_69 ;
    wire \serializer_mod_inst.shift_regZ0Z_106 ;
    wire \serializer_mod_inst.shift_regZ0Z_47 ;
    wire \serializer_mod_inst.shift_regZ0Z_94 ;
    wire \serializer_mod_inst.shift_regZ0Z_104 ;
    wire \serializer_mod_inst.shift_regZ0Z_105 ;
    wire \serializer_mod_inst.shift_regZ0Z_46 ;
    wire \serializer_mod_inst.shift_regZ0Z_91 ;
    wire \serializer_mod_inst.shift_regZ0Z_92 ;
    wire \serializer_mod_inst.shift_regZ0Z_93 ;
    wire \serializer_mod_inst.shift_regZ0Z_95 ;
    wire \serializer_mod_inst.shift_regZ0Z_96 ;
    wire \serializer_mod_inst.shift_regZ0Z_97 ;
    wire enable_config_c;
    wire elec_config_out_c;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_24 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_24_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_24 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_24;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_24;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_24_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_24 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_23;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_10;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_10 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_24;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_676 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_23 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_687 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_23 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_23_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_23 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_23;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_23;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_23_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_23 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_20 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_21;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_21;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_21_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_21;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1320 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1896 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_21_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_21 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_21 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_21_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_21 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_30;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_13;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_31;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_14;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_22_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_22 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_22;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_22_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDDZ0Z7 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_22;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_22 ;
    wire cemf_module_64ch_ctrl_inst1_data_config_20;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_30;
    wire cemf_module_64ch_ctrl_inst1_data_config_22;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_8_0_m2_ns_1_cascade_ ;
    wire N_1842_0;
    wire N_1842_0_cascade_;
    wire N_1841_0;
    wire \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C_net ;
    wire bfn_18_18_0_;
    wire \cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0 ;
    wire \cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_CO ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1 ;
    wire \cemf_module_64ch_ctrl_inst1.c_addr_RNI3UAS1_6 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2 ;
    wire \cemf_module_64ch_ctrl_inst1.c_addr_RNI50BS1_7 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93STZ0Z1 ;
    wire CONSTANT_ONE_NET;
    wire \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rstZ0 ;
    wire \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNOZ0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_3_cascade_ ;
    wire N_1975;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNOZ0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0 ;
    wire bfn_18_20_0_;
    wire \cemf_module_64ch_ctrl_inst1.paddr_fsm_1 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_2;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_3;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_4;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_5;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_6;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_7 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_8;
    wire bfn_18_21_0_;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_9;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_10;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_11;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_12;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_13;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_14;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_14 ;
    wire cemf_module_64ch_ctrl_inst1_paddr_fsm_15;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0 ;
    wire \serializer_mod_inst.shift_regZ0Z_86 ;
    wire \serializer_mod_inst.shift_regZ0Z_54 ;
    wire cemf_module_64ch_ctrl_inst1_s_data_system_o_0;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6 ;
    wire \serializer_mod_inst.shift_regZ0Z_52 ;
    wire \serializer_mod_inst.shift_regZ0Z_53 ;
    wire \serializer_mod_inst.shift_regZ0Z_87 ;
    wire \serializer_mod_inst.shift_regZ0Z_88 ;
    wire \serializer_mod_inst.shift_regZ0Z_49 ;
    wire \serializer_mod_inst.shift_regZ0Z_50 ;
    wire \serializer_mod_inst.shift_regZ0Z_89 ;
    wire \serializer_mod_inst.shift_regZ0Z_90 ;
    wire \serializer_mod_inst.shift_regZ0Z_85 ;
    wire \serializer_mod_inst.shift_regZ0Z_1 ;
    wire \serializer_mod_inst.shift_regZ0Z_101 ;
    wire \serializer_mod_inst.shift_regZ0Z_66 ;
    wire \serializer_mod_inst.shift_regZ0Z_102 ;
    wire \serializer_mod_inst.shift_regZ0Z_103 ;
    wire \serializer_mod_inst.shift_regZ0Z_84 ;
    wire \serializer_mod_inst.shift_regZ0Z_41 ;
    wire \serializer_mod_inst.shift_regZ0Z_100 ;
    wire \serializer_mod_inst.shift_regZ0Z_42 ;
    wire \serializer_mod_inst.shift_regZ0Z_43 ;
    wire \serializer_mod_inst.shift_regZ0Z_44 ;
    wire \serializer_mod_inst.shift_regZ0Z_45 ;
    wire \serializer_mod_inst.shift_regZ0Z_70 ;
    wire \serializer_mod_inst.shift_regZ0Z_71 ;
    wire \serializer_mod_inst.shift_regZ0Z_74 ;
    wire \serializer_mod_inst.shift_regZ0Z_75 ;
    wire \serializer_mod_inst.shift_regZ0Z_98 ;
    wire \serializer_mod_inst.shift_regZ0Z_99 ;
    wire \serializer_mod_inst.shift_regZ0Z_72 ;
    wire \serializer_mod_inst.shift_regZ0Z_73 ;
    wire \serializer_mod_inst.shift_regZ0Z_83 ;
    wire \serializer_mod_inst.shift_regZ0Z_82 ;
    wire \serializer_mod_inst.shift_regZ0Z_80 ;
    wire \serializer_mod_inst.shift_regZ0Z_81 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_29;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_29;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_29_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_29 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_29 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_29_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_632 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_29 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_29 ;
    wire cemf_module_64ch_ctrl_inst1_data_config_7;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_8_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_6 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_7 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_24;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_28;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_1Z0Z_26 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_27;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_7 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_7;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_8 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_8;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_8;
    wire cemf_module_64ch_ctrl_inst1_data_config_8;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_8_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8DZ0Z7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14_cascade_ ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_8;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_20 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_3 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_20;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_12;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_0_12_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_2_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_0_i_12_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_13 ;
    wire cemf_module_64ch_ctrl_inst1_data_config_13;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_13 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_5;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_6;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_7;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_8;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_12 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_config_12;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_12;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_12 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_11_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFHZ0Z5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0_cascade_ ;
    wire \I2C_top_level_inst1.s_addr1_o_1 ;
    wire \I2C_top_level_inst1.s_addr1_o_2 ;
    wire \I2C_top_level_inst1.s_addr1_o_3 ;
    wire \I2C_top_level_inst1.s_addr1_o_4 ;
    wire \I2C_top_level_inst1.s_addr1_o_5 ;
    wire \I2C_top_level_inst1.s_addr1_o_6 ;
    wire \I2C_top_level_inst1.s_addr1_o_7 ;
    wire \I2C_top_level_inst1.s_load_addr1 ;
    wire \I2C_top_level_inst1.s_addr0_o_3 ;
    wire \I2C_top_level_inst1.s_data_ireg_4 ;
    wire \I2C_top_level_inst1.s_addr0_o_4 ;
    wire \I2C_top_level_inst1.s_data_ireg_5 ;
    wire \I2C_top_level_inst1.s_addr0_o_5 ;
    wire \I2C_top_level_inst1.s_data_ireg_6 ;
    wire \I2C_top_level_inst1.s_addr0_o_6 ;
    wire \I2C_top_level_inst1.s_data_ireg_7 ;
    wire \I2C_top_level_inst1.s_addr0_o_7 ;
    wire N_396;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_3 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_4_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNOZ0Z_0_cascade_ ;
    wire \I2C_top_level_inst1.s_no_restart ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_304_0 ;
    wire \I2C_top_level_inst1.s_ack ;
    wire \serializer_mod_inst.shift_regZ0Z_6 ;
    wire \serializer_mod_inst.shift_regZ0Z_5 ;
    wire \serializer_mod_inst.shift_regZ0Z_2 ;
    wire \serializer_mod_inst.shift_regZ0Z_3 ;
    wire \serializer_mod_inst.shift_regZ0Z_4 ;
    wire \serializer_mod_inst.shift_regZ0Z_21 ;
    wire \serializer_mod_inst.shift_regZ0Z_27 ;
    wire \serializer_mod_inst.shift_regZ0Z_22 ;
    wire \serializer_mod_inst.shift_regZ0Z_23 ;
    wire \serializer_mod_inst.shift_regZ0Z_108 ;
    wire \serializer_mod_inst.shift_regZ0Z_109 ;
    wire \serializer_mod_inst.shift_regZ0Z_19 ;
    wire \serializer_mod_inst.shift_regZ0Z_20 ;
    wire \serializer_mod_inst.shift_regZ0Z_24 ;
    wire \serializer_mod_inst.shift_regZ0Z_124 ;
    wire \serializer_mod_inst.shift_regZ0Z_125 ;
    wire \serializer_mod_inst.shift_regZ0Z_122 ;
    wire \serializer_mod_inst.shift_regZ0Z_123 ;
    wire \serializer_mod_inst.shift_regZ0Z_25 ;
    wire \serializer_mod_inst.shift_regZ0Z_26 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_27;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_27_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_27 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_27 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_27_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_654 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_27 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_27 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_16;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_16;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_16_cascade_ ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_16;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_16;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_764 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_16_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_16 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_16 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_16_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_16 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_24;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_24 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_22;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_4;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_5;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_6;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_15_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_14 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_15 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_4;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_20;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_20;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_12;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_22;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_14;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_15;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_16;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_11;
    wire cemf_module_64ch_ctrl_inst1_data_config_11;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_11_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_13 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_13;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_23 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_10;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_10;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_2;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_2;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_11;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_11 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_11;
    wire bfn_20_17_0_;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_CO ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_4 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_6 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_7 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7 ;
    wire bfn_20_18_0_;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_10 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_12 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_13 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_15 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_103_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_0 ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_291_cascade_ ;
    wire \I2C_top_level_inst1.s_load_addr0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_6_0_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1378 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_1676_cascade_ ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21;
    wire c_state_RNIEVJ7_22_cascade_;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_77_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_300_6 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_FSM_inst.N_1425_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_3 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0 ;
    wire \serializer_mod_inst.shift_regZ0Z_64 ;
    wire \serializer_mod_inst.shift_regZ0Z_65 ;
    wire \serializer_mod_inst.shift_regZ0Z_128 ;
    wire \serializer_mod_inst.shift_regZ0Z_126 ;
    wire \serializer_mod_inst.shift_regZ0Z_127 ;
    wire \serializer_mod_inst.shift_regZ0Z_28 ;
    wire \serializer_mod_inst.shift_regZ0Z_29 ;
    wire \serializer_mod_inst.shift_regZ0Z_30 ;
    wire \serializer_mod_inst.shift_regZ0Z_62 ;
    wire \serializer_mod_inst.shift_regZ0Z_63 ;
    wire \serializer_mod_inst.shift_regZ0Z_58 ;
    wire \serializer_mod_inst.shift_regZ0Z_59 ;
    wire \serializer_mod_inst.shift_regZ0Z_60 ;
    wire \serializer_mod_inst.shift_regZ0Z_61 ;
    wire \serializer_mod_inst.shift_regZ0Z_56 ;
    wire \serializer_mod_inst.shift_regZ0Z_57 ;
    wire \serializer_mod_inst.un22_next_state_1_cascade_ ;
    wire \serializer_mod_inst.un22_next_state ;
    wire \serializer_mod_inst.current_stateZ0Z_1 ;
    wire \serializer_mod_inst.current_stateZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_0;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_940 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_25;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_3Z0Z_26 ;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_16 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_7;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_7 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_17_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_16 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_17;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_11 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_21_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LHZ0Z5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_21 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_21;
    wire cemf_module_64ch_ctrl_inst1_data_config_21;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_21_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDDZ0Z7 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_21;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_21;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_21 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_11;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_12;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_21;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_30;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_13;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_31;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_15;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_13;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_31;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_15;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_24;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_17;
    wire I2C_top_level_inst1_s_data_oreg_9;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_10 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_9;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_9;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i_cascade_ ;
    wire s_paddr_I2C_5;
    wire s_paddr_I2C_4;
    wire s_paddr_I2C_6;
    wire s_paddr_I2C_7;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_5 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_3 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_2_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_1_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0_cascade_ ;
    wire s_paddr_I2C_2;
    wire s_paddr_I2C_1;
    wire s_paddr_I2C_0;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_7_3_i_a2_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0 ;
    wire \I2C_top_level_inst1.s_addr1_o_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_8_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_CO ;
    wire \I2C_top_level_inst1.s_addr0_o_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1651 ;
    wire \I2C_top_level_inst1.s_addr0_o_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1652 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_0_4_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_0_1_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_279_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_0_1_7_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_268_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_10_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_18_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1605_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0 ;
    wire \I2C_top_level_inst1.s_data_ireg_0 ;
    wire \I2C_top_level_inst1.s_command_0 ;
    wire \I2C_top_level_inst1.s_data_ireg_1 ;
    wire \I2C_top_level_inst1.s_data_ireg_2 ;
    wire \I2C_top_level_inst1.s_data_ireg_3 ;
    wire scl_c_g;
    wire \I2C_top_level_inst1.s_load_command ;
    wire \serializer_mod_inst.un1_counter_srlto6_3 ;
    wire \serializer_mod_inst.un1_counter_srlto6_4_cascade_ ;
    wire \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ;
    wire \serializer_mod_inst.un22_next_state_5 ;
    wire \serializer_mod_inst.counter_srZ0Z_0 ;
    wire bfn_21_27_0_;
    wire \serializer_mod_inst.counter_srZ0Z_1 ;
    wire \serializer_mod_inst.counter_sr_cry_0 ;
    wire \serializer_mod_inst.counter_srZ0Z_2 ;
    wire \serializer_mod_inst.counter_sr_cry_1 ;
    wire \serializer_mod_inst.counter_srZ0Z_3 ;
    wire \serializer_mod_inst.counter_sr_cry_2 ;
    wire \serializer_mod_inst.counter_srZ0Z_4 ;
    wire \serializer_mod_inst.counter_sr_cry_3 ;
    wire \serializer_mod_inst.counter_srZ0Z_5 ;
    wire \serializer_mod_inst.counter_sr_cry_4 ;
    wire \serializer_mod_inst.counter_srZ0Z_6 ;
    wire \serializer_mod_inst.counter_sr_cry_5 ;
    wire \serializer_mod_inst.next_state32_i ;
    wire \serializer_mod_inst.counter_sr_cry_6 ;
    wire \serializer_mod_inst.counter_srZ0Z_7 ;
    wire \serializer_mod_inst.counter_sre_0_i ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_15;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_24;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_2Z0Z_26 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_28;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_29;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_7;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_19;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_19;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_0;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_0;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_18;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_18_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9DZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_19 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_18;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_28;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_29;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_23;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_23;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_23_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.dout_conf ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALHZ0Z5 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_21 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_22 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_23;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_23;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_23 ;
    wire cemf_module_64ch_ctrl_inst1_data_config_9;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_9;
    wire cemf_module_64ch_ctrl_inst1_data_config_10;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_10;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_10;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_10_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_10 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_9;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_8 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_9 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_2;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_3;
    wire cemf_module_64ch_ctrl_inst1_data_config_3;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_3;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_3 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_2;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_2 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_6_0_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_607 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_15_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_1_15 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_322 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_267 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_394 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_267_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_1_1_i_m2_1_9_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_101 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_1_2_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_372_cascade_ ;
    wire N_409;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_a3_1_0_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_412_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_1_14 ;
    wire N_410;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_1_0_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_25 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_24_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_11_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_11_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_2_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_86_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_95_0 ;
    wire \I2C_top_level_inst1.s_stop ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_844_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1754_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_1 ;
    wire scl_c;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0 ;
    wire \I2C_top_level_inst1.s_command_1 ;
    wire \I2C_top_level_inst1.s_command_2 ;
    wire \I2C_top_level_inst1.s_command_3 ;
    wire \I2C_top_level_inst1.s_load_wdata ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2 ;
    wire \I2C_top_level_inst1.s_start ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_1 ;
    wire \I2C_top_level_inst1.s_r_w ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_27;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_29;
    wire cemf_module_64ch_ctrl_inst1_data_config_23;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_19 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_19;
    wire cemf_module_64ch_ctrl_inst1_data_config_19;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_19 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_18;
    wire cemf_module_64ch_ctrl_inst1_data_config_18;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_18;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_18_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_18 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_25;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_25;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_25;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_25;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_25;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_25_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_25 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_25 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_25_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_665 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_25;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_25 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_25 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_16;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_17;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_17;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_17_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_17 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_16;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGHZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_15 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_16 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net ;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_31;
    wire cemf_module_64ch_ctrl_inst1_data_config_14;
    wire cemf_module_64ch_ctrl_inst1_data_config_15;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_24;
    wire cemf_module_64ch_ctrl_inst1_data_config_16;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_28;
    wire cemf_module_64ch_ctrl_inst1_data_config_17;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273 ;
    wire cemf_module_64ch_ctrl_inst1_data_config_2;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RLZ0Z7_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_2 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270 ;
    wire cemf_module_64ch_ctrl_inst1_data_clkstopmask_1;
    wire cemf_module_64ch_ctrl_inst1_data_clkctrovf_1;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_3_26 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_4093_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_26 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_g ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0 ;
    wire s_paddr_I2C_3;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_230_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_0_sqmuxa ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_2_sqmuxa ;
    wire s_paddr_I2C_8;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_230 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_4 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_365_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_4_0_a2_2_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_676_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_address ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1606_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1565_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_5_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_6_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_7_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_11_0_cascade_ ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_23_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_288 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_288_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_23 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_115 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_904 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un30_i_a2_9_a2_4_a2_0_1_2_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_291 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_0_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_232_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_2_1_cascade_ ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_20;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_4_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_232 ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_1_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_2_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_231 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_212 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_211 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1653_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_122_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_208 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_239 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_239_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_294 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_1_0_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_0_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1776 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_209 ;
    wire s_sda_i;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_0 ;
    wire I2C_top_level_inst1_s_data_oreg_16;
    wire I2C_top_level_inst1_s_data_oreg_15;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_15 ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_16 ;
    wire I2C_top_level_inst1_s_data_oreg_17;
    wire \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_19;
    wire cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_29;
    wire N_1592_0;
    wire \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0 ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_9 ;
    wire I2C_top_level_inst1_s_data_oreg_10;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_10 ;
    wire I2C_top_level_inst1_s_data_oreg_11;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_11 ;
    wire I2C_top_level_inst1_s_data_oreg_12;
    wire I2C_top_level_inst1_s_data_oreg_14;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_14 ;
    wire I2C_top_level_inst1_s_data_oreg_13;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_12 ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_13 ;
    wire \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_0;
    wire cemf_module_64ch_ctrl_inst1_data_config_0;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273 ;
    wire cemf_module_64ch_ctrl_inst1_data_interrupts_1;
    wire cemf_module_64ch_ctrl_inst1_data_config_1;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_1;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_1 ;
    wire cemf_module_64ch_ctrl_inst1_data_coarseovf_0;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2QZ0Z5_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0_cascade_ ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_0 ;
    wire \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net ;
    wire \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i ;
    wire I2C_top_level_inst1_s_data_oreg_18;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_17 ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_18 ;
    wire I2C_top_level_inst1_s_data_oreg_19;
    wire I2C_top_level_inst1_s_data_oreg_20;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_19 ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_20 ;
    wire I2C_top_level_inst1_s_data_oreg_21;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_21 ;
    wire I2C_top_level_inst1_s_data_oreg_22;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_22 ;
    wire I2C_top_level_inst1_s_data_oreg_23;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_23 ;
    wire I2C_top_level_inst1_s_data_oreg_24;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_24 ;
    wire I2C_top_level_inst1_s_data_oreg_25;
    wire \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_25 ;
    wire I2C_top_level_inst1_s_data_oreg_26;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_26 ;
    wire I2C_top_level_inst1_s_data_oreg_27;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_27 ;
    wire I2C_top_level_inst1_s_data_oreg_28;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_28 ;
    wire I2C_top_level_inst1_s_data_oreg_29;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_29 ;
    wire I2C_top_level_inst1_s_data_oreg_30;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_30 ;
    wire I2C_top_level_inst1_s_data_oreg_31;
    wire \I2C_top_level_inst1.s_sda_o_reg ;
    wire I2C_top_level_inst1_s_data_oreg_0;
    wire \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_0 ;
    wire I2C_top_level_inst1_s_data_oreg_1;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_1 ;
    wire I2C_top_level_inst1_s_data_oreg_2;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_2 ;
    wire I2C_top_level_inst1_s_data_oreg_3;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_3 ;
    wire I2C_top_level_inst1_s_data_oreg_4;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_4 ;
    wire I2C_top_level_inst1_s_data_oreg_5;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_5 ;
    wire I2C_top_level_inst1_s_data_oreg_6;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_6 ;
    wire I2C_top_level_inst1_s_data_oreg_7;
    wire \I2C_top_level_inst1.s_enable_desp_tx ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_7 ;
    wire I2C_top_level_inst1_s_data_oreg_8;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_8 ;
    wire \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ;
    wire \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0 ;
    wire rst_n_c_i_g;
    wire c_state_RNIEVJ7_22;
    wire \I2C_top_level_inst1.s_load_rdata2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o3_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1802 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1609_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0 ;
    wire \I2C_top_level_inst1.s_addr0_o_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_691 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_295_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_6 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0 ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_277 ;
    wire N_552_i;
    wire N_1838_0;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_295 ;
    wire N_73_i_0_cascade_;
    wire I2C_top_level_inst1_s_burst;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_19 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_274_cascade_ ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19 ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2 ;
    wire I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_276 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_245 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1669_cascade_ ;
    wire clock_c_g;
    wire \I2C_top_level_inst1.c_state4_0_i_g ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_2_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_0_2_cascade_ ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0 ;
    wire \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666_2 ;
    wire _gnd_net_;

    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_15,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_14,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_13,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_12,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_11,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_10,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_9,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_8,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_7,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_6,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_5,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_4,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_3,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_2,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_1,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_0}),
            .RADDR({dangling_wire_0,dangling_wire_1,dangling_wire_2,dangling_wire_3,dangling_wire_4,N__24740,N__24935,N__25112,N__25316,N__36044,N__25214}),
            .WADDR({dangling_wire_5,dangling_wire_6,dangling_wire_7,dangling_wire_8,dangling_wire_9,N__24731,N__24932,N__25109,N__25313,N__36041,N__25211}),
            .MASK({dangling_wire_10,dangling_wire_11,dangling_wire_12,dangling_wire_13,dangling_wire_14,dangling_wire_15,dangling_wire_16,dangling_wire_17,dangling_wire_18,dangling_wire_19,dangling_wire_20,dangling_wire_21,dangling_wire_22,dangling_wire_23,dangling_wire_24,dangling_wire_25}),
            .WDATA({N__23921,N__23963,N__24005,N__24042,N__24483,N__24697,N__24275,N__26186,N__33976,N__26384,N__24353,N__24392,N__23798,N__24619,N__23684,N__23721}),
            .RCLKE(),
            .RCLK(N__65640),
            .RE(N__39325),
            .WCLKE(N__24887),
            .WCLK(N__65641),
            .WE(N__39314));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_31,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_30,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_29,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_28,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_27,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_26,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_25,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_24,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_23,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_22,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_21,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_20,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_19,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_18,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_17,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_16}),
            .RADDR({dangling_wire_26,dangling_wire_27,dangling_wire_28,dangling_wire_29,dangling_wire_30,N__24728,N__24923,N__25100,N__25304,N__36032,N__25202}),
            .WADDR({dangling_wire_31,dangling_wire_32,dangling_wire_33,dangling_wire_34,dangling_wire_35,N__24719,N__24920,N__25097,N__25301,N__36029,N__25199}),
            .MASK({dangling_wire_36,dangling_wire_37,dangling_wire_38,dangling_wire_39,dangling_wire_40,dangling_wire_41,dangling_wire_42,dangling_wire_43,dangling_wire_44,dangling_wire_45,dangling_wire_46,dangling_wire_47,dangling_wire_48,dangling_wire_49,dangling_wire_50,dangling_wire_51}),
            .WDATA({N__26553,N__24666,N__24077,N__24445,N__24533,N__24158,N__24240,N__24584,N__24198,N__24317,N__24119,N__23841,N__26424,N__26469,N__26514,N__23883}),
            .RCLKE(),
            .RCLK(N__65665),
            .RE(N__39296),
            .WCLKE(N__24891),
            .WCLK(N__65666),
            .WE(N__39305));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_31,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_30,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_29,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_28,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_27,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_26,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_25,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_24,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_23,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_22,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_21,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_20,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_19,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_18,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_17,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_16}),
            .RADDR({dangling_wire_52,dangling_wire_53,dangling_wire_54,dangling_wire_55,dangling_wire_56,N__24800,N__24995,N__25172,N__25376,N__36104,N__25274}),
            .WADDR({dangling_wire_57,dangling_wire_58,dangling_wire_59,dangling_wire_60,dangling_wire_61,N__24791,N__24992,N__25169,N__25373,N__36101,N__25271}),
            .MASK({dangling_wire_62,dangling_wire_63,dangling_wire_64,dangling_wire_65,dangling_wire_66,dangling_wire_67,dangling_wire_68,dangling_wire_69,dangling_wire_70,dangling_wire_71,dangling_wire_72,dangling_wire_73,dangling_wire_74,dangling_wire_75,dangling_wire_76,dangling_wire_77}),
            .WDATA({N__26552,N__24665,N__24078,N__24459,N__24534,N__24159,N__24239,N__24588,N__24197,N__24318,N__24120,N__23840,N__26419,N__26464,N__26509,N__23882}),
            .RCLKE(),
            .RCLK(N__65524),
            .RE(N__39401),
            .WCLKE(N__23739),
            .WCLK(N__65525),
            .WE(N__39396));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_15,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_14,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_13,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_12,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_11,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_10,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_9,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_8,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_7,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_6,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_5,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_4,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_3,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_2,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_1,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_0}),
            .RADDR({dangling_wire_78,dangling_wire_79,dangling_wire_80,dangling_wire_81,dangling_wire_82,N__24807,N__25005,N__25182,N__25386,N__36114,N__25284}),
            .WADDR({dangling_wire_83,dangling_wire_84,dangling_wire_85,dangling_wire_86,dangling_wire_87,N__24803,N__25004,N__25181,N__25385,N__36113,N__25283}),
            .MASK({dangling_wire_88,dangling_wire_89,dangling_wire_90,dangling_wire_91,dangling_wire_92,dangling_wire_93,dangling_wire_94,dangling_wire_95,dangling_wire_96,dangling_wire_97,dangling_wire_98,dangling_wire_99,dangling_wire_100,dangling_wire_101,dangling_wire_102,dangling_wire_103}),
            .WDATA({N__23922,N__23964,N__24006,N__24041,N__24495,N__24702,N__24279,N__26187,N__34005,N__26385,N__24354,N__24393,N__23799,N__24624,N__23685,N__23720}),
            .RCLKE(),
            .RCLK(N__65515),
            .RE(N__39402),
            .WCLKE(N__23732),
            .WCLK(N__65516),
            .WE(N__39400));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_31,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_30,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_29,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_28,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_27,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_26,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_25,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_24,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_23,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_22,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_21,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_20,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_19,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_18,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_17,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_16}),
            .RADDR({dangling_wire_104,dangling_wire_105,dangling_wire_106,dangling_wire_107,dangling_wire_108,N__24752,N__24947,N__25124,N__25328,N__36056,N__25226}),
            .WADDR({dangling_wire_109,dangling_wire_110,dangling_wire_111,dangling_wire_112,dangling_wire_113,N__24743,N__24944,N__25121,N__25325,N__36053,N__25223}),
            .MASK({dangling_wire_114,dangling_wire_115,dangling_wire_116,dangling_wire_117,dangling_wire_118,dangling_wire_119,dangling_wire_120,dangling_wire_121,dangling_wire_122,dangling_wire_123,dangling_wire_124,dangling_wire_125,dangling_wire_126,dangling_wire_127,dangling_wire_128,dangling_wire_129}),
            .WDATA({N__26548,N__24661,N__24069,N__24430,N__24513,N__24150,N__24235,N__24564,N__24193,N__24310,N__24117,N__23836,N__26420,N__26465,N__26510,N__23878}),
            .RCLKE(),
            .RCLK(N__65614),
            .RE(N__39336),
            .WCLKE(N__24549),
            .WCLK(N__65615),
            .WE(N__39350));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_15,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_14,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_13,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_12,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_11,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_10,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_9,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_8,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_7,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_6,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_5,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_4,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_3,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_2,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_1,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_0}),
            .RADDR({dangling_wire_130,dangling_wire_131,dangling_wire_132,dangling_wire_133,dangling_wire_134,N__24788,N__24983,N__25160,N__25364,N__36092,N__25262}),
            .WADDR({dangling_wire_135,dangling_wire_136,dangling_wire_137,dangling_wire_138,dangling_wire_139,N__24779,N__24980,N__25157,N__25361,N__36089,N__25259}),
            .MASK({dangling_wire_140,dangling_wire_141,dangling_wire_142,dangling_wire_143,dangling_wire_144,dangling_wire_145,dangling_wire_146,dangling_wire_147,dangling_wire_148,dangling_wire_149,dangling_wire_150,dangling_wire_151,dangling_wire_152,dangling_wire_153,dangling_wire_154,dangling_wire_155}),
            .WDATA({N__23920,N__23961,N__23998,N__24033,N__24491,N__24698,N__24274,N__26182,N__34001,N__26380,N__24349,N__24387,N__23794,N__24620,N__23659,N__23698}),
            .RCLKE(),
            .RCLK(N__65544),
            .RE(N__39392),
            .WCLKE(N__26637),
            .WCLK(N__65545),
            .WE(N__39381));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_15,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_14,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_13,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_12,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_11,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_10,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_9,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_8,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_7,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_6,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_5,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_4,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_3,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_2,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_1,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_0}),
            .RADDR({dangling_wire_156,dangling_wire_157,dangling_wire_158,dangling_wire_159,dangling_wire_160,N__24764,N__24959,N__25136,N__25340,N__36068,N__25238}),
            .WADDR({dangling_wire_161,dangling_wire_162,dangling_wire_163,dangling_wire_164,dangling_wire_165,N__24755,N__24956,N__25133,N__25337,N__36065,N__25235}),
            .MASK({dangling_wire_166,dangling_wire_167,dangling_wire_168,dangling_wire_169,dangling_wire_170,dangling_wire_171,dangling_wire_172,dangling_wire_173,dangling_wire_174,dangling_wire_175,dangling_wire_176,dangling_wire_177,dangling_wire_178,dangling_wire_179,dangling_wire_180,dangling_wire_181}),
            .WDATA({N__23913,N__23962,N__23991,N__24037,N__24484,N__24679,N__24255,N__26169,N__33994,N__26376,N__24345,N__24391,N__23790,N__24601,N__23677,N__23716}),
            .RCLKE(),
            .RCLK(N__65594),
            .RE(N__39362),
            .WCLKE(N__24548),
            .WCLK(N__65593),
            .WE(N__39373));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical .WRITE_MODE=0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical .READ_MODE=0;
    SB_RAM40_4K \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical  (
            .RDATA({cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_31,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_30,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_29,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_28,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_27,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_26,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_25,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_24,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_23,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_22,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_21,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_20,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_19,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_18,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_17,cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_16}),
            .RADDR({dangling_wire_182,dangling_wire_183,dangling_wire_184,dangling_wire_185,dangling_wire_186,N__24776,N__24971,N__25148,N__25352,N__36080,N__25250}),
            .WADDR({dangling_wire_187,dangling_wire_188,dangling_wire_189,dangling_wire_190,dangling_wire_191,N__24767,N__24968,N__25145,N__25349,N__36077,N__25247}),
            .MASK({dangling_wire_192,dangling_wire_193,dangling_wire_194,dangling_wire_195,dangling_wire_196,dangling_wire_197,dangling_wire_198,dangling_wire_199,dangling_wire_200,dangling_wire_201,dangling_wire_202,dangling_wire_203,dangling_wire_204,dangling_wire_205,dangling_wire_206,dangling_wire_207}),
            .WDATA({N__26538,N__24657,N__24073,N__24452,N__24532,N__24154,N__24231,N__24583,N__24189,N__24292,N__24118,N__23818,N__26412,N__26457,N__26502,N__23860}),
            .RCLKE(),
            .RCLK(N__65569),
            .RE(N__39382),
            .WCLKE(N__26636),
            .WCLK(N__65570),
            .WE(N__39374));
    IO_PAD next_sequence_obuf_iopad (
            .OE(N__67138),
            .DIN(N__67137),
            .DOUT(N__67136),
            .PACKAGEPIN(next_sequence));
    defparam next_sequence_obuf_preio.NEG_TRIGGER=1'b0;
    defparam next_sequence_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO next_sequence_obuf_preio (
            .PADOEN(N__67138),
            .PADOUT(N__67137),
            .PADIN(N__67136),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__31524),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD stop_fpga2_obuf_iopad (
            .OE(N__67129),
            .DIN(N__67128),
            .DOUT(N__67127),
            .PACKAGEPIN(stop_fpga2));
    defparam stop_fpga2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam stop_fpga2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO stop_fpga2_obuf_preio (
            .PADOEN(N__67129),
            .PADOUT(N__67128),
            .PADIN(N__67127),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__33015),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD stop1_obuf_iopad (
            .OE(N__67120),
            .DIN(N__67119),
            .DOUT(N__67118),
            .PACKAGEPIN(stop1));
    defparam stop1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam stop1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO stop1_obuf_preio (
            .PADOEN(N__67120),
            .PADOUT(N__67119),
            .PADIN(N__67118),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s0_obuf_iopad (
            .OE(N__67111),
            .DIN(N__67110),
            .DOUT(N__67109),
            .PACKAGEPIN(s0));
    defparam s0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s0_obuf_preio (
            .PADOEN(N__67111),
            .PADOUT(N__67110),
            .PADIN(N__67109),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD mcu_data_obuf_iopad (
            .OE(N__67102),
            .DIN(N__67101),
            .DOUT(N__67100),
            .PACKAGEPIN(mcu_data));
    defparam mcu_data_obuf_preio.NEG_TRIGGER=1'b0;
    defparam mcu_data_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO mcu_data_obuf_preio (
            .PADOEN(N__67102),
            .PADOUT(N__67101),
            .PADIN(N__67100),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22536),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start1_obuf_iopad (
            .OE(N__67093),
            .DIN(N__67092),
            .DOUT(N__67091),
            .PACKAGEPIN(start1));
    defparam start1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam start1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO start1_obuf_preio (
            .PADOEN(N__67093),
            .PADOUT(N__67092),
            .PADIN(N__67091),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD rst_n_ibuf_iopad (
            .OE(N__67084),
            .DIN(N__67083),
            .DOUT(N__67082),
            .PACKAGEPIN(rst_n));
    defparam rst_n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam rst_n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO rst_n_ibuf_preio (
            .PADOEN(N__67084),
            .PADOUT(N__67083),
            .PADIN(N__67082),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(rst_n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD scl_ibuf_iopad (
            .OE(N__67075),
            .DIN(N__67074),
            .DOUT(N__67073),
            .PACKAGEPIN(scl));
    defparam scl_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam scl_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO scl_ibuf_preio (
            .PADOEN(N__67075),
            .PADOUT(N__67074),
            .PADIN(N__67073),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(scl_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout0_obuf_iopad (
            .OE(N__67066),
            .DIN(N__67065),
            .DOUT(N__67064),
            .PACKAGEPIN(dout0));
    defparam dout0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam dout0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO dout0_obuf_preio (
            .PADOEN(N__67066),
            .PADOUT(N__67065),
            .PADIN(N__67064),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23139),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD stop0_obuf_iopad (
            .OE(N__67057),
            .DIN(N__67056),
            .DOUT(N__67055),
            .PACKAGEPIN(stop0));
    defparam stop0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam stop0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO stop0_obuf_preio (
            .PADOEN(N__67057),
            .PADOUT(N__67056),
            .PADIN(N__67055),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s2_obuf_iopad (
            .OE(N__67048),
            .DIN(N__67047),
            .DOUT(N__67046),
            .PACKAGEPIN(s2));
    defparam s2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s2_obuf_preio (
            .PADOEN(N__67048),
            .PADOUT(N__67047),
            .PADIN(N__67046),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24840),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD mcu_sclk_obuf_iopad (
            .OE(N__67039),
            .DIN(N__67038),
            .DOUT(N__67037),
            .PACKAGEPIN(mcu_sclk));
    defparam mcu_sclk_obuf_preio.NEG_TRIGGER=1'b0;
    defparam mcu_sclk_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO mcu_sclk_obuf_preio (
            .PADOEN(N__67039),
            .PADOUT(N__67038),
            .PADIN(N__67037),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22359),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD frame_sync_obuf_iopad (
            .OE(N__67030),
            .DIN(N__67029),
            .DOUT(N__67028),
            .PACKAGEPIN(frame_sync));
    defparam frame_sync_obuf_preio.NEG_TRIGGER=1'b0;
    defparam frame_sync_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO frame_sync_obuf_preio (
            .PADOEN(N__67030),
            .PADOUT(N__67029),
            .PADIN(N__67028),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sdin0_ibuf_iopad (
            .OE(N__67021),
            .DIN(N__67020),
            .DOUT(N__67019),
            .PACKAGEPIN(sdin0));
    defparam sdin0_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam sdin0_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO sdin0_ibuf_preio (
            .PADOEN(N__67021),
            .PADOUT(N__67020),
            .PADIN(N__67019),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sdin0_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sdin1_ibuf_iopad (
            .OE(N__67012),
            .DIN(N__67011),
            .DOUT(N__67010),
            .PACKAGEPIN(sdin1));
    defparam sdin1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam sdin1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO sdin1_ibuf_preio (
            .PADOEN(N__67012),
            .PADOUT(N__67011),
            .PADIN(N__67010),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sdin1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD dout1_obuf_iopad (
            .OE(N__67003),
            .DIN(N__67002),
            .DOUT(N__67001),
            .PACKAGEPIN(dout1));
    defparam dout1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam dout1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO dout1_obuf_preio (
            .PADOEN(N__67003),
            .PADOUT(N__67002),
            .PADIN(N__67001),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23265),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD csb1_obuf_iopad (
            .OE(N__66994),
            .DIN(N__66993),
            .DOUT(N__66992),
            .PACKAGEPIN(csb1));
    defparam csb1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam csb1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO csb1_obuf_preio (
            .PADOEN(N__66994),
            .PADOUT(N__66993),
            .PADIN(N__66992),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__25653),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sclk1_obuf_iopad (
            .OE(N__66985),
            .DIN(N__66984),
            .DOUT(N__66983),
            .PACKAGEPIN(sclk1));
    defparam sclk1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sclk1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sclk1_obuf_preio (
            .PADOEN(N__66985),
            .PADOUT(N__66984),
            .PADIN(N__66983),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22899),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sclk0_obuf_iopad (
            .OE(N__66976),
            .DIN(N__66975),
            .DOUT(N__66974),
            .PACKAGEPIN(sclk0));
    defparam sclk0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam sclk0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO sclk0_obuf_preio (
            .PADOEN(N__66976),
            .PADOUT(N__66975),
            .PADIN(N__66974),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__22593),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s1_obuf_iopad (
            .OE(N__66967),
            .DIN(N__66966),
            .DOUT(N__66965),
            .PACKAGEPIN(s1));
    defparam s1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s1_obuf_preio (
            .PADOEN(N__66967),
            .PADOUT(N__66966),
            .PADIN(N__66965),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__24836),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD enable_config_obuf_iopad (
            .OE(N__66958),
            .DIN(N__66957),
            .DOUT(N__66956),
            .PACKAGEPIN(enable_config));
    defparam enable_config_obuf_preio.NEG_TRIGGER=1'b0;
    defparam enable_config_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO enable_config_obuf_preio (
            .PADOEN(N__66958),
            .PADOUT(N__66957),
            .PADIN(N__66956),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37449),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD sync_50hz_ibuf_iopad (
            .OE(N__66949),
            .DIN(N__66948),
            .DOUT(N__66947),
            .PACKAGEPIN(sync_50hz));
    defparam sync_50hz_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam sync_50hz_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO sync_50hz_ibuf_preio (
            .PADOEN(N__66949),
            .PADOUT(N__66948),
            .PADIN(N__66947),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(sync_50hz_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD serial_out_testing_obuf_iopad (
            .OE(N__66940),
            .DIN(N__66939),
            .DOUT(N__66938),
            .PACKAGEPIN(serial_out_testing));
    defparam serial_out_testing_obuf_preio.NEG_TRIGGER=1'b0;
    defparam serial_out_testing_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO serial_out_testing_obuf_preio (
            .PADOEN(N__66940),
            .PADOUT(N__66939),
            .PADIN(N__66938),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__35508),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD start0_obuf_iopad (
            .OE(N__66931),
            .DIN(N__66930),
            .DOUT(N__66929),
            .PACKAGEPIN(start0));
    defparam start0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam start0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO start0_obuf_preio (
            .PADOEN(N__66931),
            .PADOUT(N__66930),
            .PADIN(N__66929),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD s3_obuf_iopad (
            .OE(N__66922),
            .DIN(N__66921),
            .DOUT(N__66920),
            .PACKAGEPIN(s3));
    defparam s3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam s3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO s3_obuf_preio (
            .PADOEN(N__66922),
            .PADOUT(N__66921),
            .PADIN(N__66920),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD elec_config_out_obuf_iopad (
            .OE(N__66913),
            .DIN(N__66912),
            .DOUT(N__66911),
            .PACKAGEPIN(elec_config_out));
    defparam elec_config_out_obuf_preio.NEG_TRIGGER=1'b0;
    defparam elec_config_out_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO elec_config_out_obuf_preio (
            .PADOEN(N__66913),
            .PADOUT(N__66912),
            .PADIN(N__66911),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__37437),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD csb0_obuf_iopad (
            .OE(N__66904),
            .DIN(N__66903),
            .DOUT(N__66902),
            .PACKAGEPIN(csb0));
    defparam csb0_obuf_preio.NEG_TRIGGER=1'b0;
    defparam csb0_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO csb0_obuf_preio (
            .PADOEN(N__66904),
            .PADOUT(N__66903),
            .PADIN(N__66902),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__23064),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam IO_PIN_INST_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD IO_PIN_INST_iopad (
            .OE(N__66895),
            .DIN(N__66894),
            .DOUT(N__66893),
            .PACKAGEPIN(sda));
    defparam IO_PIN_INST_preio.PIN_TYPE=6'b101001;
    defparam IO_PIN_INST_preio.NEG_TRIGGER=1'b0;
    PRE_IO IO_PIN_INST_preio (
            .PADOEN(N__66895),
            .PADOUT(N__66894),
            .PADIN(N__66893),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(N__29340),
            .DIN0(s_sda_i),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD clock_ibuf_gb_io_iopad (
            .OE(N__66886),
            .DIN(N__66885),
            .DOUT(N__66884),
            .PACKAGEPIN(clock));
    defparam clock_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clock_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clock_ibuf_gb_io_preio (
            .PADOEN(N__66886),
            .PADOUT(N__66885),
            .PADIN(N__66884),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clock_ibuf_gb_io_gb_input),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__16711 (
            .O(N__66867),
            .I(N__66863));
    InMux I__16710 (
            .O(N__66866),
            .I(N__66860));
    LocalMux I__16709 (
            .O(N__66863),
            .I(N__66857));
    LocalMux I__16708 (
            .O(N__66860),
            .I(N__66854));
    Span4Mux_h I__16707 (
            .O(N__66857),
            .I(N__66847));
    Span4Mux_v I__16706 (
            .O(N__66854),
            .I(N__66844));
    InMux I__16705 (
            .O(N__66853),
            .I(N__66839));
    InMux I__16704 (
            .O(N__66852),
            .I(N__66839));
    InMux I__16703 (
            .O(N__66851),
            .I(N__66834));
    InMux I__16702 (
            .O(N__66850),
            .I(N__66834));
    Odrv4 I__16701 (
            .O(N__66847),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0 ));
    Odrv4 I__16700 (
            .O(N__66844),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0 ));
    LocalMux I__16699 (
            .O(N__66839),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0 ));
    LocalMux I__16698 (
            .O(N__66834),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0 ));
    CascadeMux I__16697 (
            .O(N__66825),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0_cascade_ ));
    CascadeMux I__16696 (
            .O(N__66822),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_0_2_cascade_ ));
    CascadeMux I__16695 (
            .O(N__66819),
            .I(N__66816));
    InMux I__16694 (
            .O(N__66816),
            .I(N__66806));
    InMux I__16693 (
            .O(N__66815),
            .I(N__66806));
    InMux I__16692 (
            .O(N__66814),
            .I(N__66806));
    CascadeMux I__16691 (
            .O(N__66813),
            .I(N__66803));
    LocalMux I__16690 (
            .O(N__66806),
            .I(N__66800));
    InMux I__16689 (
            .O(N__66803),
            .I(N__66795));
    Span4Mux_v I__16688 (
            .O(N__66800),
            .I(N__66791));
    InMux I__16687 (
            .O(N__66799),
            .I(N__66784));
    InMux I__16686 (
            .O(N__66798),
            .I(N__66781));
    LocalMux I__16685 (
            .O(N__66795),
            .I(N__66776));
    InMux I__16684 (
            .O(N__66794),
            .I(N__66773));
    Span4Mux_v I__16683 (
            .O(N__66791),
            .I(N__66770));
    InMux I__16682 (
            .O(N__66790),
            .I(N__66764));
    InMux I__16681 (
            .O(N__66789),
            .I(N__66764));
    InMux I__16680 (
            .O(N__66788),
            .I(N__66759));
    InMux I__16679 (
            .O(N__66787),
            .I(N__66759));
    LocalMux I__16678 (
            .O(N__66784),
            .I(N__66756));
    LocalMux I__16677 (
            .O(N__66781),
            .I(N__66752));
    InMux I__16676 (
            .O(N__66780),
            .I(N__66747));
    InMux I__16675 (
            .O(N__66779),
            .I(N__66747));
    Span4Mux_v I__16674 (
            .O(N__66776),
            .I(N__66744));
    LocalMux I__16673 (
            .O(N__66773),
            .I(N__66739));
    Span4Mux_h I__16672 (
            .O(N__66770),
            .I(N__66739));
    InMux I__16671 (
            .O(N__66769),
            .I(N__66736));
    LocalMux I__16670 (
            .O(N__66764),
            .I(N__66731));
    LocalMux I__16669 (
            .O(N__66759),
            .I(N__66731));
    Span4Mux_h I__16668 (
            .O(N__66756),
            .I(N__66728));
    InMux I__16667 (
            .O(N__66755),
            .I(N__66725));
    Span4Mux_h I__16666 (
            .O(N__66752),
            .I(N__66720));
    LocalMux I__16665 (
            .O(N__66747),
            .I(N__66720));
    Span4Mux_h I__16664 (
            .O(N__66744),
            .I(N__66715));
    Span4Mux_h I__16663 (
            .O(N__66739),
            .I(N__66715));
    LocalMux I__16662 (
            .O(N__66736),
            .I(N__66708));
    Span4Mux_v I__16661 (
            .O(N__66731),
            .I(N__66708));
    Span4Mux_v I__16660 (
            .O(N__66728),
            .I(N__66708));
    LocalMux I__16659 (
            .O(N__66725),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8 ));
    Odrv4 I__16658 (
            .O(N__66720),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8 ));
    Odrv4 I__16657 (
            .O(N__66715),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8 ));
    Odrv4 I__16656 (
            .O(N__66708),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8 ));
    InMux I__16655 (
            .O(N__66699),
            .I(N__66696));
    LocalMux I__16654 (
            .O(N__66696),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_2 ));
    CascadeMux I__16653 (
            .O(N__66693),
            .I(N__66688));
    InMux I__16652 (
            .O(N__66692),
            .I(N__66684));
    InMux I__16651 (
            .O(N__66691),
            .I(N__66681));
    InMux I__16650 (
            .O(N__66688),
            .I(N__66677));
    InMux I__16649 (
            .O(N__66687),
            .I(N__66670));
    LocalMux I__16648 (
            .O(N__66684),
            .I(N__66665));
    LocalMux I__16647 (
            .O(N__66681),
            .I(N__66665));
    InMux I__16646 (
            .O(N__66680),
            .I(N__66662));
    LocalMux I__16645 (
            .O(N__66677),
            .I(N__66659));
    CascadeMux I__16644 (
            .O(N__66676),
            .I(N__66655));
    InMux I__16643 (
            .O(N__66675),
            .I(N__66650));
    InMux I__16642 (
            .O(N__66674),
            .I(N__66645));
    InMux I__16641 (
            .O(N__66673),
            .I(N__66645));
    LocalMux I__16640 (
            .O(N__66670),
            .I(N__66640));
    Span4Mux_v I__16639 (
            .O(N__66665),
            .I(N__66640));
    LocalMux I__16638 (
            .O(N__66662),
            .I(N__66637));
    Span4Mux_h I__16637 (
            .O(N__66659),
            .I(N__66634));
    InMux I__16636 (
            .O(N__66658),
            .I(N__66627));
    InMux I__16635 (
            .O(N__66655),
            .I(N__66627));
    InMux I__16634 (
            .O(N__66654),
            .I(N__66627));
    InMux I__16633 (
            .O(N__66653),
            .I(N__66624));
    LocalMux I__16632 (
            .O(N__66650),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    LocalMux I__16631 (
            .O(N__66645),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    Odrv4 I__16630 (
            .O(N__66640),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    Odrv12 I__16629 (
            .O(N__66637),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    Odrv4 I__16628 (
            .O(N__66634),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    LocalMux I__16627 (
            .O(N__66627),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    LocalMux I__16626 (
            .O(N__66624),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ));
    CascadeMux I__16625 (
            .O(N__66609),
            .I(N__66604));
    InMux I__16624 (
            .O(N__66608),
            .I(N__66599));
    InMux I__16623 (
            .O(N__66607),
            .I(N__66594));
    InMux I__16622 (
            .O(N__66604),
            .I(N__66594));
    InMux I__16621 (
            .O(N__66603),
            .I(N__66590));
    InMux I__16620 (
            .O(N__66602),
            .I(N__66587));
    LocalMux I__16619 (
            .O(N__66599),
            .I(N__66582));
    LocalMux I__16618 (
            .O(N__66594),
            .I(N__66582));
    InMux I__16617 (
            .O(N__66593),
            .I(N__66579));
    LocalMux I__16616 (
            .O(N__66590),
            .I(N__66574));
    LocalMux I__16615 (
            .O(N__66587),
            .I(N__66574));
    Span4Mux_h I__16614 (
            .O(N__66582),
            .I(N__66571));
    LocalMux I__16613 (
            .O(N__66579),
            .I(N__66568));
    Odrv4 I__16612 (
            .O(N__66574),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0 ));
    Odrv4 I__16611 (
            .O(N__66571),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0 ));
    Odrv12 I__16610 (
            .O(N__66568),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0 ));
    InMux I__16609 (
            .O(N__66561),
            .I(N__66556));
    InMux I__16608 (
            .O(N__66560),
            .I(N__66545));
    InMux I__16607 (
            .O(N__66559),
            .I(N__66542));
    LocalMux I__16606 (
            .O(N__66556),
            .I(N__66539));
    InMux I__16605 (
            .O(N__66555),
            .I(N__66536));
    InMux I__16604 (
            .O(N__66554),
            .I(N__66533));
    InMux I__16603 (
            .O(N__66553),
            .I(N__66522));
    InMux I__16602 (
            .O(N__66552),
            .I(N__66522));
    InMux I__16601 (
            .O(N__66551),
            .I(N__66522));
    InMux I__16600 (
            .O(N__66550),
            .I(N__66522));
    InMux I__16599 (
            .O(N__66549),
            .I(N__66522));
    InMux I__16598 (
            .O(N__66548),
            .I(N__66519));
    LocalMux I__16597 (
            .O(N__66545),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    LocalMux I__16596 (
            .O(N__66542),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    Odrv4 I__16595 (
            .O(N__66539),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    LocalMux I__16594 (
            .O(N__66536),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    LocalMux I__16593 (
            .O(N__66533),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    LocalMux I__16592 (
            .O(N__66522),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    LocalMux I__16591 (
            .O(N__66519),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ));
    InMux I__16590 (
            .O(N__66504),
            .I(N__66499));
    InMux I__16589 (
            .O(N__66503),
            .I(N__66489));
    InMux I__16588 (
            .O(N__66502),
            .I(N__66486));
    LocalMux I__16587 (
            .O(N__66499),
            .I(N__66483));
    InMux I__16586 (
            .O(N__66498),
            .I(N__66478));
    InMux I__16585 (
            .O(N__66497),
            .I(N__66478));
    InMux I__16584 (
            .O(N__66496),
            .I(N__66471));
    InMux I__16583 (
            .O(N__66495),
            .I(N__66471));
    InMux I__16582 (
            .O(N__66494),
            .I(N__66471));
    InMux I__16581 (
            .O(N__66493),
            .I(N__66466));
    InMux I__16580 (
            .O(N__66492),
            .I(N__66466));
    LocalMux I__16579 (
            .O(N__66489),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ));
    LocalMux I__16578 (
            .O(N__66486),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ));
    Odrv4 I__16577 (
            .O(N__66483),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ));
    LocalMux I__16576 (
            .O(N__66478),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ));
    LocalMux I__16575 (
            .O(N__66471),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ));
    LocalMux I__16574 (
            .O(N__66466),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ));
    InMux I__16573 (
            .O(N__66453),
            .I(N__66450));
    LocalMux I__16572 (
            .O(N__66450),
            .I(N__66446));
    CascadeMux I__16571 (
            .O(N__66449),
            .I(N__66443));
    Span4Mux_v I__16570 (
            .O(N__66446),
            .I(N__66440));
    InMux I__16569 (
            .O(N__66443),
            .I(N__66437));
    Span4Mux_v I__16568 (
            .O(N__66440),
            .I(N__66432));
    LocalMux I__16567 (
            .O(N__66437),
            .I(N__66432));
    Span4Mux_v I__16566 (
            .O(N__66432),
            .I(N__66428));
    InMux I__16565 (
            .O(N__66431),
            .I(N__66425));
    Odrv4 I__16564 (
            .O(N__66428),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0 ));
    LocalMux I__16563 (
            .O(N__66425),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0 ));
    InMux I__16562 (
            .O(N__66420),
            .I(N__66416));
    CascadeMux I__16561 (
            .O(N__66419),
            .I(N__66413));
    LocalMux I__16560 (
            .O(N__66416),
            .I(N__66407));
    InMux I__16559 (
            .O(N__66413),
            .I(N__66402));
    InMux I__16558 (
            .O(N__66412),
            .I(N__66402));
    InMux I__16557 (
            .O(N__66411),
            .I(N__66397));
    InMux I__16556 (
            .O(N__66410),
            .I(N__66397));
    Span4Mux_v I__16555 (
            .O(N__66407),
            .I(N__66394));
    LocalMux I__16554 (
            .O(N__66402),
            .I(N__66389));
    LocalMux I__16553 (
            .O(N__66397),
            .I(N__66389));
    Odrv4 I__16552 (
            .O(N__66394),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0 ));
    Odrv4 I__16551 (
            .O(N__66389),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0 ));
    InMux I__16550 (
            .O(N__66384),
            .I(N__66379));
    InMux I__16549 (
            .O(N__66383),
            .I(N__66370));
    InMux I__16548 (
            .O(N__66382),
            .I(N__66370));
    LocalMux I__16547 (
            .O(N__66379),
            .I(N__66367));
    InMux I__16546 (
            .O(N__66378),
            .I(N__66364));
    InMux I__16545 (
            .O(N__66377),
            .I(N__66361));
    InMux I__16544 (
            .O(N__66376),
            .I(N__66356));
    InMux I__16543 (
            .O(N__66375),
            .I(N__66356));
    LocalMux I__16542 (
            .O(N__66370),
            .I(N__66353));
    Span4Mux_h I__16541 (
            .O(N__66367),
            .I(N__66346));
    LocalMux I__16540 (
            .O(N__66364),
            .I(N__66346));
    LocalMux I__16539 (
            .O(N__66361),
            .I(N__66346));
    LocalMux I__16538 (
            .O(N__66356),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0 ));
    Odrv12 I__16537 (
            .O(N__66353),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0 ));
    Odrv4 I__16536 (
            .O(N__66346),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0 ));
    InMux I__16535 (
            .O(N__66339),
            .I(N__66336));
    LocalMux I__16534 (
            .O(N__66336),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1666_2 ));
    CascadeMux I__16533 (
            .O(N__66333),
            .I(N__66330));
    InMux I__16532 (
            .O(N__66330),
            .I(N__66321));
    InMux I__16531 (
            .O(N__66329),
            .I(N__66312));
    InMux I__16530 (
            .O(N__66328),
            .I(N__66312));
    InMux I__16529 (
            .O(N__66327),
            .I(N__66312));
    InMux I__16528 (
            .O(N__66326),
            .I(N__66312));
    InMux I__16527 (
            .O(N__66325),
            .I(N__66309));
    InMux I__16526 (
            .O(N__66324),
            .I(N__66306));
    LocalMux I__16525 (
            .O(N__66321),
            .I(N__66303));
    LocalMux I__16524 (
            .O(N__66312),
            .I(N__66300));
    LocalMux I__16523 (
            .O(N__66309),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17 ));
    LocalMux I__16522 (
            .O(N__66306),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17 ));
    Odrv12 I__16521 (
            .O(N__66303),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17 ));
    Odrv4 I__16520 (
            .O(N__66300),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17 ));
    InMux I__16519 (
            .O(N__66291),
            .I(N__66287));
    InMux I__16518 (
            .O(N__66290),
            .I(N__66284));
    LocalMux I__16517 (
            .O(N__66287),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_295 ));
    LocalMux I__16516 (
            .O(N__66284),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_295 ));
    CascadeMux I__16515 (
            .O(N__66279),
            .I(N_73_i_0_cascade_));
    InMux I__16514 (
            .O(N__66276),
            .I(N__66268));
    InMux I__16513 (
            .O(N__66275),
            .I(N__66268));
    InMux I__16512 (
            .O(N__66274),
            .I(N__66265));
    InMux I__16511 (
            .O(N__66273),
            .I(N__66261));
    LocalMux I__16510 (
            .O(N__66268),
            .I(N__66256));
    LocalMux I__16509 (
            .O(N__66265),
            .I(N__66256));
    InMux I__16508 (
            .O(N__66264),
            .I(N__66252));
    LocalMux I__16507 (
            .O(N__66261),
            .I(N__66248));
    Span4Mux_v I__16506 (
            .O(N__66256),
            .I(N__66245));
    InMux I__16505 (
            .O(N__66255),
            .I(N__66240));
    LocalMux I__16504 (
            .O(N__66252),
            .I(N__66237));
    InMux I__16503 (
            .O(N__66251),
            .I(N__66234));
    Span4Mux_v I__16502 (
            .O(N__66248),
            .I(N__66229));
    Span4Mux_h I__16501 (
            .O(N__66245),
            .I(N__66229));
    InMux I__16500 (
            .O(N__66244),
            .I(N__66226));
    InMux I__16499 (
            .O(N__66243),
            .I(N__66223));
    LocalMux I__16498 (
            .O(N__66240),
            .I(N__66220));
    Span4Mux_h I__16497 (
            .O(N__66237),
            .I(N__66215));
    LocalMux I__16496 (
            .O(N__66234),
            .I(N__66215));
    Span4Mux_h I__16495 (
            .O(N__66229),
            .I(N__66210));
    LocalMux I__16494 (
            .O(N__66226),
            .I(N__66210));
    LocalMux I__16493 (
            .O(N__66223),
            .I(I2C_top_level_inst1_s_burst));
    Odrv12 I__16492 (
            .O(N__66220),
            .I(I2C_top_level_inst1_s_burst));
    Odrv4 I__16491 (
            .O(N__66215),
            .I(I2C_top_level_inst1_s_burst));
    Odrv4 I__16490 (
            .O(N__66210),
            .I(I2C_top_level_inst1_s_burst));
    InMux I__16489 (
            .O(N__66201),
            .I(N__66198));
    LocalMux I__16488 (
            .O(N__66198),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_19 ));
    CascadeMux I__16487 (
            .O(N__66195),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_274_cascade_ ));
    CascadeMux I__16486 (
            .O(N__66192),
            .I(N__66188));
    InMux I__16485 (
            .O(N__66191),
            .I(N__66175));
    InMux I__16484 (
            .O(N__66188),
            .I(N__66175));
    InMux I__16483 (
            .O(N__66187),
            .I(N__66175));
    InMux I__16482 (
            .O(N__66186),
            .I(N__66175));
    InMux I__16481 (
            .O(N__66185),
            .I(N__66169));
    InMux I__16480 (
            .O(N__66184),
            .I(N__66169));
    LocalMux I__16479 (
            .O(N__66175),
            .I(N__66160));
    InMux I__16478 (
            .O(N__66174),
            .I(N__66157));
    LocalMux I__16477 (
            .O(N__66169),
            .I(N__66151));
    InMux I__16476 (
            .O(N__66168),
            .I(N__66143));
    InMux I__16475 (
            .O(N__66167),
            .I(N__66143));
    InMux I__16474 (
            .O(N__66166),
            .I(N__66143));
    InMux I__16473 (
            .O(N__66165),
            .I(N__66138));
    InMux I__16472 (
            .O(N__66164),
            .I(N__66138));
    InMux I__16471 (
            .O(N__66163),
            .I(N__66135));
    Span4Mux_h I__16470 (
            .O(N__66160),
            .I(N__66130));
    LocalMux I__16469 (
            .O(N__66157),
            .I(N__66130));
    CascadeMux I__16468 (
            .O(N__66156),
            .I(N__66126));
    CascadeMux I__16467 (
            .O(N__66155),
            .I(N__66122));
    CascadeMux I__16466 (
            .O(N__66154),
            .I(N__66119));
    Span4Mux_v I__16465 (
            .O(N__66151),
            .I(N__66115));
    InMux I__16464 (
            .O(N__66150),
            .I(N__66112));
    LocalMux I__16463 (
            .O(N__66143),
            .I(N__66106));
    LocalMux I__16462 (
            .O(N__66138),
            .I(N__66102));
    LocalMux I__16461 (
            .O(N__66135),
            .I(N__66099));
    Span4Mux_h I__16460 (
            .O(N__66130),
            .I(N__66096));
    InMux I__16459 (
            .O(N__66129),
            .I(N__66086));
    InMux I__16458 (
            .O(N__66126),
            .I(N__66086));
    InMux I__16457 (
            .O(N__66125),
            .I(N__66086));
    InMux I__16456 (
            .O(N__66122),
            .I(N__66079));
    InMux I__16455 (
            .O(N__66119),
            .I(N__66079));
    InMux I__16454 (
            .O(N__66118),
            .I(N__66079));
    Span4Mux_v I__16453 (
            .O(N__66115),
            .I(N__66074));
    LocalMux I__16452 (
            .O(N__66112),
            .I(N__66074));
    InMux I__16451 (
            .O(N__66111),
            .I(N__66067));
    InMux I__16450 (
            .O(N__66110),
            .I(N__66067));
    InMux I__16449 (
            .O(N__66109),
            .I(N__66067));
    Span4Mux_v I__16448 (
            .O(N__66106),
            .I(N__66064));
    InMux I__16447 (
            .O(N__66105),
            .I(N__66061));
    Span4Mux_h I__16446 (
            .O(N__66102),
            .I(N__66054));
    Span4Mux_h I__16445 (
            .O(N__66099),
            .I(N__66054));
    Span4Mux_v I__16444 (
            .O(N__66096),
            .I(N__66054));
    InMux I__16443 (
            .O(N__66095),
            .I(N__66051));
    InMux I__16442 (
            .O(N__66094),
            .I(N__66046));
    InMux I__16441 (
            .O(N__66093),
            .I(N__66046));
    LocalMux I__16440 (
            .O(N__66086),
            .I(N__66041));
    LocalMux I__16439 (
            .O(N__66079),
            .I(N__66041));
    Span4Mux_h I__16438 (
            .O(N__66074),
            .I(N__66038));
    LocalMux I__16437 (
            .O(N__66067),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    Odrv4 I__16436 (
            .O(N__66064),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    LocalMux I__16435 (
            .O(N__66061),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    Odrv4 I__16434 (
            .O(N__66054),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    LocalMux I__16433 (
            .O(N__66051),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    LocalMux I__16432 (
            .O(N__66046),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    Odrv4 I__16431 (
            .O(N__66041),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    Odrv4 I__16430 (
            .O(N__66038),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2));
    InMux I__16429 (
            .O(N__66021),
            .I(N__66012));
    InMux I__16428 (
            .O(N__66020),
            .I(N__66012));
    InMux I__16427 (
            .O(N__66019),
            .I(N__66009));
    InMux I__16426 (
            .O(N__66018),
            .I(N__66006));
    InMux I__16425 (
            .O(N__66017),
            .I(N__66003));
    LocalMux I__16424 (
            .O(N__66012),
            .I(N__65998));
    LocalMux I__16423 (
            .O(N__66009),
            .I(N__65998));
    LocalMux I__16422 (
            .O(N__66006),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19 ));
    LocalMux I__16421 (
            .O(N__66003),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19 ));
    Odrv4 I__16420 (
            .O(N__65998),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19 ));
    InMux I__16419 (
            .O(N__65991),
            .I(N__65988));
    LocalMux I__16418 (
            .O(N__65988),
            .I(N__65982));
    CascadeMux I__16417 (
            .O(N__65987),
            .I(N__65979));
    CascadeMux I__16416 (
            .O(N__65986),
            .I(N__65975));
    InMux I__16415 (
            .O(N__65985),
            .I(N__65971));
    Span4Mux_v I__16414 (
            .O(N__65982),
            .I(N__65968));
    InMux I__16413 (
            .O(N__65979),
            .I(N__65965));
    InMux I__16412 (
            .O(N__65978),
            .I(N__65962));
    InMux I__16411 (
            .O(N__65975),
            .I(N__65957));
    InMux I__16410 (
            .O(N__65974),
            .I(N__65957));
    LocalMux I__16409 (
            .O(N__65971),
            .I(N__65946));
    Sp12to4 I__16408 (
            .O(N__65968),
            .I(N__65946));
    LocalMux I__16407 (
            .O(N__65965),
            .I(N__65946));
    LocalMux I__16406 (
            .O(N__65962),
            .I(N__65946));
    LocalMux I__16405 (
            .O(N__65957),
            .I(N__65946));
    Span12Mux_h I__16404 (
            .O(N__65946),
            .I(N__65942));
    InMux I__16403 (
            .O(N__65945),
            .I(N__65939));
    Odrv12 I__16402 (
            .O(N__65942),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6));
    LocalMux I__16401 (
            .O(N__65939),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6));
    InMux I__16400 (
            .O(N__65934),
            .I(N__65927));
    InMux I__16399 (
            .O(N__65933),
            .I(N__65927));
    CascadeMux I__16398 (
            .O(N__65932),
            .I(N__65923));
    LocalMux I__16397 (
            .O(N__65927),
            .I(N__65920));
    InMux I__16396 (
            .O(N__65926),
            .I(N__65915));
    InMux I__16395 (
            .O(N__65923),
            .I(N__65915));
    Span4Mux_h I__16394 (
            .O(N__65920),
            .I(N__65909));
    LocalMux I__16393 (
            .O(N__65915),
            .I(N__65909));
    InMux I__16392 (
            .O(N__65914),
            .I(N__65906));
    Span4Mux_h I__16391 (
            .O(N__65909),
            .I(N__65903));
    LocalMux I__16390 (
            .O(N__65906),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2 ));
    Odrv4 I__16389 (
            .O(N__65903),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2 ));
    CascadeMux I__16388 (
            .O(N__65898),
            .I(N__65894));
    InMux I__16387 (
            .O(N__65897),
            .I(N__65889));
    InMux I__16386 (
            .O(N__65894),
            .I(N__65884));
    InMux I__16385 (
            .O(N__65893),
            .I(N__65884));
    InMux I__16384 (
            .O(N__65892),
            .I(N__65881));
    LocalMux I__16383 (
            .O(N__65889),
            .I(N__65878));
    LocalMux I__16382 (
            .O(N__65884),
            .I(N__65873));
    LocalMux I__16381 (
            .O(N__65881),
            .I(N__65873));
    Span4Mux_v I__16380 (
            .O(N__65878),
            .I(N__65866));
    Span4Mux_v I__16379 (
            .O(N__65873),
            .I(N__65866));
    InMux I__16378 (
            .O(N__65872),
            .I(N__65861));
    InMux I__16377 (
            .O(N__65871),
            .I(N__65861));
    Odrv4 I__16376 (
            .O(N__65866),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2));
    LocalMux I__16375 (
            .O(N__65861),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2));
    InMux I__16374 (
            .O(N__65856),
            .I(N__65853));
    LocalMux I__16373 (
            .O(N__65853),
            .I(N__65849));
    InMux I__16372 (
            .O(N__65852),
            .I(N__65845));
    Span4Mux_v I__16371 (
            .O(N__65849),
            .I(N__65842));
    InMux I__16370 (
            .O(N__65848),
            .I(N__65839));
    LocalMux I__16369 (
            .O(N__65845),
            .I(N__65836));
    Odrv4 I__16368 (
            .O(N__65842),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2 ));
    LocalMux I__16367 (
            .O(N__65839),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2 ));
    Odrv4 I__16366 (
            .O(N__65836),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2 ));
    InMux I__16365 (
            .O(N__65829),
            .I(N__65826));
    LocalMux I__16364 (
            .O(N__65826),
            .I(N__65823));
    Odrv4 I__16363 (
            .O(N__65823),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_276 ));
    InMux I__16362 (
            .O(N__65820),
            .I(N__65816));
    InMux I__16361 (
            .O(N__65819),
            .I(N__65813));
    LocalMux I__16360 (
            .O(N__65816),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1 ));
    LocalMux I__16359 (
            .O(N__65813),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1 ));
    CascadeMux I__16358 (
            .O(N__65808),
            .I(N__65804));
    CascadeMux I__16357 (
            .O(N__65807),
            .I(N__65801));
    InMux I__16356 (
            .O(N__65804),
            .I(N__65797));
    InMux I__16355 (
            .O(N__65801),
            .I(N__65792));
    InMux I__16354 (
            .O(N__65800),
            .I(N__65792));
    LocalMux I__16353 (
            .O(N__65797),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_245 ));
    LocalMux I__16352 (
            .O(N__65792),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_245 ));
    InMux I__16351 (
            .O(N__65787),
            .I(N__65784));
    LocalMux I__16350 (
            .O(N__65784),
            .I(N__65780));
    InMux I__16349 (
            .O(N__65783),
            .I(N__65777));
    Odrv4 I__16348 (
            .O(N__65780),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0 ));
    LocalMux I__16347 (
            .O(N__65777),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0 ));
    CascadeMux I__16346 (
            .O(N__65772),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1669_cascade_ ));
    InMux I__16345 (
            .O(N__65769),
            .I(N__65764));
    InMux I__16344 (
            .O(N__65768),
            .I(N__65761));
    InMux I__16343 (
            .O(N__65767),
            .I(N__65758));
    LocalMux I__16342 (
            .O(N__65764),
            .I(N__65755));
    LocalMux I__16341 (
            .O(N__65761),
            .I(N__65710));
    LocalMux I__16340 (
            .O(N__65758),
            .I(N__65707));
    Glb2LocalMux I__16339 (
            .O(N__65755),
            .I(N__65034));
    ClkMux I__16338 (
            .O(N__65754),
            .I(N__65034));
    ClkMux I__16337 (
            .O(N__65753),
            .I(N__65034));
    ClkMux I__16336 (
            .O(N__65752),
            .I(N__65034));
    ClkMux I__16335 (
            .O(N__65751),
            .I(N__65034));
    ClkMux I__16334 (
            .O(N__65750),
            .I(N__65034));
    ClkMux I__16333 (
            .O(N__65749),
            .I(N__65034));
    ClkMux I__16332 (
            .O(N__65748),
            .I(N__65034));
    ClkMux I__16331 (
            .O(N__65747),
            .I(N__65034));
    ClkMux I__16330 (
            .O(N__65746),
            .I(N__65034));
    ClkMux I__16329 (
            .O(N__65745),
            .I(N__65034));
    ClkMux I__16328 (
            .O(N__65744),
            .I(N__65034));
    ClkMux I__16327 (
            .O(N__65743),
            .I(N__65034));
    ClkMux I__16326 (
            .O(N__65742),
            .I(N__65034));
    ClkMux I__16325 (
            .O(N__65741),
            .I(N__65034));
    ClkMux I__16324 (
            .O(N__65740),
            .I(N__65034));
    ClkMux I__16323 (
            .O(N__65739),
            .I(N__65034));
    ClkMux I__16322 (
            .O(N__65738),
            .I(N__65034));
    ClkMux I__16321 (
            .O(N__65737),
            .I(N__65034));
    ClkMux I__16320 (
            .O(N__65736),
            .I(N__65034));
    ClkMux I__16319 (
            .O(N__65735),
            .I(N__65034));
    ClkMux I__16318 (
            .O(N__65734),
            .I(N__65034));
    ClkMux I__16317 (
            .O(N__65733),
            .I(N__65034));
    ClkMux I__16316 (
            .O(N__65732),
            .I(N__65034));
    ClkMux I__16315 (
            .O(N__65731),
            .I(N__65034));
    ClkMux I__16314 (
            .O(N__65730),
            .I(N__65034));
    ClkMux I__16313 (
            .O(N__65729),
            .I(N__65034));
    ClkMux I__16312 (
            .O(N__65728),
            .I(N__65034));
    ClkMux I__16311 (
            .O(N__65727),
            .I(N__65034));
    ClkMux I__16310 (
            .O(N__65726),
            .I(N__65034));
    ClkMux I__16309 (
            .O(N__65725),
            .I(N__65034));
    ClkMux I__16308 (
            .O(N__65724),
            .I(N__65034));
    ClkMux I__16307 (
            .O(N__65723),
            .I(N__65034));
    ClkMux I__16306 (
            .O(N__65722),
            .I(N__65034));
    ClkMux I__16305 (
            .O(N__65721),
            .I(N__65034));
    ClkMux I__16304 (
            .O(N__65720),
            .I(N__65034));
    ClkMux I__16303 (
            .O(N__65719),
            .I(N__65034));
    ClkMux I__16302 (
            .O(N__65718),
            .I(N__65034));
    ClkMux I__16301 (
            .O(N__65717),
            .I(N__65034));
    ClkMux I__16300 (
            .O(N__65716),
            .I(N__65034));
    ClkMux I__16299 (
            .O(N__65715),
            .I(N__65034));
    ClkMux I__16298 (
            .O(N__65714),
            .I(N__65034));
    ClkMux I__16297 (
            .O(N__65713),
            .I(N__65034));
    Glb2LocalMux I__16296 (
            .O(N__65710),
            .I(N__65034));
    Glb2LocalMux I__16295 (
            .O(N__65707),
            .I(N__65034));
    ClkMux I__16294 (
            .O(N__65706),
            .I(N__65034));
    ClkMux I__16293 (
            .O(N__65705),
            .I(N__65034));
    ClkMux I__16292 (
            .O(N__65704),
            .I(N__65034));
    ClkMux I__16291 (
            .O(N__65703),
            .I(N__65034));
    ClkMux I__16290 (
            .O(N__65702),
            .I(N__65034));
    ClkMux I__16289 (
            .O(N__65701),
            .I(N__65034));
    ClkMux I__16288 (
            .O(N__65700),
            .I(N__65034));
    ClkMux I__16287 (
            .O(N__65699),
            .I(N__65034));
    ClkMux I__16286 (
            .O(N__65698),
            .I(N__65034));
    ClkMux I__16285 (
            .O(N__65697),
            .I(N__65034));
    ClkMux I__16284 (
            .O(N__65696),
            .I(N__65034));
    ClkMux I__16283 (
            .O(N__65695),
            .I(N__65034));
    ClkMux I__16282 (
            .O(N__65694),
            .I(N__65034));
    ClkMux I__16281 (
            .O(N__65693),
            .I(N__65034));
    ClkMux I__16280 (
            .O(N__65692),
            .I(N__65034));
    ClkMux I__16279 (
            .O(N__65691),
            .I(N__65034));
    ClkMux I__16278 (
            .O(N__65690),
            .I(N__65034));
    ClkMux I__16277 (
            .O(N__65689),
            .I(N__65034));
    ClkMux I__16276 (
            .O(N__65688),
            .I(N__65034));
    ClkMux I__16275 (
            .O(N__65687),
            .I(N__65034));
    ClkMux I__16274 (
            .O(N__65686),
            .I(N__65034));
    ClkMux I__16273 (
            .O(N__65685),
            .I(N__65034));
    ClkMux I__16272 (
            .O(N__65684),
            .I(N__65034));
    ClkMux I__16271 (
            .O(N__65683),
            .I(N__65034));
    ClkMux I__16270 (
            .O(N__65682),
            .I(N__65034));
    ClkMux I__16269 (
            .O(N__65681),
            .I(N__65034));
    ClkMux I__16268 (
            .O(N__65680),
            .I(N__65034));
    ClkMux I__16267 (
            .O(N__65679),
            .I(N__65034));
    ClkMux I__16266 (
            .O(N__65678),
            .I(N__65034));
    ClkMux I__16265 (
            .O(N__65677),
            .I(N__65034));
    ClkMux I__16264 (
            .O(N__65676),
            .I(N__65034));
    ClkMux I__16263 (
            .O(N__65675),
            .I(N__65034));
    ClkMux I__16262 (
            .O(N__65674),
            .I(N__65034));
    ClkMux I__16261 (
            .O(N__65673),
            .I(N__65034));
    ClkMux I__16260 (
            .O(N__65672),
            .I(N__65034));
    ClkMux I__16259 (
            .O(N__65671),
            .I(N__65034));
    ClkMux I__16258 (
            .O(N__65670),
            .I(N__65034));
    ClkMux I__16257 (
            .O(N__65669),
            .I(N__65034));
    ClkMux I__16256 (
            .O(N__65668),
            .I(N__65034));
    ClkMux I__16255 (
            .O(N__65667),
            .I(N__65034));
    ClkMux I__16254 (
            .O(N__65666),
            .I(N__65034));
    ClkMux I__16253 (
            .O(N__65665),
            .I(N__65034));
    ClkMux I__16252 (
            .O(N__65664),
            .I(N__65034));
    ClkMux I__16251 (
            .O(N__65663),
            .I(N__65034));
    ClkMux I__16250 (
            .O(N__65662),
            .I(N__65034));
    ClkMux I__16249 (
            .O(N__65661),
            .I(N__65034));
    ClkMux I__16248 (
            .O(N__65660),
            .I(N__65034));
    ClkMux I__16247 (
            .O(N__65659),
            .I(N__65034));
    ClkMux I__16246 (
            .O(N__65658),
            .I(N__65034));
    ClkMux I__16245 (
            .O(N__65657),
            .I(N__65034));
    ClkMux I__16244 (
            .O(N__65656),
            .I(N__65034));
    ClkMux I__16243 (
            .O(N__65655),
            .I(N__65034));
    ClkMux I__16242 (
            .O(N__65654),
            .I(N__65034));
    ClkMux I__16241 (
            .O(N__65653),
            .I(N__65034));
    ClkMux I__16240 (
            .O(N__65652),
            .I(N__65034));
    ClkMux I__16239 (
            .O(N__65651),
            .I(N__65034));
    ClkMux I__16238 (
            .O(N__65650),
            .I(N__65034));
    ClkMux I__16237 (
            .O(N__65649),
            .I(N__65034));
    ClkMux I__16236 (
            .O(N__65648),
            .I(N__65034));
    ClkMux I__16235 (
            .O(N__65647),
            .I(N__65034));
    ClkMux I__16234 (
            .O(N__65646),
            .I(N__65034));
    ClkMux I__16233 (
            .O(N__65645),
            .I(N__65034));
    ClkMux I__16232 (
            .O(N__65644),
            .I(N__65034));
    ClkMux I__16231 (
            .O(N__65643),
            .I(N__65034));
    ClkMux I__16230 (
            .O(N__65642),
            .I(N__65034));
    ClkMux I__16229 (
            .O(N__65641),
            .I(N__65034));
    ClkMux I__16228 (
            .O(N__65640),
            .I(N__65034));
    ClkMux I__16227 (
            .O(N__65639),
            .I(N__65034));
    ClkMux I__16226 (
            .O(N__65638),
            .I(N__65034));
    ClkMux I__16225 (
            .O(N__65637),
            .I(N__65034));
    ClkMux I__16224 (
            .O(N__65636),
            .I(N__65034));
    ClkMux I__16223 (
            .O(N__65635),
            .I(N__65034));
    ClkMux I__16222 (
            .O(N__65634),
            .I(N__65034));
    ClkMux I__16221 (
            .O(N__65633),
            .I(N__65034));
    ClkMux I__16220 (
            .O(N__65632),
            .I(N__65034));
    ClkMux I__16219 (
            .O(N__65631),
            .I(N__65034));
    ClkMux I__16218 (
            .O(N__65630),
            .I(N__65034));
    ClkMux I__16217 (
            .O(N__65629),
            .I(N__65034));
    ClkMux I__16216 (
            .O(N__65628),
            .I(N__65034));
    ClkMux I__16215 (
            .O(N__65627),
            .I(N__65034));
    ClkMux I__16214 (
            .O(N__65626),
            .I(N__65034));
    ClkMux I__16213 (
            .O(N__65625),
            .I(N__65034));
    ClkMux I__16212 (
            .O(N__65624),
            .I(N__65034));
    ClkMux I__16211 (
            .O(N__65623),
            .I(N__65034));
    ClkMux I__16210 (
            .O(N__65622),
            .I(N__65034));
    ClkMux I__16209 (
            .O(N__65621),
            .I(N__65034));
    ClkMux I__16208 (
            .O(N__65620),
            .I(N__65034));
    ClkMux I__16207 (
            .O(N__65619),
            .I(N__65034));
    ClkMux I__16206 (
            .O(N__65618),
            .I(N__65034));
    ClkMux I__16205 (
            .O(N__65617),
            .I(N__65034));
    ClkMux I__16204 (
            .O(N__65616),
            .I(N__65034));
    ClkMux I__16203 (
            .O(N__65615),
            .I(N__65034));
    ClkMux I__16202 (
            .O(N__65614),
            .I(N__65034));
    ClkMux I__16201 (
            .O(N__65613),
            .I(N__65034));
    ClkMux I__16200 (
            .O(N__65612),
            .I(N__65034));
    ClkMux I__16199 (
            .O(N__65611),
            .I(N__65034));
    ClkMux I__16198 (
            .O(N__65610),
            .I(N__65034));
    ClkMux I__16197 (
            .O(N__65609),
            .I(N__65034));
    ClkMux I__16196 (
            .O(N__65608),
            .I(N__65034));
    ClkMux I__16195 (
            .O(N__65607),
            .I(N__65034));
    ClkMux I__16194 (
            .O(N__65606),
            .I(N__65034));
    ClkMux I__16193 (
            .O(N__65605),
            .I(N__65034));
    ClkMux I__16192 (
            .O(N__65604),
            .I(N__65034));
    ClkMux I__16191 (
            .O(N__65603),
            .I(N__65034));
    ClkMux I__16190 (
            .O(N__65602),
            .I(N__65034));
    ClkMux I__16189 (
            .O(N__65601),
            .I(N__65034));
    ClkMux I__16188 (
            .O(N__65600),
            .I(N__65034));
    ClkMux I__16187 (
            .O(N__65599),
            .I(N__65034));
    ClkMux I__16186 (
            .O(N__65598),
            .I(N__65034));
    ClkMux I__16185 (
            .O(N__65597),
            .I(N__65034));
    ClkMux I__16184 (
            .O(N__65596),
            .I(N__65034));
    ClkMux I__16183 (
            .O(N__65595),
            .I(N__65034));
    ClkMux I__16182 (
            .O(N__65594),
            .I(N__65034));
    ClkMux I__16181 (
            .O(N__65593),
            .I(N__65034));
    ClkMux I__16180 (
            .O(N__65592),
            .I(N__65034));
    ClkMux I__16179 (
            .O(N__65591),
            .I(N__65034));
    ClkMux I__16178 (
            .O(N__65590),
            .I(N__65034));
    ClkMux I__16177 (
            .O(N__65589),
            .I(N__65034));
    ClkMux I__16176 (
            .O(N__65588),
            .I(N__65034));
    ClkMux I__16175 (
            .O(N__65587),
            .I(N__65034));
    ClkMux I__16174 (
            .O(N__65586),
            .I(N__65034));
    ClkMux I__16173 (
            .O(N__65585),
            .I(N__65034));
    ClkMux I__16172 (
            .O(N__65584),
            .I(N__65034));
    ClkMux I__16171 (
            .O(N__65583),
            .I(N__65034));
    ClkMux I__16170 (
            .O(N__65582),
            .I(N__65034));
    ClkMux I__16169 (
            .O(N__65581),
            .I(N__65034));
    ClkMux I__16168 (
            .O(N__65580),
            .I(N__65034));
    ClkMux I__16167 (
            .O(N__65579),
            .I(N__65034));
    ClkMux I__16166 (
            .O(N__65578),
            .I(N__65034));
    ClkMux I__16165 (
            .O(N__65577),
            .I(N__65034));
    ClkMux I__16164 (
            .O(N__65576),
            .I(N__65034));
    ClkMux I__16163 (
            .O(N__65575),
            .I(N__65034));
    ClkMux I__16162 (
            .O(N__65574),
            .I(N__65034));
    ClkMux I__16161 (
            .O(N__65573),
            .I(N__65034));
    ClkMux I__16160 (
            .O(N__65572),
            .I(N__65034));
    ClkMux I__16159 (
            .O(N__65571),
            .I(N__65034));
    ClkMux I__16158 (
            .O(N__65570),
            .I(N__65034));
    ClkMux I__16157 (
            .O(N__65569),
            .I(N__65034));
    ClkMux I__16156 (
            .O(N__65568),
            .I(N__65034));
    ClkMux I__16155 (
            .O(N__65567),
            .I(N__65034));
    ClkMux I__16154 (
            .O(N__65566),
            .I(N__65034));
    ClkMux I__16153 (
            .O(N__65565),
            .I(N__65034));
    ClkMux I__16152 (
            .O(N__65564),
            .I(N__65034));
    ClkMux I__16151 (
            .O(N__65563),
            .I(N__65034));
    ClkMux I__16150 (
            .O(N__65562),
            .I(N__65034));
    ClkMux I__16149 (
            .O(N__65561),
            .I(N__65034));
    ClkMux I__16148 (
            .O(N__65560),
            .I(N__65034));
    ClkMux I__16147 (
            .O(N__65559),
            .I(N__65034));
    ClkMux I__16146 (
            .O(N__65558),
            .I(N__65034));
    ClkMux I__16145 (
            .O(N__65557),
            .I(N__65034));
    ClkMux I__16144 (
            .O(N__65556),
            .I(N__65034));
    ClkMux I__16143 (
            .O(N__65555),
            .I(N__65034));
    ClkMux I__16142 (
            .O(N__65554),
            .I(N__65034));
    ClkMux I__16141 (
            .O(N__65553),
            .I(N__65034));
    ClkMux I__16140 (
            .O(N__65552),
            .I(N__65034));
    ClkMux I__16139 (
            .O(N__65551),
            .I(N__65034));
    ClkMux I__16138 (
            .O(N__65550),
            .I(N__65034));
    ClkMux I__16137 (
            .O(N__65549),
            .I(N__65034));
    ClkMux I__16136 (
            .O(N__65548),
            .I(N__65034));
    ClkMux I__16135 (
            .O(N__65547),
            .I(N__65034));
    ClkMux I__16134 (
            .O(N__65546),
            .I(N__65034));
    ClkMux I__16133 (
            .O(N__65545),
            .I(N__65034));
    ClkMux I__16132 (
            .O(N__65544),
            .I(N__65034));
    ClkMux I__16131 (
            .O(N__65543),
            .I(N__65034));
    ClkMux I__16130 (
            .O(N__65542),
            .I(N__65034));
    ClkMux I__16129 (
            .O(N__65541),
            .I(N__65034));
    ClkMux I__16128 (
            .O(N__65540),
            .I(N__65034));
    ClkMux I__16127 (
            .O(N__65539),
            .I(N__65034));
    ClkMux I__16126 (
            .O(N__65538),
            .I(N__65034));
    ClkMux I__16125 (
            .O(N__65537),
            .I(N__65034));
    ClkMux I__16124 (
            .O(N__65536),
            .I(N__65034));
    ClkMux I__16123 (
            .O(N__65535),
            .I(N__65034));
    ClkMux I__16122 (
            .O(N__65534),
            .I(N__65034));
    ClkMux I__16121 (
            .O(N__65533),
            .I(N__65034));
    ClkMux I__16120 (
            .O(N__65532),
            .I(N__65034));
    ClkMux I__16119 (
            .O(N__65531),
            .I(N__65034));
    ClkMux I__16118 (
            .O(N__65530),
            .I(N__65034));
    ClkMux I__16117 (
            .O(N__65529),
            .I(N__65034));
    ClkMux I__16116 (
            .O(N__65528),
            .I(N__65034));
    ClkMux I__16115 (
            .O(N__65527),
            .I(N__65034));
    ClkMux I__16114 (
            .O(N__65526),
            .I(N__65034));
    ClkMux I__16113 (
            .O(N__65525),
            .I(N__65034));
    ClkMux I__16112 (
            .O(N__65524),
            .I(N__65034));
    ClkMux I__16111 (
            .O(N__65523),
            .I(N__65034));
    ClkMux I__16110 (
            .O(N__65522),
            .I(N__65034));
    ClkMux I__16109 (
            .O(N__65521),
            .I(N__65034));
    ClkMux I__16108 (
            .O(N__65520),
            .I(N__65034));
    ClkMux I__16107 (
            .O(N__65519),
            .I(N__65034));
    ClkMux I__16106 (
            .O(N__65518),
            .I(N__65034));
    ClkMux I__16105 (
            .O(N__65517),
            .I(N__65034));
    ClkMux I__16104 (
            .O(N__65516),
            .I(N__65034));
    ClkMux I__16103 (
            .O(N__65515),
            .I(N__65034));
    ClkMux I__16102 (
            .O(N__65514),
            .I(N__65034));
    ClkMux I__16101 (
            .O(N__65513),
            .I(N__65034));
    GlobalMux I__16100 (
            .O(N__65034),
            .I(N__65031));
    gio2CtrlBuf I__16099 (
            .O(N__65031),
            .I(clock_c_g));
    SRMux I__16098 (
            .O(N__65028),
            .I(N__64830));
    SRMux I__16097 (
            .O(N__65027),
            .I(N__64830));
    SRMux I__16096 (
            .O(N__65026),
            .I(N__64830));
    SRMux I__16095 (
            .O(N__65025),
            .I(N__64830));
    SRMux I__16094 (
            .O(N__65024),
            .I(N__64830));
    SRMux I__16093 (
            .O(N__65023),
            .I(N__64830));
    SRMux I__16092 (
            .O(N__65022),
            .I(N__64830));
    SRMux I__16091 (
            .O(N__65021),
            .I(N__64830));
    SRMux I__16090 (
            .O(N__65020),
            .I(N__64830));
    SRMux I__16089 (
            .O(N__65019),
            .I(N__64830));
    SRMux I__16088 (
            .O(N__65018),
            .I(N__64830));
    SRMux I__16087 (
            .O(N__65017),
            .I(N__64830));
    SRMux I__16086 (
            .O(N__65016),
            .I(N__64830));
    SRMux I__16085 (
            .O(N__65015),
            .I(N__64830));
    SRMux I__16084 (
            .O(N__65014),
            .I(N__64830));
    SRMux I__16083 (
            .O(N__65013),
            .I(N__64830));
    SRMux I__16082 (
            .O(N__65012),
            .I(N__64830));
    SRMux I__16081 (
            .O(N__65011),
            .I(N__64830));
    SRMux I__16080 (
            .O(N__65010),
            .I(N__64830));
    SRMux I__16079 (
            .O(N__65009),
            .I(N__64830));
    SRMux I__16078 (
            .O(N__65008),
            .I(N__64830));
    SRMux I__16077 (
            .O(N__65007),
            .I(N__64830));
    SRMux I__16076 (
            .O(N__65006),
            .I(N__64830));
    SRMux I__16075 (
            .O(N__65005),
            .I(N__64830));
    SRMux I__16074 (
            .O(N__65004),
            .I(N__64830));
    SRMux I__16073 (
            .O(N__65003),
            .I(N__64830));
    SRMux I__16072 (
            .O(N__65002),
            .I(N__64830));
    SRMux I__16071 (
            .O(N__65001),
            .I(N__64830));
    SRMux I__16070 (
            .O(N__65000),
            .I(N__64830));
    SRMux I__16069 (
            .O(N__64999),
            .I(N__64830));
    SRMux I__16068 (
            .O(N__64998),
            .I(N__64830));
    SRMux I__16067 (
            .O(N__64997),
            .I(N__64830));
    SRMux I__16066 (
            .O(N__64996),
            .I(N__64830));
    SRMux I__16065 (
            .O(N__64995),
            .I(N__64830));
    SRMux I__16064 (
            .O(N__64994),
            .I(N__64830));
    SRMux I__16063 (
            .O(N__64993),
            .I(N__64830));
    SRMux I__16062 (
            .O(N__64992),
            .I(N__64830));
    SRMux I__16061 (
            .O(N__64991),
            .I(N__64830));
    SRMux I__16060 (
            .O(N__64990),
            .I(N__64830));
    SRMux I__16059 (
            .O(N__64989),
            .I(N__64830));
    SRMux I__16058 (
            .O(N__64988),
            .I(N__64830));
    SRMux I__16057 (
            .O(N__64987),
            .I(N__64830));
    SRMux I__16056 (
            .O(N__64986),
            .I(N__64830));
    SRMux I__16055 (
            .O(N__64985),
            .I(N__64830));
    SRMux I__16054 (
            .O(N__64984),
            .I(N__64830));
    SRMux I__16053 (
            .O(N__64983),
            .I(N__64830));
    SRMux I__16052 (
            .O(N__64982),
            .I(N__64830));
    SRMux I__16051 (
            .O(N__64981),
            .I(N__64830));
    SRMux I__16050 (
            .O(N__64980),
            .I(N__64830));
    SRMux I__16049 (
            .O(N__64979),
            .I(N__64830));
    SRMux I__16048 (
            .O(N__64978),
            .I(N__64830));
    SRMux I__16047 (
            .O(N__64977),
            .I(N__64830));
    SRMux I__16046 (
            .O(N__64976),
            .I(N__64830));
    SRMux I__16045 (
            .O(N__64975),
            .I(N__64830));
    SRMux I__16044 (
            .O(N__64974),
            .I(N__64830));
    SRMux I__16043 (
            .O(N__64973),
            .I(N__64830));
    SRMux I__16042 (
            .O(N__64972),
            .I(N__64830));
    SRMux I__16041 (
            .O(N__64971),
            .I(N__64830));
    SRMux I__16040 (
            .O(N__64970),
            .I(N__64830));
    SRMux I__16039 (
            .O(N__64969),
            .I(N__64830));
    SRMux I__16038 (
            .O(N__64968),
            .I(N__64830));
    SRMux I__16037 (
            .O(N__64967),
            .I(N__64830));
    SRMux I__16036 (
            .O(N__64966),
            .I(N__64830));
    SRMux I__16035 (
            .O(N__64965),
            .I(N__64830));
    SRMux I__16034 (
            .O(N__64964),
            .I(N__64830));
    SRMux I__16033 (
            .O(N__64963),
            .I(N__64830));
    GlobalMux I__16032 (
            .O(N__64830),
            .I(N__64827));
    gio2CtrlBuf I__16031 (
            .O(N__64827),
            .I(\I2C_top_level_inst1.c_state4_0_i_g ));
    CascadeMux I__16030 (
            .O(N__64824),
            .I(N__64821));
    InMux I__16029 (
            .O(N__64821),
            .I(N__64818));
    LocalMux I__16028 (
            .O(N__64818),
            .I(N__64815));
    Span4Mux_h I__16027 (
            .O(N__64815),
            .I(N__64812));
    Odrv4 I__16026 (
            .O(N__64812),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1666 ));
    InMux I__16025 (
            .O(N__64809),
            .I(N__64806));
    LocalMux I__16024 (
            .O(N__64806),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_1 ));
    InMux I__16023 (
            .O(N__64803),
            .I(N__64798));
    InMux I__16022 (
            .O(N__64802),
            .I(N__64795));
    CascadeMux I__16021 (
            .O(N__64801),
            .I(N__64791));
    LocalMux I__16020 (
            .O(N__64798),
            .I(N__64784));
    LocalMux I__16019 (
            .O(N__64795),
            .I(N__64781));
    InMux I__16018 (
            .O(N__64794),
            .I(N__64778));
    InMux I__16017 (
            .O(N__64791),
            .I(N__64775));
    InMux I__16016 (
            .O(N__64790),
            .I(N__64772));
    CascadeMux I__16015 (
            .O(N__64789),
            .I(N__64769));
    InMux I__16014 (
            .O(N__64788),
            .I(N__64766));
    InMux I__16013 (
            .O(N__64787),
            .I(N__64763));
    Span4Mux_v I__16012 (
            .O(N__64784),
            .I(N__64756));
    Span4Mux_v I__16011 (
            .O(N__64781),
            .I(N__64756));
    LocalMux I__16010 (
            .O(N__64778),
            .I(N__64756));
    LocalMux I__16009 (
            .O(N__64775),
            .I(N__64751));
    LocalMux I__16008 (
            .O(N__64772),
            .I(N__64751));
    InMux I__16007 (
            .O(N__64769),
            .I(N__64748));
    LocalMux I__16006 (
            .O(N__64766),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ));
    LocalMux I__16005 (
            .O(N__64763),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ));
    Odrv4 I__16004 (
            .O(N__64756),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ));
    Odrv4 I__16003 (
            .O(N__64751),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ));
    LocalMux I__16002 (
            .O(N__64748),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ));
    CascadeMux I__16001 (
            .O(N__64737),
            .I(N__64734));
    InMux I__16000 (
            .O(N__64734),
            .I(N__64731));
    LocalMux I__15999 (
            .O(N__64731),
            .I(N__64728));
    Span4Mux_h I__15998 (
            .O(N__64728),
            .I(N__64725));
    Odrv4 I__15997 (
            .O(N__64725),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_2_1 ));
    InMux I__15996 (
            .O(N__64722),
            .I(N__64716));
    InMux I__15995 (
            .O(N__64721),
            .I(N__64716));
    LocalMux I__15994 (
            .O(N__64716),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0 ));
    InMux I__15993 (
            .O(N__64713),
            .I(N__64709));
    InMux I__15992 (
            .O(N__64712),
            .I(N__64701));
    LocalMux I__15991 (
            .O(N__64709),
            .I(N__64698));
    InMux I__15990 (
            .O(N__64708),
            .I(N__64693));
    InMux I__15989 (
            .O(N__64707),
            .I(N__64688));
    InMux I__15988 (
            .O(N__64706),
            .I(N__64688));
    InMux I__15987 (
            .O(N__64705),
            .I(N__64680));
    InMux I__15986 (
            .O(N__64704),
            .I(N__64680));
    LocalMux I__15985 (
            .O(N__64701),
            .I(N__64674));
    Span4Mux_h I__15984 (
            .O(N__64698),
            .I(N__64674));
    InMux I__15983 (
            .O(N__64697),
            .I(N__64669));
    InMux I__15982 (
            .O(N__64696),
            .I(N__64669));
    LocalMux I__15981 (
            .O(N__64693),
            .I(N__64664));
    LocalMux I__15980 (
            .O(N__64688),
            .I(N__64664));
    InMux I__15979 (
            .O(N__64687),
            .I(N__64657));
    InMux I__15978 (
            .O(N__64686),
            .I(N__64657));
    InMux I__15977 (
            .O(N__64685),
            .I(N__64657));
    LocalMux I__15976 (
            .O(N__64680),
            .I(N__64654));
    InMux I__15975 (
            .O(N__64679),
            .I(N__64651));
    Span4Mux_h I__15974 (
            .O(N__64674),
            .I(N__64648));
    LocalMux I__15973 (
            .O(N__64669),
            .I(N__64641));
    Span4Mux_v I__15972 (
            .O(N__64664),
            .I(N__64641));
    LocalMux I__15971 (
            .O(N__64657),
            .I(N__64641));
    Span4Mux_h I__15970 (
            .O(N__64654),
            .I(N__64638));
    LocalMux I__15969 (
            .O(N__64651),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7 ));
    Odrv4 I__15968 (
            .O(N__64648),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7 ));
    Odrv4 I__15967 (
            .O(N__64641),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7 ));
    Odrv4 I__15966 (
            .O(N__64638),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7 ));
    InMux I__15965 (
            .O(N__64629),
            .I(N__64626));
    LocalMux I__15964 (
            .O(N__64626),
            .I(N__64623));
    Span4Mux_h I__15963 (
            .O(N__64623),
            .I(N__64620));
    Odrv4 I__15962 (
            .O(N__64620),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o3_1 ));
    CascadeMux I__15961 (
            .O(N__64617),
            .I(N__64614));
    InMux I__15960 (
            .O(N__64614),
            .I(N__64611));
    LocalMux I__15959 (
            .O(N__64611),
            .I(N__64608));
    Odrv4 I__15958 (
            .O(N__64608),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1802 ));
    InMux I__15957 (
            .O(N__64605),
            .I(N__64602));
    LocalMux I__15956 (
            .O(N__64602),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1609_0 ));
    InMux I__15955 (
            .O(N__64599),
            .I(N__64596));
    LocalMux I__15954 (
            .O(N__64596),
            .I(N__64593));
    Span4Mux_v I__15953 (
            .O(N__64593),
            .I(N__64590));
    Span4Mux_h I__15952 (
            .O(N__64590),
            .I(N__64587));
    Odrv4 I__15951 (
            .O(N__64587),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa ));
    CascadeMux I__15950 (
            .O(N__64584),
            .I(N__64578));
    InMux I__15949 (
            .O(N__64583),
            .I(N__64561));
    InMux I__15948 (
            .O(N__64582),
            .I(N__64561));
    InMux I__15947 (
            .O(N__64581),
            .I(N__64561));
    InMux I__15946 (
            .O(N__64578),
            .I(N__64561));
    InMux I__15945 (
            .O(N__64577),
            .I(N__64552));
    InMux I__15944 (
            .O(N__64576),
            .I(N__64552));
    InMux I__15943 (
            .O(N__64575),
            .I(N__64552));
    InMux I__15942 (
            .O(N__64574),
            .I(N__64552));
    InMux I__15941 (
            .O(N__64573),
            .I(N__64542));
    InMux I__15940 (
            .O(N__64572),
            .I(N__64542));
    InMux I__15939 (
            .O(N__64571),
            .I(N__64542));
    InMux I__15938 (
            .O(N__64570),
            .I(N__64542));
    LocalMux I__15937 (
            .O(N__64561),
            .I(N__64539));
    LocalMux I__15936 (
            .O(N__64552),
            .I(N__64536));
    InMux I__15935 (
            .O(N__64551),
            .I(N__64533));
    LocalMux I__15934 (
            .O(N__64542),
            .I(N__64526));
    Span4Mux_v I__15933 (
            .O(N__64539),
            .I(N__64526));
    Span4Mux_v I__15932 (
            .O(N__64536),
            .I(N__64526));
    LocalMux I__15931 (
            .O(N__64533),
            .I(N__64523));
    Span4Mux_h I__15930 (
            .O(N__64526),
            .I(N__64518));
    Span4Mux_v I__15929 (
            .O(N__64523),
            .I(N__64518));
    Odrv4 I__15928 (
            .O(N__64518),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0 ));
    CascadeMux I__15927 (
            .O(N__64515),
            .I(N__64512));
    InMux I__15926 (
            .O(N__64512),
            .I(N__64509));
    LocalMux I__15925 (
            .O(N__64509),
            .I(N__64506));
    Span4Mux_h I__15924 (
            .O(N__64506),
            .I(N__64503));
    Span4Mux_h I__15923 (
            .O(N__64503),
            .I(N__64500));
    Odrv4 I__15922 (
            .O(N__64500),
            .I(\I2C_top_level_inst1.s_addr0_o_0 ));
    InMux I__15921 (
            .O(N__64497),
            .I(N__64493));
    InMux I__15920 (
            .O(N__64496),
            .I(N__64490));
    LocalMux I__15919 (
            .O(N__64493),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_691 ));
    LocalMux I__15918 (
            .O(N__64490),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_691 ));
    InMux I__15917 (
            .O(N__64485),
            .I(N__64482));
    LocalMux I__15916 (
            .O(N__64482),
            .I(N__64479));
    Odrv12 I__15915 (
            .O(N__64479),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_0 ));
    CascadeMux I__15914 (
            .O(N__64476),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_295_cascade_ ));
    InMux I__15913 (
            .O(N__64473),
            .I(N__64469));
    InMux I__15912 (
            .O(N__64472),
            .I(N__64466));
    LocalMux I__15911 (
            .O(N__64469),
            .I(N__64462));
    LocalMux I__15910 (
            .O(N__64466),
            .I(N__64459));
    InMux I__15909 (
            .O(N__64465),
            .I(N__64454));
    Span4Mux_v I__15908 (
            .O(N__64462),
            .I(N__64449));
    Span4Mux_h I__15907 (
            .O(N__64459),
            .I(N__64449));
    InMux I__15906 (
            .O(N__64458),
            .I(N__64444));
    InMux I__15905 (
            .O(N__64457),
            .I(N__64444));
    LocalMux I__15904 (
            .O(N__64454),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3 ));
    Odrv4 I__15903 (
            .O(N__64449),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3 ));
    LocalMux I__15902 (
            .O(N__64444),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3 ));
    CascadeMux I__15901 (
            .O(N__64437),
            .I(N__64434));
    InMux I__15900 (
            .O(N__64434),
            .I(N__64429));
    InMux I__15899 (
            .O(N__64433),
            .I(N__64426));
    InMux I__15898 (
            .O(N__64432),
            .I(N__64422));
    LocalMux I__15897 (
            .O(N__64429),
            .I(N__64417));
    LocalMux I__15896 (
            .O(N__64426),
            .I(N__64414));
    InMux I__15895 (
            .O(N__64425),
            .I(N__64411));
    LocalMux I__15894 (
            .O(N__64422),
            .I(N__64408));
    InMux I__15893 (
            .O(N__64421),
            .I(N__64401));
    InMux I__15892 (
            .O(N__64420),
            .I(N__64401));
    Span4Mux_h I__15891 (
            .O(N__64417),
            .I(N__64398));
    Span4Mux_h I__15890 (
            .O(N__64414),
            .I(N__64393));
    LocalMux I__15889 (
            .O(N__64411),
            .I(N__64393));
    Span4Mux_h I__15888 (
            .O(N__64408),
            .I(N__64390));
    InMux I__15887 (
            .O(N__64407),
            .I(N__64385));
    InMux I__15886 (
            .O(N__64406),
            .I(N__64385));
    LocalMux I__15885 (
            .O(N__64401),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ));
    Odrv4 I__15884 (
            .O(N__64398),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ));
    Odrv4 I__15883 (
            .O(N__64393),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ));
    Odrv4 I__15882 (
            .O(N__64390),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ));
    LocalMux I__15881 (
            .O(N__64385),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ));
    InMux I__15880 (
            .O(N__64374),
            .I(N__64371));
    LocalMux I__15879 (
            .O(N__64371),
            .I(N__64368));
    Span4Mux_h I__15878 (
            .O(N__64368),
            .I(N__64365));
    Span4Mux_h I__15877 (
            .O(N__64365),
            .I(N__64362));
    Odrv4 I__15876 (
            .O(N__64362),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_6 ));
    InMux I__15875 (
            .O(N__64359),
            .I(N__64356));
    LocalMux I__15874 (
            .O(N__64356),
            .I(N__64352));
    InMux I__15873 (
            .O(N__64355),
            .I(N__64349));
    Odrv4 I__15872 (
            .O(N__64352),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0 ));
    LocalMux I__15871 (
            .O(N__64349),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0 ));
    InMux I__15870 (
            .O(N__64344),
            .I(N__64340));
    InMux I__15869 (
            .O(N__64343),
            .I(N__64337));
    LocalMux I__15868 (
            .O(N__64340),
            .I(N__64334));
    LocalMux I__15867 (
            .O(N__64337),
            .I(N__64331));
    Span4Mux_h I__15866 (
            .O(N__64334),
            .I(N__64328));
    Odrv4 I__15865 (
            .O(N__64331),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2));
    Odrv4 I__15864 (
            .O(N__64328),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2));
    InMux I__15863 (
            .O(N__64323),
            .I(N__64320));
    LocalMux I__15862 (
            .O(N__64320),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_277 ));
    CascadeMux I__15861 (
            .O(N__64317),
            .I(N__64313));
    InMux I__15860 (
            .O(N__64316),
            .I(N__64309));
    InMux I__15859 (
            .O(N__64313),
            .I(N__64306));
    InMux I__15858 (
            .O(N__64312),
            .I(N__64303));
    LocalMux I__15857 (
            .O(N__64309),
            .I(N__64300));
    LocalMux I__15856 (
            .O(N__64306),
            .I(N__64296));
    LocalMux I__15855 (
            .O(N__64303),
            .I(N__64293));
    Span4Mux_v I__15854 (
            .O(N__64300),
            .I(N__64290));
    InMux I__15853 (
            .O(N__64299),
            .I(N__64287));
    Span12Mux_h I__15852 (
            .O(N__64296),
            .I(N__64284));
    Span4Mux_v I__15851 (
            .O(N__64293),
            .I(N__64281));
    Sp12to4 I__15850 (
            .O(N__64290),
            .I(N__64274));
    LocalMux I__15849 (
            .O(N__64287),
            .I(N__64274));
    Span12Mux_v I__15848 (
            .O(N__64284),
            .I(N__64274));
    Odrv4 I__15847 (
            .O(N__64281),
            .I(N_552_i));
    Odrv12 I__15846 (
            .O(N__64274),
            .I(N_552_i));
    InMux I__15845 (
            .O(N__64269),
            .I(N__64262));
    InMux I__15844 (
            .O(N__64268),
            .I(N__64256));
    InMux I__15843 (
            .O(N__64267),
            .I(N__64253));
    InMux I__15842 (
            .O(N__64266),
            .I(N__64240));
    InMux I__15841 (
            .O(N__64265),
            .I(N__64237));
    LocalMux I__15840 (
            .O(N__64262),
            .I(N__64231));
    InMux I__15839 (
            .O(N__64261),
            .I(N__64225));
    InMux I__15838 (
            .O(N__64260),
            .I(N__64220));
    InMux I__15837 (
            .O(N__64259),
            .I(N__64220));
    LocalMux I__15836 (
            .O(N__64256),
            .I(N__64210));
    LocalMux I__15835 (
            .O(N__64253),
            .I(N__64198));
    InMux I__15834 (
            .O(N__64252),
            .I(N__64193));
    InMux I__15833 (
            .O(N__64251),
            .I(N__64193));
    InMux I__15832 (
            .O(N__64250),
            .I(N__64190));
    InMux I__15831 (
            .O(N__64249),
            .I(N__64175));
    InMux I__15830 (
            .O(N__64248),
            .I(N__64175));
    InMux I__15829 (
            .O(N__64247),
            .I(N__64175));
    InMux I__15828 (
            .O(N__64246),
            .I(N__64175));
    InMux I__15827 (
            .O(N__64245),
            .I(N__64175));
    InMux I__15826 (
            .O(N__64244),
            .I(N__64175));
    InMux I__15825 (
            .O(N__64243),
            .I(N__64175));
    LocalMux I__15824 (
            .O(N__64240),
            .I(N__64169));
    LocalMux I__15823 (
            .O(N__64237),
            .I(N__64166));
    InMux I__15822 (
            .O(N__64236),
            .I(N__64161));
    InMux I__15821 (
            .O(N__64235),
            .I(N__64161));
    InMux I__15820 (
            .O(N__64234),
            .I(N__64158));
    Span4Mux_h I__15819 (
            .O(N__64231),
            .I(N__64154));
    InMux I__15818 (
            .O(N__64230),
            .I(N__64149));
    InMux I__15817 (
            .O(N__64229),
            .I(N__64144));
    InMux I__15816 (
            .O(N__64228),
            .I(N__64144));
    LocalMux I__15815 (
            .O(N__64225),
            .I(N__64139));
    LocalMux I__15814 (
            .O(N__64220),
            .I(N__64139));
    InMux I__15813 (
            .O(N__64219),
            .I(N__64124));
    InMux I__15812 (
            .O(N__64218),
            .I(N__64124));
    InMux I__15811 (
            .O(N__64217),
            .I(N__64124));
    InMux I__15810 (
            .O(N__64216),
            .I(N__64124));
    InMux I__15809 (
            .O(N__64215),
            .I(N__64124));
    InMux I__15808 (
            .O(N__64214),
            .I(N__64124));
    InMux I__15807 (
            .O(N__64213),
            .I(N__64124));
    Span4Mux_h I__15806 (
            .O(N__64210),
            .I(N__64121));
    CascadeMux I__15805 (
            .O(N__64209),
            .I(N__64118));
    InMux I__15804 (
            .O(N__64208),
            .I(N__64100));
    InMux I__15803 (
            .O(N__64207),
            .I(N__64100));
    InMux I__15802 (
            .O(N__64206),
            .I(N__64100));
    InMux I__15801 (
            .O(N__64205),
            .I(N__64100));
    InMux I__15800 (
            .O(N__64204),
            .I(N__64100));
    InMux I__15799 (
            .O(N__64203),
            .I(N__64100));
    InMux I__15798 (
            .O(N__64202),
            .I(N__64100));
    InMux I__15797 (
            .O(N__64201),
            .I(N__64100));
    Span4Mux_h I__15796 (
            .O(N__64198),
            .I(N__64095));
    LocalMux I__15795 (
            .O(N__64193),
            .I(N__64095));
    LocalMux I__15794 (
            .O(N__64190),
            .I(N__64092));
    LocalMux I__15793 (
            .O(N__64175),
            .I(N__64089));
    InMux I__15792 (
            .O(N__64174),
            .I(N__64082));
    InMux I__15791 (
            .O(N__64173),
            .I(N__64082));
    InMux I__15790 (
            .O(N__64172),
            .I(N__64082));
    Span4Mux_h I__15789 (
            .O(N__64169),
            .I(N__64078));
    Span4Mux_h I__15788 (
            .O(N__64166),
            .I(N__64075));
    LocalMux I__15787 (
            .O(N__64161),
            .I(N__64061));
    LocalMux I__15786 (
            .O(N__64158),
            .I(N__64061));
    InMux I__15785 (
            .O(N__64157),
            .I(N__64058));
    Span4Mux_h I__15784 (
            .O(N__64154),
            .I(N__64055));
    InMux I__15783 (
            .O(N__64153),
            .I(N__64050));
    InMux I__15782 (
            .O(N__64152),
            .I(N__64050));
    LocalMux I__15781 (
            .O(N__64149),
            .I(N__64043));
    LocalMux I__15780 (
            .O(N__64144),
            .I(N__64043));
    Span4Mux_v I__15779 (
            .O(N__64139),
            .I(N__64043));
    LocalMux I__15778 (
            .O(N__64124),
            .I(N__64038));
    Span4Mux_v I__15777 (
            .O(N__64121),
            .I(N__64038));
    InMux I__15776 (
            .O(N__64118),
            .I(N__64033));
    InMux I__15775 (
            .O(N__64117),
            .I(N__64033));
    LocalMux I__15774 (
            .O(N__64100),
            .I(N__64028));
    Span4Mux_v I__15773 (
            .O(N__64095),
            .I(N__64028));
    Span4Mux_h I__15772 (
            .O(N__64092),
            .I(N__64021));
    Span4Mux_v I__15771 (
            .O(N__64089),
            .I(N__64021));
    LocalMux I__15770 (
            .O(N__64082),
            .I(N__64021));
    InMux I__15769 (
            .O(N__64081),
            .I(N__64018));
    Span4Mux_h I__15768 (
            .O(N__64078),
            .I(N__64013));
    Span4Mux_h I__15767 (
            .O(N__64075),
            .I(N__64013));
    InMux I__15766 (
            .O(N__64074),
            .I(N__64010));
    InMux I__15765 (
            .O(N__64073),
            .I(N__64007));
    InMux I__15764 (
            .O(N__64072),
            .I(N__64000));
    InMux I__15763 (
            .O(N__64071),
            .I(N__64000));
    InMux I__15762 (
            .O(N__64070),
            .I(N__64000));
    InMux I__15761 (
            .O(N__64069),
            .I(N__63991));
    InMux I__15760 (
            .O(N__64068),
            .I(N__63991));
    InMux I__15759 (
            .O(N__64067),
            .I(N__63991));
    InMux I__15758 (
            .O(N__64066),
            .I(N__63991));
    Span4Mux_v I__15757 (
            .O(N__64061),
            .I(N__63988));
    LocalMux I__15756 (
            .O(N__64058),
            .I(N__63977));
    Span4Mux_v I__15755 (
            .O(N__64055),
            .I(N__63977));
    LocalMux I__15754 (
            .O(N__64050),
            .I(N__63977));
    Span4Mux_h I__15753 (
            .O(N__64043),
            .I(N__63977));
    Span4Mux_v I__15752 (
            .O(N__64038),
            .I(N__63977));
    LocalMux I__15751 (
            .O(N__64033),
            .I(N__63970));
    Span4Mux_h I__15750 (
            .O(N__64028),
            .I(N__63970));
    Span4Mux_v I__15749 (
            .O(N__64021),
            .I(N__63970));
    LocalMux I__15748 (
            .O(N__64018),
            .I(N_1838_0));
    Odrv4 I__15747 (
            .O(N__64013),
            .I(N_1838_0));
    LocalMux I__15746 (
            .O(N__64010),
            .I(N_1838_0));
    LocalMux I__15745 (
            .O(N__64007),
            .I(N_1838_0));
    LocalMux I__15744 (
            .O(N__64000),
            .I(N_1838_0));
    LocalMux I__15743 (
            .O(N__63991),
            .I(N_1838_0));
    Odrv4 I__15742 (
            .O(N__63988),
            .I(N_1838_0));
    Odrv4 I__15741 (
            .O(N__63977),
            .I(N_1838_0));
    Odrv4 I__15740 (
            .O(N__63970),
            .I(N_1838_0));
    InMux I__15739 (
            .O(N__63951),
            .I(N__63948));
    LocalMux I__15738 (
            .O(N__63948),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_2 ));
    InMux I__15737 (
            .O(N__63945),
            .I(N__63941));
    InMux I__15736 (
            .O(N__63944),
            .I(N__63936));
    LocalMux I__15735 (
            .O(N__63941),
            .I(N__63933));
    InMux I__15734 (
            .O(N__63940),
            .I(N__63930));
    InMux I__15733 (
            .O(N__63939),
            .I(N__63927));
    LocalMux I__15732 (
            .O(N__63936),
            .I(N__63924));
    Span4Mux_v I__15731 (
            .O(N__63933),
            .I(N__63918));
    LocalMux I__15730 (
            .O(N__63930),
            .I(N__63918));
    LocalMux I__15729 (
            .O(N__63927),
            .I(N__63915));
    Span4Mux_v I__15728 (
            .O(N__63924),
            .I(N__63911));
    InMux I__15727 (
            .O(N__63923),
            .I(N__63906));
    Span4Mux_v I__15726 (
            .O(N__63918),
            .I(N__63902));
    Span4Mux_v I__15725 (
            .O(N__63915),
            .I(N__63899));
    InMux I__15724 (
            .O(N__63914),
            .I(N__63896));
    Span4Mux_v I__15723 (
            .O(N__63911),
            .I(N__63893));
    InMux I__15722 (
            .O(N__63910),
            .I(N__63890));
    InMux I__15721 (
            .O(N__63909),
            .I(N__63887));
    LocalMux I__15720 (
            .O(N__63906),
            .I(N__63884));
    InMux I__15719 (
            .O(N__63905),
            .I(N__63881));
    Span4Mux_h I__15718 (
            .O(N__63902),
            .I(N__63878));
    Span4Mux_h I__15717 (
            .O(N__63899),
            .I(N__63873));
    LocalMux I__15716 (
            .O(N__63896),
            .I(N__63873));
    Sp12to4 I__15715 (
            .O(N__63893),
            .I(N__63870));
    LocalMux I__15714 (
            .O(N__63890),
            .I(N__63867));
    LocalMux I__15713 (
            .O(N__63887),
            .I(N__63864));
    Span4Mux_v I__15712 (
            .O(N__63884),
            .I(N__63859));
    LocalMux I__15711 (
            .O(N__63881),
            .I(N__63859));
    Span4Mux_h I__15710 (
            .O(N__63878),
            .I(N__63854));
    Span4Mux_v I__15709 (
            .O(N__63873),
            .I(N__63854));
    Span12Mux_h I__15708 (
            .O(N__63870),
            .I(N__63851));
    Span4Mux_v I__15707 (
            .O(N__63867),
            .I(N__63844));
    Span4Mux_v I__15706 (
            .O(N__63864),
            .I(N__63844));
    Span4Mux_h I__15705 (
            .O(N__63859),
            .I(N__63844));
    Odrv4 I__15704 (
            .O(N__63854),
            .I(I2C_top_level_inst1_s_data_oreg_3));
    Odrv12 I__15703 (
            .O(N__63851),
            .I(I2C_top_level_inst1_s_data_oreg_3));
    Odrv4 I__15702 (
            .O(N__63844),
            .I(I2C_top_level_inst1_s_data_oreg_3));
    InMux I__15701 (
            .O(N__63837),
            .I(N__63834));
    LocalMux I__15700 (
            .O(N__63834),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_3 ));
    CascadeMux I__15699 (
            .O(N__63831),
            .I(N__63828));
    InMux I__15698 (
            .O(N__63828),
            .I(N__63823));
    InMux I__15697 (
            .O(N__63827),
            .I(N__63819));
    InMux I__15696 (
            .O(N__63826),
            .I(N__63816));
    LocalMux I__15695 (
            .O(N__63823),
            .I(N__63813));
    InMux I__15694 (
            .O(N__63822),
            .I(N__63810));
    LocalMux I__15693 (
            .O(N__63819),
            .I(N__63806));
    LocalMux I__15692 (
            .O(N__63816),
            .I(N__63803));
    Span4Mux_v I__15691 (
            .O(N__63813),
            .I(N__63800));
    LocalMux I__15690 (
            .O(N__63810),
            .I(N__63796));
    InMux I__15689 (
            .O(N__63809),
            .I(N__63793));
    Span4Mux_v I__15688 (
            .O(N__63806),
            .I(N__63790));
    Span4Mux_h I__15687 (
            .O(N__63803),
            .I(N__63786));
    Span4Mux_h I__15686 (
            .O(N__63800),
            .I(N__63782));
    InMux I__15685 (
            .O(N__63799),
            .I(N__63779));
    Span4Mux_h I__15684 (
            .O(N__63796),
            .I(N__63776));
    LocalMux I__15683 (
            .O(N__63793),
            .I(N__63770));
    Span4Mux_h I__15682 (
            .O(N__63790),
            .I(N__63770));
    InMux I__15681 (
            .O(N__63789),
            .I(N__63767));
    Sp12to4 I__15680 (
            .O(N__63786),
            .I(N__63764));
    InMux I__15679 (
            .O(N__63785),
            .I(N__63761));
    Span4Mux_h I__15678 (
            .O(N__63782),
            .I(N__63756));
    LocalMux I__15677 (
            .O(N__63779),
            .I(N__63756));
    Span4Mux_h I__15676 (
            .O(N__63776),
            .I(N__63753));
    InMux I__15675 (
            .O(N__63775),
            .I(N__63750));
    Span4Mux_v I__15674 (
            .O(N__63770),
            .I(N__63747));
    LocalMux I__15673 (
            .O(N__63767),
            .I(N__63742));
    Span12Mux_v I__15672 (
            .O(N__63764),
            .I(N__63742));
    LocalMux I__15671 (
            .O(N__63761),
            .I(N__63739));
    Span4Mux_v I__15670 (
            .O(N__63756),
            .I(N__63736));
    Span4Mux_v I__15669 (
            .O(N__63753),
            .I(N__63733));
    LocalMux I__15668 (
            .O(N__63750),
            .I(N__63730));
    Span4Mux_h I__15667 (
            .O(N__63747),
            .I(N__63727));
    Span12Mux_h I__15666 (
            .O(N__63742),
            .I(N__63724));
    Span4Mux_v I__15665 (
            .O(N__63739),
            .I(N__63719));
    Span4Mux_v I__15664 (
            .O(N__63736),
            .I(N__63719));
    Odrv4 I__15663 (
            .O(N__63733),
            .I(I2C_top_level_inst1_s_data_oreg_4));
    Odrv4 I__15662 (
            .O(N__63730),
            .I(I2C_top_level_inst1_s_data_oreg_4));
    Odrv4 I__15661 (
            .O(N__63727),
            .I(I2C_top_level_inst1_s_data_oreg_4));
    Odrv12 I__15660 (
            .O(N__63724),
            .I(I2C_top_level_inst1_s_data_oreg_4));
    Odrv4 I__15659 (
            .O(N__63719),
            .I(I2C_top_level_inst1_s_data_oreg_4));
    InMux I__15658 (
            .O(N__63708),
            .I(N__63705));
    LocalMux I__15657 (
            .O(N__63705),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_4 ));
    InMux I__15656 (
            .O(N__63702),
            .I(N__63698));
    InMux I__15655 (
            .O(N__63701),
            .I(N__63694));
    LocalMux I__15654 (
            .O(N__63698),
            .I(N__63691));
    CascadeMux I__15653 (
            .O(N__63697),
            .I(N__63688));
    LocalMux I__15652 (
            .O(N__63694),
            .I(N__63684));
    Span4Mux_v I__15651 (
            .O(N__63691),
            .I(N__63681));
    InMux I__15650 (
            .O(N__63688),
            .I(N__63678));
    InMux I__15649 (
            .O(N__63687),
            .I(N__63674));
    Span4Mux_h I__15648 (
            .O(N__63684),
            .I(N__63671));
    Span4Mux_h I__15647 (
            .O(N__63681),
            .I(N__63665));
    LocalMux I__15646 (
            .O(N__63678),
            .I(N__63665));
    InMux I__15645 (
            .O(N__63677),
            .I(N__63662));
    LocalMux I__15644 (
            .O(N__63674),
            .I(N__63658));
    Span4Mux_v I__15643 (
            .O(N__63671),
            .I(N__63654));
    CascadeMux I__15642 (
            .O(N__63670),
            .I(N__63651));
    Span4Mux_v I__15641 (
            .O(N__63665),
            .I(N__63646));
    LocalMux I__15640 (
            .O(N__63662),
            .I(N__63646));
    InMux I__15639 (
            .O(N__63661),
            .I(N__63642));
    Span4Mux_v I__15638 (
            .O(N__63658),
            .I(N__63639));
    InMux I__15637 (
            .O(N__63657),
            .I(N__63636));
    Sp12to4 I__15636 (
            .O(N__63654),
            .I(N__63633));
    InMux I__15635 (
            .O(N__63651),
            .I(N__63630));
    Span4Mux_h I__15634 (
            .O(N__63646),
            .I(N__63627));
    InMux I__15633 (
            .O(N__63645),
            .I(N__63624));
    LocalMux I__15632 (
            .O(N__63642),
            .I(N__63621));
    Sp12to4 I__15631 (
            .O(N__63639),
            .I(N__63612));
    LocalMux I__15630 (
            .O(N__63636),
            .I(N__63612));
    Span12Mux_v I__15629 (
            .O(N__63633),
            .I(N__63612));
    LocalMux I__15628 (
            .O(N__63630),
            .I(N__63612));
    Span4Mux_h I__15627 (
            .O(N__63627),
            .I(N__63609));
    LocalMux I__15626 (
            .O(N__63624),
            .I(N__63606));
    Span4Mux_h I__15625 (
            .O(N__63621),
            .I(N__63603));
    Span12Mux_h I__15624 (
            .O(N__63612),
            .I(N__63600));
    Odrv4 I__15623 (
            .O(N__63609),
            .I(I2C_top_level_inst1_s_data_oreg_5));
    Odrv12 I__15622 (
            .O(N__63606),
            .I(I2C_top_level_inst1_s_data_oreg_5));
    Odrv4 I__15621 (
            .O(N__63603),
            .I(I2C_top_level_inst1_s_data_oreg_5));
    Odrv12 I__15620 (
            .O(N__63600),
            .I(I2C_top_level_inst1_s_data_oreg_5));
    InMux I__15619 (
            .O(N__63591),
            .I(N__63588));
    LocalMux I__15618 (
            .O(N__63588),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_5 ));
    InMux I__15617 (
            .O(N__63585),
            .I(N__63577));
    InMux I__15616 (
            .O(N__63584),
            .I(N__63574));
    InMux I__15615 (
            .O(N__63583),
            .I(N__63569));
    InMux I__15614 (
            .O(N__63582),
            .I(N__63569));
    InMux I__15613 (
            .O(N__63581),
            .I(N__63565));
    InMux I__15612 (
            .O(N__63580),
            .I(N__63562));
    LocalMux I__15611 (
            .O(N__63577),
            .I(N__63559));
    LocalMux I__15610 (
            .O(N__63574),
            .I(N__63556));
    LocalMux I__15609 (
            .O(N__63569),
            .I(N__63553));
    InMux I__15608 (
            .O(N__63568),
            .I(N__63550));
    LocalMux I__15607 (
            .O(N__63565),
            .I(N__63547));
    LocalMux I__15606 (
            .O(N__63562),
            .I(N__63544));
    Span4Mux_v I__15605 (
            .O(N__63559),
            .I(N__63540));
    Span4Mux_v I__15604 (
            .O(N__63556),
            .I(N__63537));
    Span4Mux_h I__15603 (
            .O(N__63553),
            .I(N__63532));
    LocalMux I__15602 (
            .O(N__63550),
            .I(N__63532));
    Span4Mux_h I__15601 (
            .O(N__63547),
            .I(N__63527));
    Span4Mux_v I__15600 (
            .O(N__63544),
            .I(N__63527));
    InMux I__15599 (
            .O(N__63543),
            .I(N__63523));
    Sp12to4 I__15598 (
            .O(N__63540),
            .I(N__63520));
    Span4Mux_h I__15597 (
            .O(N__63537),
            .I(N__63517));
    Span4Mux_h I__15596 (
            .O(N__63532),
            .I(N__63514));
    Span4Mux_h I__15595 (
            .O(N__63527),
            .I(N__63511));
    InMux I__15594 (
            .O(N__63526),
            .I(N__63508));
    LocalMux I__15593 (
            .O(N__63523),
            .I(N__63503));
    Span12Mux_h I__15592 (
            .O(N__63520),
            .I(N__63503));
    Span4Mux_v I__15591 (
            .O(N__63517),
            .I(N__63498));
    Span4Mux_v I__15590 (
            .O(N__63514),
            .I(N__63498));
    Odrv4 I__15589 (
            .O(N__63511),
            .I(I2C_top_level_inst1_s_data_oreg_6));
    LocalMux I__15588 (
            .O(N__63508),
            .I(I2C_top_level_inst1_s_data_oreg_6));
    Odrv12 I__15587 (
            .O(N__63503),
            .I(I2C_top_level_inst1_s_data_oreg_6));
    Odrv4 I__15586 (
            .O(N__63498),
            .I(I2C_top_level_inst1_s_data_oreg_6));
    InMux I__15585 (
            .O(N__63489),
            .I(N__63486));
    LocalMux I__15584 (
            .O(N__63486),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_6 ));
    InMux I__15583 (
            .O(N__63483),
            .I(N__63478));
    InMux I__15582 (
            .O(N__63482),
            .I(N__63473));
    InMux I__15581 (
            .O(N__63481),
            .I(N__63468));
    LocalMux I__15580 (
            .O(N__63478),
            .I(N__63464));
    InMux I__15579 (
            .O(N__63477),
            .I(N__63461));
    InMux I__15578 (
            .O(N__63476),
            .I(N__63458));
    LocalMux I__15577 (
            .O(N__63473),
            .I(N__63455));
    CascadeMux I__15576 (
            .O(N__63472),
            .I(N__63452));
    InMux I__15575 (
            .O(N__63471),
            .I(N__63449));
    LocalMux I__15574 (
            .O(N__63468),
            .I(N__63445));
    InMux I__15573 (
            .O(N__63467),
            .I(N__63442));
    Span4Mux_v I__15572 (
            .O(N__63464),
            .I(N__63439));
    LocalMux I__15571 (
            .O(N__63461),
            .I(N__63436));
    LocalMux I__15570 (
            .O(N__63458),
            .I(N__63433));
    Span4Mux_v I__15569 (
            .O(N__63455),
            .I(N__63430));
    InMux I__15568 (
            .O(N__63452),
            .I(N__63427));
    LocalMux I__15567 (
            .O(N__63449),
            .I(N__63424));
    InMux I__15566 (
            .O(N__63448),
            .I(N__63421));
    Span4Mux_v I__15565 (
            .O(N__63445),
            .I(N__63418));
    LocalMux I__15564 (
            .O(N__63442),
            .I(N__63407));
    Sp12to4 I__15563 (
            .O(N__63439),
            .I(N__63407));
    Span12Mux_v I__15562 (
            .O(N__63436),
            .I(N__63407));
    Sp12to4 I__15561 (
            .O(N__63433),
            .I(N__63407));
    Sp12to4 I__15560 (
            .O(N__63430),
            .I(N__63407));
    LocalMux I__15559 (
            .O(N__63427),
            .I(N__63400));
    Span12Mux_v I__15558 (
            .O(N__63424),
            .I(N__63400));
    LocalMux I__15557 (
            .O(N__63421),
            .I(N__63400));
    Span4Mux_h I__15556 (
            .O(N__63418),
            .I(N__63397));
    Span12Mux_h I__15555 (
            .O(N__63407),
            .I(N__63394));
    Span12Mux_h I__15554 (
            .O(N__63400),
            .I(N__63391));
    Odrv4 I__15553 (
            .O(N__63397),
            .I(I2C_top_level_inst1_s_data_oreg_7));
    Odrv12 I__15552 (
            .O(N__63394),
            .I(I2C_top_level_inst1_s_data_oreg_7));
    Odrv12 I__15551 (
            .O(N__63391),
            .I(I2C_top_level_inst1_s_data_oreg_7));
    InMux I__15550 (
            .O(N__63384),
            .I(N__63359));
    InMux I__15549 (
            .O(N__63383),
            .I(N__63359));
    InMux I__15548 (
            .O(N__63382),
            .I(N__63359));
    InMux I__15547 (
            .O(N__63381),
            .I(N__63359));
    InMux I__15546 (
            .O(N__63380),
            .I(N__63359));
    InMux I__15545 (
            .O(N__63379),
            .I(N__63359));
    InMux I__15544 (
            .O(N__63378),
            .I(N__63359));
    InMux I__15543 (
            .O(N__63377),
            .I(N__63359));
    CascadeMux I__15542 (
            .O(N__63376),
            .I(N__63356));
    LocalMux I__15541 (
            .O(N__63359),
            .I(N__63338));
    InMux I__15540 (
            .O(N__63356),
            .I(N__63327));
    InMux I__15539 (
            .O(N__63355),
            .I(N__63327));
    InMux I__15538 (
            .O(N__63354),
            .I(N__63327));
    InMux I__15537 (
            .O(N__63353),
            .I(N__63327));
    InMux I__15536 (
            .O(N__63352),
            .I(N__63327));
    InMux I__15535 (
            .O(N__63351),
            .I(N__63310));
    InMux I__15534 (
            .O(N__63350),
            .I(N__63310));
    InMux I__15533 (
            .O(N__63349),
            .I(N__63310));
    InMux I__15532 (
            .O(N__63348),
            .I(N__63310));
    InMux I__15531 (
            .O(N__63347),
            .I(N__63310));
    InMux I__15530 (
            .O(N__63346),
            .I(N__63310));
    InMux I__15529 (
            .O(N__63345),
            .I(N__63310));
    InMux I__15528 (
            .O(N__63344),
            .I(N__63310));
    InMux I__15527 (
            .O(N__63343),
            .I(N__63303));
    InMux I__15526 (
            .O(N__63342),
            .I(N__63303));
    InMux I__15525 (
            .O(N__63341),
            .I(N__63303));
    Span4Mux_v I__15524 (
            .O(N__63338),
            .I(N__63285));
    LocalMux I__15523 (
            .O(N__63327),
            .I(N__63285));
    LocalMux I__15522 (
            .O(N__63310),
            .I(N__63285));
    LocalMux I__15521 (
            .O(N__63303),
            .I(N__63282));
    CascadeMux I__15520 (
            .O(N__63302),
            .I(N__63278));
    CascadeMux I__15519 (
            .O(N__63301),
            .I(N__63275));
    InMux I__15518 (
            .O(N__63300),
            .I(N__63270));
    InMux I__15517 (
            .O(N__63299),
            .I(N__63255));
    InMux I__15516 (
            .O(N__63298),
            .I(N__63255));
    InMux I__15515 (
            .O(N__63297),
            .I(N__63255));
    InMux I__15514 (
            .O(N__63296),
            .I(N__63255));
    InMux I__15513 (
            .O(N__63295),
            .I(N__63255));
    InMux I__15512 (
            .O(N__63294),
            .I(N__63255));
    InMux I__15511 (
            .O(N__63293),
            .I(N__63255));
    InMux I__15510 (
            .O(N__63292),
            .I(N__63252));
    Span4Mux_v I__15509 (
            .O(N__63285),
            .I(N__63247));
    Span4Mux_v I__15508 (
            .O(N__63282),
            .I(N__63247));
    InMux I__15507 (
            .O(N__63281),
            .I(N__63243));
    InMux I__15506 (
            .O(N__63278),
            .I(N__63238));
    InMux I__15505 (
            .O(N__63275),
            .I(N__63238));
    CascadeMux I__15504 (
            .O(N__63274),
            .I(N__63235));
    CascadeMux I__15503 (
            .O(N__63273),
            .I(N__63232));
    LocalMux I__15502 (
            .O(N__63270),
            .I(N__63225));
    LocalMux I__15501 (
            .O(N__63255),
            .I(N__63225));
    LocalMux I__15500 (
            .O(N__63252),
            .I(N__63222));
    Span4Mux_h I__15499 (
            .O(N__63247),
            .I(N__63219));
    InMux I__15498 (
            .O(N__63246),
            .I(N__63216));
    LocalMux I__15497 (
            .O(N__63243),
            .I(N__63211));
    LocalMux I__15496 (
            .O(N__63238),
            .I(N__63211));
    InMux I__15495 (
            .O(N__63235),
            .I(N__63202));
    InMux I__15494 (
            .O(N__63232),
            .I(N__63202));
    InMux I__15493 (
            .O(N__63231),
            .I(N__63202));
    InMux I__15492 (
            .O(N__63230),
            .I(N__63202));
    Span4Mux_h I__15491 (
            .O(N__63225),
            .I(N__63199));
    Span4Mux_v I__15490 (
            .O(N__63222),
            .I(N__63194));
    Sp12to4 I__15489 (
            .O(N__63219),
            .I(N__63191));
    LocalMux I__15488 (
            .O(N__63216),
            .I(N__63188));
    Span4Mux_h I__15487 (
            .O(N__63211),
            .I(N__63183));
    LocalMux I__15486 (
            .O(N__63202),
            .I(N__63183));
    Span4Mux_v I__15485 (
            .O(N__63199),
            .I(N__63180));
    InMux I__15484 (
            .O(N__63198),
            .I(N__63175));
    InMux I__15483 (
            .O(N__63197),
            .I(N__63175));
    Sp12to4 I__15482 (
            .O(N__63194),
            .I(N__63170));
    Span12Mux_v I__15481 (
            .O(N__63191),
            .I(N__63170));
    Span4Mux_v I__15480 (
            .O(N__63188),
            .I(N__63163));
    Span4Mux_v I__15479 (
            .O(N__63183),
            .I(N__63163));
    Span4Mux_h I__15478 (
            .O(N__63180),
            .I(N__63163));
    LocalMux I__15477 (
            .O(N__63175),
            .I(\I2C_top_level_inst1.s_enable_desp_tx ));
    Odrv12 I__15476 (
            .O(N__63170),
            .I(\I2C_top_level_inst1.s_enable_desp_tx ));
    Odrv4 I__15475 (
            .O(N__63163),
            .I(\I2C_top_level_inst1.s_enable_desp_tx ));
    InMux I__15474 (
            .O(N__63156),
            .I(N__63153));
    LocalMux I__15473 (
            .O(N__63153),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_7 ));
    InMux I__15472 (
            .O(N__63150),
            .I(N__63146));
    InMux I__15471 (
            .O(N__63149),
            .I(N__63141));
    LocalMux I__15470 (
            .O(N__63146),
            .I(N__63138));
    InMux I__15469 (
            .O(N__63145),
            .I(N__63135));
    InMux I__15468 (
            .O(N__63144),
            .I(N__63131));
    LocalMux I__15467 (
            .O(N__63141),
            .I(N__63128));
    Span4Mux_v I__15466 (
            .O(N__63138),
            .I(N__63123));
    LocalMux I__15465 (
            .O(N__63135),
            .I(N__63123));
    CascadeMux I__15464 (
            .O(N__63134),
            .I(N__63120));
    LocalMux I__15463 (
            .O(N__63131),
            .I(N__63115));
    Span4Mux_v I__15462 (
            .O(N__63128),
            .I(N__63110));
    Span4Mux_v I__15461 (
            .O(N__63123),
            .I(N__63110));
    InMux I__15460 (
            .O(N__63120),
            .I(N__63107));
    InMux I__15459 (
            .O(N__63119),
            .I(N__63104));
    InMux I__15458 (
            .O(N__63118),
            .I(N__63099));
    Span4Mux_v I__15457 (
            .O(N__63115),
            .I(N__63094));
    Span4Mux_h I__15456 (
            .O(N__63110),
            .I(N__63094));
    LocalMux I__15455 (
            .O(N__63107),
            .I(N__63091));
    LocalMux I__15454 (
            .O(N__63104),
            .I(N__63088));
    InMux I__15453 (
            .O(N__63103),
            .I(N__63083));
    InMux I__15452 (
            .O(N__63102),
            .I(N__63083));
    LocalMux I__15451 (
            .O(N__63099),
            .I(N__63080));
    Span4Mux_h I__15450 (
            .O(N__63094),
            .I(N__63077));
    Span4Mux_h I__15449 (
            .O(N__63091),
            .I(N__63074));
    Span4Mux_v I__15448 (
            .O(N__63088),
            .I(N__63071));
    LocalMux I__15447 (
            .O(N__63083),
            .I(N__63068));
    Span12Mux_v I__15446 (
            .O(N__63080),
            .I(N__63065));
    Span4Mux_v I__15445 (
            .O(N__63077),
            .I(N__63062));
    Span4Mux_h I__15444 (
            .O(N__63074),
            .I(N__63059));
    Span4Mux_h I__15443 (
            .O(N__63071),
            .I(N__63054));
    Span4Mux_v I__15442 (
            .O(N__63068),
            .I(N__63054));
    Odrv12 I__15441 (
            .O(N__63065),
            .I(I2C_top_level_inst1_s_data_oreg_8));
    Odrv4 I__15440 (
            .O(N__63062),
            .I(I2C_top_level_inst1_s_data_oreg_8));
    Odrv4 I__15439 (
            .O(N__63059),
            .I(I2C_top_level_inst1_s_data_oreg_8));
    Odrv4 I__15438 (
            .O(N__63054),
            .I(I2C_top_level_inst1_s_data_oreg_8));
    InMux I__15437 (
            .O(N__63045),
            .I(N__63042));
    LocalMux I__15436 (
            .O(N__63042),
            .I(N__63039));
    Span4Mux_h I__15435 (
            .O(N__63039),
            .I(N__63036));
    Span4Mux_h I__15434 (
            .O(N__63036),
            .I(N__63033));
    Odrv4 I__15433 (
            .O(N__63033),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_8 ));
    CEMux I__15432 (
            .O(N__63030),
            .I(N__63026));
    CEMux I__15431 (
            .O(N__63029),
            .I(N__63022));
    LocalMux I__15430 (
            .O(N__63026),
            .I(N__63019));
    CEMux I__15429 (
            .O(N__63025),
            .I(N__63016));
    LocalMux I__15428 (
            .O(N__63022),
            .I(N__63012));
    Span4Mux_h I__15427 (
            .O(N__63019),
            .I(N__63007));
    LocalMux I__15426 (
            .O(N__63016),
            .I(N__63007));
    CEMux I__15425 (
            .O(N__63015),
            .I(N__63004));
    Span4Mux_v I__15424 (
            .O(N__63012),
            .I(N__62999));
    Span4Mux_v I__15423 (
            .O(N__63007),
            .I(N__62994));
    LocalMux I__15422 (
            .O(N__63004),
            .I(N__62994));
    CEMux I__15421 (
            .O(N__63003),
            .I(N__62991));
    CEMux I__15420 (
            .O(N__63002),
            .I(N__62988));
    Span4Mux_h I__15419 (
            .O(N__62999),
            .I(N__62985));
    Span4Mux_v I__15418 (
            .O(N__62994),
            .I(N__62980));
    LocalMux I__15417 (
            .O(N__62991),
            .I(N__62980));
    LocalMux I__15416 (
            .O(N__62988),
            .I(N__62977));
    Span4Mux_v I__15415 (
            .O(N__62985),
            .I(N__62974));
    Span4Mux_h I__15414 (
            .O(N__62980),
            .I(N__62971));
    Span4Mux_v I__15413 (
            .O(N__62977),
            .I(N__62968));
    Odrv4 I__15412 (
            .O(N__62974),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0 ));
    Odrv4 I__15411 (
            .O(N__62971),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0 ));
    Odrv4 I__15410 (
            .O(N__62968),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0 ));
    SRMux I__15409 (
            .O(N__62961),
            .I(N__62487));
    SRMux I__15408 (
            .O(N__62960),
            .I(N__62487));
    SRMux I__15407 (
            .O(N__62959),
            .I(N__62487));
    SRMux I__15406 (
            .O(N__62958),
            .I(N__62487));
    SRMux I__15405 (
            .O(N__62957),
            .I(N__62487));
    SRMux I__15404 (
            .O(N__62956),
            .I(N__62487));
    SRMux I__15403 (
            .O(N__62955),
            .I(N__62487));
    SRMux I__15402 (
            .O(N__62954),
            .I(N__62487));
    SRMux I__15401 (
            .O(N__62953),
            .I(N__62487));
    SRMux I__15400 (
            .O(N__62952),
            .I(N__62487));
    SRMux I__15399 (
            .O(N__62951),
            .I(N__62487));
    SRMux I__15398 (
            .O(N__62950),
            .I(N__62487));
    SRMux I__15397 (
            .O(N__62949),
            .I(N__62487));
    SRMux I__15396 (
            .O(N__62948),
            .I(N__62487));
    SRMux I__15395 (
            .O(N__62947),
            .I(N__62487));
    SRMux I__15394 (
            .O(N__62946),
            .I(N__62487));
    SRMux I__15393 (
            .O(N__62945),
            .I(N__62487));
    SRMux I__15392 (
            .O(N__62944),
            .I(N__62487));
    SRMux I__15391 (
            .O(N__62943),
            .I(N__62487));
    SRMux I__15390 (
            .O(N__62942),
            .I(N__62487));
    SRMux I__15389 (
            .O(N__62941),
            .I(N__62487));
    SRMux I__15388 (
            .O(N__62940),
            .I(N__62487));
    SRMux I__15387 (
            .O(N__62939),
            .I(N__62487));
    SRMux I__15386 (
            .O(N__62938),
            .I(N__62487));
    SRMux I__15385 (
            .O(N__62937),
            .I(N__62487));
    SRMux I__15384 (
            .O(N__62936),
            .I(N__62487));
    SRMux I__15383 (
            .O(N__62935),
            .I(N__62487));
    SRMux I__15382 (
            .O(N__62934),
            .I(N__62487));
    SRMux I__15381 (
            .O(N__62933),
            .I(N__62487));
    SRMux I__15380 (
            .O(N__62932),
            .I(N__62487));
    SRMux I__15379 (
            .O(N__62931),
            .I(N__62487));
    SRMux I__15378 (
            .O(N__62930),
            .I(N__62487));
    SRMux I__15377 (
            .O(N__62929),
            .I(N__62487));
    SRMux I__15376 (
            .O(N__62928),
            .I(N__62487));
    SRMux I__15375 (
            .O(N__62927),
            .I(N__62487));
    SRMux I__15374 (
            .O(N__62926),
            .I(N__62487));
    SRMux I__15373 (
            .O(N__62925),
            .I(N__62487));
    SRMux I__15372 (
            .O(N__62924),
            .I(N__62487));
    SRMux I__15371 (
            .O(N__62923),
            .I(N__62487));
    SRMux I__15370 (
            .O(N__62922),
            .I(N__62487));
    SRMux I__15369 (
            .O(N__62921),
            .I(N__62487));
    SRMux I__15368 (
            .O(N__62920),
            .I(N__62487));
    SRMux I__15367 (
            .O(N__62919),
            .I(N__62487));
    SRMux I__15366 (
            .O(N__62918),
            .I(N__62487));
    SRMux I__15365 (
            .O(N__62917),
            .I(N__62487));
    SRMux I__15364 (
            .O(N__62916),
            .I(N__62487));
    SRMux I__15363 (
            .O(N__62915),
            .I(N__62487));
    SRMux I__15362 (
            .O(N__62914),
            .I(N__62487));
    SRMux I__15361 (
            .O(N__62913),
            .I(N__62487));
    SRMux I__15360 (
            .O(N__62912),
            .I(N__62487));
    SRMux I__15359 (
            .O(N__62911),
            .I(N__62487));
    SRMux I__15358 (
            .O(N__62910),
            .I(N__62487));
    SRMux I__15357 (
            .O(N__62909),
            .I(N__62487));
    SRMux I__15356 (
            .O(N__62908),
            .I(N__62487));
    SRMux I__15355 (
            .O(N__62907),
            .I(N__62487));
    SRMux I__15354 (
            .O(N__62906),
            .I(N__62487));
    SRMux I__15353 (
            .O(N__62905),
            .I(N__62487));
    SRMux I__15352 (
            .O(N__62904),
            .I(N__62487));
    SRMux I__15351 (
            .O(N__62903),
            .I(N__62487));
    SRMux I__15350 (
            .O(N__62902),
            .I(N__62487));
    SRMux I__15349 (
            .O(N__62901),
            .I(N__62487));
    SRMux I__15348 (
            .O(N__62900),
            .I(N__62487));
    SRMux I__15347 (
            .O(N__62899),
            .I(N__62487));
    SRMux I__15346 (
            .O(N__62898),
            .I(N__62487));
    SRMux I__15345 (
            .O(N__62897),
            .I(N__62487));
    SRMux I__15344 (
            .O(N__62896),
            .I(N__62487));
    SRMux I__15343 (
            .O(N__62895),
            .I(N__62487));
    SRMux I__15342 (
            .O(N__62894),
            .I(N__62487));
    SRMux I__15341 (
            .O(N__62893),
            .I(N__62487));
    SRMux I__15340 (
            .O(N__62892),
            .I(N__62487));
    SRMux I__15339 (
            .O(N__62891),
            .I(N__62487));
    SRMux I__15338 (
            .O(N__62890),
            .I(N__62487));
    SRMux I__15337 (
            .O(N__62889),
            .I(N__62487));
    SRMux I__15336 (
            .O(N__62888),
            .I(N__62487));
    SRMux I__15335 (
            .O(N__62887),
            .I(N__62487));
    SRMux I__15334 (
            .O(N__62886),
            .I(N__62487));
    SRMux I__15333 (
            .O(N__62885),
            .I(N__62487));
    SRMux I__15332 (
            .O(N__62884),
            .I(N__62487));
    SRMux I__15331 (
            .O(N__62883),
            .I(N__62487));
    SRMux I__15330 (
            .O(N__62882),
            .I(N__62487));
    SRMux I__15329 (
            .O(N__62881),
            .I(N__62487));
    SRMux I__15328 (
            .O(N__62880),
            .I(N__62487));
    SRMux I__15327 (
            .O(N__62879),
            .I(N__62487));
    SRMux I__15326 (
            .O(N__62878),
            .I(N__62487));
    SRMux I__15325 (
            .O(N__62877),
            .I(N__62487));
    SRMux I__15324 (
            .O(N__62876),
            .I(N__62487));
    SRMux I__15323 (
            .O(N__62875),
            .I(N__62487));
    SRMux I__15322 (
            .O(N__62874),
            .I(N__62487));
    SRMux I__15321 (
            .O(N__62873),
            .I(N__62487));
    SRMux I__15320 (
            .O(N__62872),
            .I(N__62487));
    SRMux I__15319 (
            .O(N__62871),
            .I(N__62487));
    SRMux I__15318 (
            .O(N__62870),
            .I(N__62487));
    SRMux I__15317 (
            .O(N__62869),
            .I(N__62487));
    SRMux I__15316 (
            .O(N__62868),
            .I(N__62487));
    SRMux I__15315 (
            .O(N__62867),
            .I(N__62487));
    SRMux I__15314 (
            .O(N__62866),
            .I(N__62487));
    SRMux I__15313 (
            .O(N__62865),
            .I(N__62487));
    SRMux I__15312 (
            .O(N__62864),
            .I(N__62487));
    SRMux I__15311 (
            .O(N__62863),
            .I(N__62487));
    SRMux I__15310 (
            .O(N__62862),
            .I(N__62487));
    SRMux I__15309 (
            .O(N__62861),
            .I(N__62487));
    SRMux I__15308 (
            .O(N__62860),
            .I(N__62487));
    SRMux I__15307 (
            .O(N__62859),
            .I(N__62487));
    SRMux I__15306 (
            .O(N__62858),
            .I(N__62487));
    SRMux I__15305 (
            .O(N__62857),
            .I(N__62487));
    SRMux I__15304 (
            .O(N__62856),
            .I(N__62487));
    SRMux I__15303 (
            .O(N__62855),
            .I(N__62487));
    SRMux I__15302 (
            .O(N__62854),
            .I(N__62487));
    SRMux I__15301 (
            .O(N__62853),
            .I(N__62487));
    SRMux I__15300 (
            .O(N__62852),
            .I(N__62487));
    SRMux I__15299 (
            .O(N__62851),
            .I(N__62487));
    SRMux I__15298 (
            .O(N__62850),
            .I(N__62487));
    SRMux I__15297 (
            .O(N__62849),
            .I(N__62487));
    SRMux I__15296 (
            .O(N__62848),
            .I(N__62487));
    SRMux I__15295 (
            .O(N__62847),
            .I(N__62487));
    SRMux I__15294 (
            .O(N__62846),
            .I(N__62487));
    SRMux I__15293 (
            .O(N__62845),
            .I(N__62487));
    SRMux I__15292 (
            .O(N__62844),
            .I(N__62487));
    SRMux I__15291 (
            .O(N__62843),
            .I(N__62487));
    SRMux I__15290 (
            .O(N__62842),
            .I(N__62487));
    SRMux I__15289 (
            .O(N__62841),
            .I(N__62487));
    SRMux I__15288 (
            .O(N__62840),
            .I(N__62487));
    SRMux I__15287 (
            .O(N__62839),
            .I(N__62487));
    SRMux I__15286 (
            .O(N__62838),
            .I(N__62487));
    SRMux I__15285 (
            .O(N__62837),
            .I(N__62487));
    SRMux I__15284 (
            .O(N__62836),
            .I(N__62487));
    SRMux I__15283 (
            .O(N__62835),
            .I(N__62487));
    SRMux I__15282 (
            .O(N__62834),
            .I(N__62487));
    SRMux I__15281 (
            .O(N__62833),
            .I(N__62487));
    SRMux I__15280 (
            .O(N__62832),
            .I(N__62487));
    SRMux I__15279 (
            .O(N__62831),
            .I(N__62487));
    SRMux I__15278 (
            .O(N__62830),
            .I(N__62487));
    SRMux I__15277 (
            .O(N__62829),
            .I(N__62487));
    SRMux I__15276 (
            .O(N__62828),
            .I(N__62487));
    SRMux I__15275 (
            .O(N__62827),
            .I(N__62487));
    SRMux I__15274 (
            .O(N__62826),
            .I(N__62487));
    SRMux I__15273 (
            .O(N__62825),
            .I(N__62487));
    SRMux I__15272 (
            .O(N__62824),
            .I(N__62487));
    SRMux I__15271 (
            .O(N__62823),
            .I(N__62487));
    SRMux I__15270 (
            .O(N__62822),
            .I(N__62487));
    SRMux I__15269 (
            .O(N__62821),
            .I(N__62487));
    SRMux I__15268 (
            .O(N__62820),
            .I(N__62487));
    SRMux I__15267 (
            .O(N__62819),
            .I(N__62487));
    SRMux I__15266 (
            .O(N__62818),
            .I(N__62487));
    SRMux I__15265 (
            .O(N__62817),
            .I(N__62487));
    SRMux I__15264 (
            .O(N__62816),
            .I(N__62487));
    SRMux I__15263 (
            .O(N__62815),
            .I(N__62487));
    SRMux I__15262 (
            .O(N__62814),
            .I(N__62487));
    SRMux I__15261 (
            .O(N__62813),
            .I(N__62487));
    SRMux I__15260 (
            .O(N__62812),
            .I(N__62487));
    SRMux I__15259 (
            .O(N__62811),
            .I(N__62487));
    SRMux I__15258 (
            .O(N__62810),
            .I(N__62487));
    SRMux I__15257 (
            .O(N__62809),
            .I(N__62487));
    SRMux I__15256 (
            .O(N__62808),
            .I(N__62487));
    SRMux I__15255 (
            .O(N__62807),
            .I(N__62487));
    SRMux I__15254 (
            .O(N__62806),
            .I(N__62487));
    SRMux I__15253 (
            .O(N__62805),
            .I(N__62487));
    SRMux I__15252 (
            .O(N__62804),
            .I(N__62487));
    GlobalMux I__15251 (
            .O(N__62487),
            .I(N__62484));
    gio2CtrlBuf I__15250 (
            .O(N__62484),
            .I(rst_n_c_i_g));
    InMux I__15249 (
            .O(N__62481),
            .I(N__62476));
    InMux I__15248 (
            .O(N__62480),
            .I(N__62473));
    InMux I__15247 (
            .O(N__62479),
            .I(N__62469));
    LocalMux I__15246 (
            .O(N__62476),
            .I(N__62466));
    LocalMux I__15245 (
            .O(N__62473),
            .I(N__62463));
    InMux I__15244 (
            .O(N__62472),
            .I(N__62460));
    LocalMux I__15243 (
            .O(N__62469),
            .I(N__62457));
    Span4Mux_v I__15242 (
            .O(N__62466),
            .I(N__62452));
    Span4Mux_v I__15241 (
            .O(N__62463),
            .I(N__62447));
    LocalMux I__15240 (
            .O(N__62460),
            .I(N__62447));
    Span4Mux_h I__15239 (
            .O(N__62457),
            .I(N__62444));
    InMux I__15238 (
            .O(N__62456),
            .I(N__62441));
    InMux I__15237 (
            .O(N__62455),
            .I(N__62438));
    Span4Mux_h I__15236 (
            .O(N__62452),
            .I(N__62433));
    Span4Mux_h I__15235 (
            .O(N__62447),
            .I(N__62433));
    Span4Mux_v I__15234 (
            .O(N__62444),
            .I(N__62428));
    LocalMux I__15233 (
            .O(N__62441),
            .I(N__62428));
    LocalMux I__15232 (
            .O(N__62438),
            .I(c_state_RNIEVJ7_22));
    Odrv4 I__15231 (
            .O(N__62433),
            .I(c_state_RNIEVJ7_22));
    Odrv4 I__15230 (
            .O(N__62428),
            .I(c_state_RNIEVJ7_22));
    InMux I__15229 (
            .O(N__62421),
            .I(N__62417));
    InMux I__15228 (
            .O(N__62420),
            .I(N__62414));
    LocalMux I__15227 (
            .O(N__62417),
            .I(N__62411));
    LocalMux I__15226 (
            .O(N__62414),
            .I(\I2C_top_level_inst1.s_load_rdata2 ));
    Odrv4 I__15225 (
            .O(N__62411),
            .I(\I2C_top_level_inst1.s_load_rdata2 ));
    InMux I__15224 (
            .O(N__62406),
            .I(N__62403));
    LocalMux I__15223 (
            .O(N__62403),
            .I(N__62399));
    InMux I__15222 (
            .O(N__62402),
            .I(N__62396));
    Span4Mux_v I__15221 (
            .O(N__62399),
            .I(N__62393));
    LocalMux I__15220 (
            .O(N__62396),
            .I(N__62390));
    Span4Mux_h I__15219 (
            .O(N__62393),
            .I(N__62387));
    Odrv4 I__15218 (
            .O(N__62390),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0 ));
    Odrv4 I__15217 (
            .O(N__62387),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0 ));
    InMux I__15216 (
            .O(N__62382),
            .I(N__62379));
    LocalMux I__15215 (
            .O(N__62379),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_27 ));
    CascadeMux I__15214 (
            .O(N__62376),
            .I(N__62373));
    InMux I__15213 (
            .O(N__62373),
            .I(N__62370));
    LocalMux I__15212 (
            .O(N__62370),
            .I(N__62364));
    InMux I__15211 (
            .O(N__62369),
            .I(N__62361));
    InMux I__15210 (
            .O(N__62368),
            .I(N__62358));
    InMux I__15209 (
            .O(N__62367),
            .I(N__62353));
    Span4Mux_v I__15208 (
            .O(N__62364),
            .I(N__62350));
    LocalMux I__15207 (
            .O(N__62361),
            .I(N__62347));
    LocalMux I__15206 (
            .O(N__62358),
            .I(N__62344));
    InMux I__15205 (
            .O(N__62357),
            .I(N__62341));
    InMux I__15204 (
            .O(N__62356),
            .I(N__62338));
    LocalMux I__15203 (
            .O(N__62353),
            .I(N__62333));
    Span4Mux_v I__15202 (
            .O(N__62350),
            .I(N__62330));
    Span4Mux_h I__15201 (
            .O(N__62347),
            .I(N__62327));
    Span4Mux_v I__15200 (
            .O(N__62344),
            .I(N__62320));
    LocalMux I__15199 (
            .O(N__62341),
            .I(N__62320));
    LocalMux I__15198 (
            .O(N__62338),
            .I(N__62320));
    InMux I__15197 (
            .O(N__62337),
            .I(N__62317));
    InMux I__15196 (
            .O(N__62336),
            .I(N__62314));
    Span4Mux_v I__15195 (
            .O(N__62333),
            .I(N__62311));
    Span4Mux_h I__15194 (
            .O(N__62330),
            .I(N__62306));
    Span4Mux_v I__15193 (
            .O(N__62327),
            .I(N__62306));
    Span4Mux_h I__15192 (
            .O(N__62320),
            .I(N__62303));
    LocalMux I__15191 (
            .O(N__62317),
            .I(N__62300));
    LocalMux I__15190 (
            .O(N__62314),
            .I(N__62295));
    Sp12to4 I__15189 (
            .O(N__62311),
            .I(N__62295));
    Span4Mux_h I__15188 (
            .O(N__62306),
            .I(N__62292));
    Span4Mux_v I__15187 (
            .O(N__62303),
            .I(N__62289));
    Span4Mux_v I__15186 (
            .O(N__62300),
            .I(N__62286));
    Span12Mux_h I__15185 (
            .O(N__62295),
            .I(N__62281));
    Sp12to4 I__15184 (
            .O(N__62292),
            .I(N__62281));
    Span4Mux_h I__15183 (
            .O(N__62289),
            .I(N__62276));
    Span4Mux_h I__15182 (
            .O(N__62286),
            .I(N__62276));
    Odrv12 I__15181 (
            .O(N__62281),
            .I(I2C_top_level_inst1_s_data_oreg_28));
    Odrv4 I__15180 (
            .O(N__62276),
            .I(I2C_top_level_inst1_s_data_oreg_28));
    InMux I__15179 (
            .O(N__62271),
            .I(N__62268));
    LocalMux I__15178 (
            .O(N__62268),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_28 ));
    InMux I__15177 (
            .O(N__62265),
            .I(N__62256));
    InMux I__15176 (
            .O(N__62264),
            .I(N__62253));
    InMux I__15175 (
            .O(N__62263),
            .I(N__62250));
    InMux I__15174 (
            .O(N__62262),
            .I(N__62247));
    InMux I__15173 (
            .O(N__62261),
            .I(N__62243));
    InMux I__15172 (
            .O(N__62260),
            .I(N__62240));
    InMux I__15171 (
            .O(N__62259),
            .I(N__62237));
    LocalMux I__15170 (
            .O(N__62256),
            .I(N__62234));
    LocalMux I__15169 (
            .O(N__62253),
            .I(N__62231));
    LocalMux I__15168 (
            .O(N__62250),
            .I(N__62226));
    LocalMux I__15167 (
            .O(N__62247),
            .I(N__62226));
    InMux I__15166 (
            .O(N__62246),
            .I(N__62223));
    LocalMux I__15165 (
            .O(N__62243),
            .I(N__62218));
    LocalMux I__15164 (
            .O(N__62240),
            .I(N__62218));
    LocalMux I__15163 (
            .O(N__62237),
            .I(N__62215));
    Sp12to4 I__15162 (
            .O(N__62234),
            .I(N__62212));
    Span4Mux_v I__15161 (
            .O(N__62231),
            .I(N__62209));
    Span4Mux_v I__15160 (
            .O(N__62226),
            .I(N__62206));
    LocalMux I__15159 (
            .O(N__62223),
            .I(N__62197));
    Span12Mux_v I__15158 (
            .O(N__62218),
            .I(N__62197));
    Span12Mux_v I__15157 (
            .O(N__62215),
            .I(N__62197));
    Span12Mux_s11_h I__15156 (
            .O(N__62212),
            .I(N__62197));
    Odrv4 I__15155 (
            .O(N__62209),
            .I(I2C_top_level_inst1_s_data_oreg_29));
    Odrv4 I__15154 (
            .O(N__62206),
            .I(I2C_top_level_inst1_s_data_oreg_29));
    Odrv12 I__15153 (
            .O(N__62197),
            .I(I2C_top_level_inst1_s_data_oreg_29));
    InMux I__15152 (
            .O(N__62190),
            .I(N__62187));
    LocalMux I__15151 (
            .O(N__62187),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_29 ));
    InMux I__15150 (
            .O(N__62184),
            .I(N__62180));
    CascadeMux I__15149 (
            .O(N__62183),
            .I(N__62176));
    LocalMux I__15148 (
            .O(N__62180),
            .I(N__62173));
    InMux I__15147 (
            .O(N__62179),
            .I(N__62170));
    InMux I__15146 (
            .O(N__62176),
            .I(N__62166));
    Span4Mux_v I__15145 (
            .O(N__62173),
            .I(N__62160));
    LocalMux I__15144 (
            .O(N__62170),
            .I(N__62160));
    InMux I__15143 (
            .O(N__62169),
            .I(N__62157));
    LocalMux I__15142 (
            .O(N__62166),
            .I(N__62154));
    InMux I__15141 (
            .O(N__62165),
            .I(N__62151));
    Span4Mux_h I__15140 (
            .O(N__62160),
            .I(N__62148));
    LocalMux I__15139 (
            .O(N__62157),
            .I(N__62144));
    Span4Mux_h I__15138 (
            .O(N__62154),
            .I(N__62139));
    LocalMux I__15137 (
            .O(N__62151),
            .I(N__62139));
    Span4Mux_v I__15136 (
            .O(N__62148),
            .I(N__62136));
    InMux I__15135 (
            .O(N__62147),
            .I(N__62133));
    Span4Mux_v I__15134 (
            .O(N__62144),
            .I(N__62129));
    Span4Mux_v I__15133 (
            .O(N__62139),
            .I(N__62126));
    Span4Mux_h I__15132 (
            .O(N__62136),
            .I(N__62120));
    LocalMux I__15131 (
            .O(N__62133),
            .I(N__62120));
    InMux I__15130 (
            .O(N__62132),
            .I(N__62117));
    Span4Mux_v I__15129 (
            .O(N__62129),
            .I(N__62114));
    Span4Mux_v I__15128 (
            .O(N__62126),
            .I(N__62111));
    InMux I__15127 (
            .O(N__62125),
            .I(N__62108));
    Span4Mux_h I__15126 (
            .O(N__62120),
            .I(N__62105));
    LocalMux I__15125 (
            .O(N__62117),
            .I(N__62102));
    Sp12to4 I__15124 (
            .O(N__62114),
            .I(N__62097));
    Sp12to4 I__15123 (
            .O(N__62111),
            .I(N__62097));
    LocalMux I__15122 (
            .O(N__62108),
            .I(N__62090));
    Span4Mux_v I__15121 (
            .O(N__62105),
            .I(N__62090));
    Span4Mux_v I__15120 (
            .O(N__62102),
            .I(N__62090));
    Span12Mux_h I__15119 (
            .O(N__62097),
            .I(N__62087));
    Span4Mux_h I__15118 (
            .O(N__62090),
            .I(N__62084));
    Odrv12 I__15117 (
            .O(N__62087),
            .I(I2C_top_level_inst1_s_data_oreg_30));
    Odrv4 I__15116 (
            .O(N__62084),
            .I(I2C_top_level_inst1_s_data_oreg_30));
    InMux I__15115 (
            .O(N__62079),
            .I(N__62076));
    LocalMux I__15114 (
            .O(N__62076),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_30 ));
    InMux I__15113 (
            .O(N__62073),
            .I(N__62067));
    InMux I__15112 (
            .O(N__62072),
            .I(N__62064));
    InMux I__15111 (
            .O(N__62071),
            .I(N__62061));
    InMux I__15110 (
            .O(N__62070),
            .I(N__62056));
    LocalMux I__15109 (
            .O(N__62067),
            .I(N__62051));
    LocalMux I__15108 (
            .O(N__62064),
            .I(N__62051));
    LocalMux I__15107 (
            .O(N__62061),
            .I(N__62048));
    CascadeMux I__15106 (
            .O(N__62060),
            .I(N__62045));
    InMux I__15105 (
            .O(N__62059),
            .I(N__62041));
    LocalMux I__15104 (
            .O(N__62056),
            .I(N__62038));
    Span4Mux_v I__15103 (
            .O(N__62051),
            .I(N__62033));
    Span4Mux_h I__15102 (
            .O(N__62048),
            .I(N__62033));
    InMux I__15101 (
            .O(N__62045),
            .I(N__62028));
    InMux I__15100 (
            .O(N__62044),
            .I(N__62028));
    LocalMux I__15099 (
            .O(N__62041),
            .I(N__62025));
    Span4Mux_v I__15098 (
            .O(N__62038),
            .I(N__62019));
    Span4Mux_h I__15097 (
            .O(N__62033),
            .I(N__62019));
    LocalMux I__15096 (
            .O(N__62028),
            .I(N__62016));
    Span12Mux_v I__15095 (
            .O(N__62025),
            .I(N__62013));
    InMux I__15094 (
            .O(N__62024),
            .I(N__62010));
    Span4Mux_h I__15093 (
            .O(N__62019),
            .I(N__62007));
    Span4Mux_h I__15092 (
            .O(N__62016),
            .I(N__62004));
    Span12Mux_h I__15091 (
            .O(N__62013),
            .I(N__62001));
    LocalMux I__15090 (
            .O(N__62010),
            .I(N__61994));
    Span4Mux_v I__15089 (
            .O(N__62007),
            .I(N__61994));
    Span4Mux_v I__15088 (
            .O(N__62004),
            .I(N__61994));
    Odrv12 I__15087 (
            .O(N__62001),
            .I(I2C_top_level_inst1_s_data_oreg_31));
    Odrv4 I__15086 (
            .O(N__61994),
            .I(I2C_top_level_inst1_s_data_oreg_31));
    InMux I__15085 (
            .O(N__61989),
            .I(N__61986));
    LocalMux I__15084 (
            .O(N__61986),
            .I(N__61983));
    Span4Mux_v I__15083 (
            .O(N__61983),
            .I(N__61980));
    Span4Mux_h I__15082 (
            .O(N__61980),
            .I(N__61977));
    Span4Mux_h I__15081 (
            .O(N__61977),
            .I(N__61974));
    Odrv4 I__15080 (
            .O(N__61974),
            .I(\I2C_top_level_inst1.s_sda_o_reg ));
    InMux I__15079 (
            .O(N__61971),
            .I(N__61965));
    InMux I__15078 (
            .O(N__61970),
            .I(N__61960));
    InMux I__15077 (
            .O(N__61969),
            .I(N__61956));
    InMux I__15076 (
            .O(N__61968),
            .I(N__61953));
    LocalMux I__15075 (
            .O(N__61965),
            .I(N__61950));
    InMux I__15074 (
            .O(N__61964),
            .I(N__61947));
    InMux I__15073 (
            .O(N__61963),
            .I(N__61944));
    LocalMux I__15072 (
            .O(N__61960),
            .I(N__61940));
    InMux I__15071 (
            .O(N__61959),
            .I(N__61937));
    LocalMux I__15070 (
            .O(N__61956),
            .I(N__61934));
    LocalMux I__15069 (
            .O(N__61953),
            .I(N__61931));
    Span4Mux_v I__15068 (
            .O(N__61950),
            .I(N__61927));
    LocalMux I__15067 (
            .O(N__61947),
            .I(N__61922));
    LocalMux I__15066 (
            .O(N__61944),
            .I(N__61922));
    InMux I__15065 (
            .O(N__61943),
            .I(N__61919));
    Span4Mux_v I__15064 (
            .O(N__61940),
            .I(N__61910));
    LocalMux I__15063 (
            .O(N__61937),
            .I(N__61910));
    Span4Mux_h I__15062 (
            .O(N__61934),
            .I(N__61910));
    Span4Mux_v I__15061 (
            .O(N__61931),
            .I(N__61910));
    InMux I__15060 (
            .O(N__61930),
            .I(N__61907));
    Sp12to4 I__15059 (
            .O(N__61927),
            .I(N__61904));
    Span12Mux_s9_v I__15058 (
            .O(N__61922),
            .I(N__61901));
    LocalMux I__15057 (
            .O(N__61919),
            .I(N__61898));
    Span4Mux_v I__15056 (
            .O(N__61910),
            .I(N__61895));
    LocalMux I__15055 (
            .O(N__61907),
            .I(N__61890));
    Span12Mux_h I__15054 (
            .O(N__61904),
            .I(N__61890));
    Span12Mux_h I__15053 (
            .O(N__61901),
            .I(N__61887));
    Odrv4 I__15052 (
            .O(N__61898),
            .I(I2C_top_level_inst1_s_data_oreg_0));
    Odrv4 I__15051 (
            .O(N__61895),
            .I(I2C_top_level_inst1_s_data_oreg_0));
    Odrv12 I__15050 (
            .O(N__61890),
            .I(I2C_top_level_inst1_s_data_oreg_0));
    Odrv12 I__15049 (
            .O(N__61887),
            .I(I2C_top_level_inst1_s_data_oreg_0));
    InMux I__15048 (
            .O(N__61878),
            .I(N__61875));
    LocalMux I__15047 (
            .O(N__61875),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_0 ));
    InMux I__15046 (
            .O(N__61872),
            .I(N__61868));
    InMux I__15045 (
            .O(N__61871),
            .I(N__61864));
    LocalMux I__15044 (
            .O(N__61868),
            .I(N__61856));
    InMux I__15043 (
            .O(N__61867),
            .I(N__61853));
    LocalMux I__15042 (
            .O(N__61864),
            .I(N__61850));
    InMux I__15041 (
            .O(N__61863),
            .I(N__61847));
    CascadeMux I__15040 (
            .O(N__61862),
            .I(N__61844));
    InMux I__15039 (
            .O(N__61861),
            .I(N__61841));
    InMux I__15038 (
            .O(N__61860),
            .I(N__61838));
    InMux I__15037 (
            .O(N__61859),
            .I(N__61835));
    Span4Mux_v I__15036 (
            .O(N__61856),
            .I(N__61832));
    LocalMux I__15035 (
            .O(N__61853),
            .I(N__61827));
    Span4Mux_v I__15034 (
            .O(N__61850),
            .I(N__61827));
    LocalMux I__15033 (
            .O(N__61847),
            .I(N__61824));
    InMux I__15032 (
            .O(N__61844),
            .I(N__61821));
    LocalMux I__15031 (
            .O(N__61841),
            .I(N__61817));
    LocalMux I__15030 (
            .O(N__61838),
            .I(N__61814));
    LocalMux I__15029 (
            .O(N__61835),
            .I(N__61811));
    Span4Mux_v I__15028 (
            .O(N__61832),
            .I(N__61808));
    Span4Mux_h I__15027 (
            .O(N__61827),
            .I(N__61803));
    Span4Mux_v I__15026 (
            .O(N__61824),
            .I(N__61803));
    LocalMux I__15025 (
            .O(N__61821),
            .I(N__61800));
    InMux I__15024 (
            .O(N__61820),
            .I(N__61797));
    Span4Mux_v I__15023 (
            .O(N__61817),
            .I(N__61794));
    Span4Mux_v I__15022 (
            .O(N__61814),
            .I(N__61791));
    Span4Mux_v I__15021 (
            .O(N__61811),
            .I(N__61788));
    Sp12to4 I__15020 (
            .O(N__61808),
            .I(N__61785));
    Span4Mux_h I__15019 (
            .O(N__61803),
            .I(N__61782));
    Span4Mux_h I__15018 (
            .O(N__61800),
            .I(N__61779));
    LocalMux I__15017 (
            .O(N__61797),
            .I(N__61776));
    Span4Mux_h I__15016 (
            .O(N__61794),
            .I(N__61773));
    Sp12to4 I__15015 (
            .O(N__61791),
            .I(N__61766));
    Sp12to4 I__15014 (
            .O(N__61788),
            .I(N__61766));
    Span12Mux_s10_h I__15013 (
            .O(N__61785),
            .I(N__61766));
    Span4Mux_v I__15012 (
            .O(N__61782),
            .I(N__61759));
    Span4Mux_v I__15011 (
            .O(N__61779),
            .I(N__61759));
    Span4Mux_h I__15010 (
            .O(N__61776),
            .I(N__61759));
    Odrv4 I__15009 (
            .O(N__61773),
            .I(I2C_top_level_inst1_s_data_oreg_1));
    Odrv12 I__15008 (
            .O(N__61766),
            .I(I2C_top_level_inst1_s_data_oreg_1));
    Odrv4 I__15007 (
            .O(N__61759),
            .I(I2C_top_level_inst1_s_data_oreg_1));
    InMux I__15006 (
            .O(N__61752),
            .I(N__61749));
    LocalMux I__15005 (
            .O(N__61749),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_1 ));
    InMux I__15004 (
            .O(N__61746),
            .I(N__61742));
    InMux I__15003 (
            .O(N__61745),
            .I(N__61739));
    LocalMux I__15002 (
            .O(N__61742),
            .I(N__61734));
    LocalMux I__15001 (
            .O(N__61739),
            .I(N__61731));
    InMux I__15000 (
            .O(N__61738),
            .I(N__61726));
    InMux I__14999 (
            .O(N__61737),
            .I(N__61723));
    Span4Mux_v I__14998 (
            .O(N__61734),
            .I(N__61720));
    Span4Mux_h I__14997 (
            .O(N__61731),
            .I(N__61716));
    InMux I__14996 (
            .O(N__61730),
            .I(N__61713));
    InMux I__14995 (
            .O(N__61729),
            .I(N__61708));
    LocalMux I__14994 (
            .O(N__61726),
            .I(N__61705));
    LocalMux I__14993 (
            .O(N__61723),
            .I(N__61700));
    Span4Mux_h I__14992 (
            .O(N__61720),
            .I(N__61700));
    InMux I__14991 (
            .O(N__61719),
            .I(N__61697));
    Span4Mux_v I__14990 (
            .O(N__61716),
            .I(N__61694));
    LocalMux I__14989 (
            .O(N__61713),
            .I(N__61691));
    CascadeMux I__14988 (
            .O(N__61712),
            .I(N__61688));
    InMux I__14987 (
            .O(N__61711),
            .I(N__61685));
    LocalMux I__14986 (
            .O(N__61708),
            .I(N__61682));
    Sp12to4 I__14985 (
            .O(N__61705),
            .I(N__61675));
    Sp12to4 I__14984 (
            .O(N__61700),
            .I(N__61675));
    LocalMux I__14983 (
            .O(N__61697),
            .I(N__61675));
    Span4Mux_h I__14982 (
            .O(N__61694),
            .I(N__61670));
    Span4Mux_h I__14981 (
            .O(N__61691),
            .I(N__61670));
    InMux I__14980 (
            .O(N__61688),
            .I(N__61667));
    LocalMux I__14979 (
            .O(N__61685),
            .I(N__61662));
    Sp12to4 I__14978 (
            .O(N__61682),
            .I(N__61662));
    Span12Mux_v I__14977 (
            .O(N__61675),
            .I(N__61659));
    Span4Mux_h I__14976 (
            .O(N__61670),
            .I(N__61656));
    LocalMux I__14975 (
            .O(N__61667),
            .I(I2C_top_level_inst1_s_data_oreg_2));
    Odrv12 I__14974 (
            .O(N__61662),
            .I(I2C_top_level_inst1_s_data_oreg_2));
    Odrv12 I__14973 (
            .O(N__61659),
            .I(I2C_top_level_inst1_s_data_oreg_2));
    Odrv4 I__14972 (
            .O(N__61656),
            .I(I2C_top_level_inst1_s_data_oreg_2));
    InMux I__14971 (
            .O(N__61647),
            .I(N__61641));
    InMux I__14970 (
            .O(N__61646),
            .I(N__61636));
    InMux I__14969 (
            .O(N__61645),
            .I(N__61633));
    InMux I__14968 (
            .O(N__61644),
            .I(N__61628));
    LocalMux I__14967 (
            .O(N__61641),
            .I(N__61625));
    InMux I__14966 (
            .O(N__61640),
            .I(N__61622));
    InMux I__14965 (
            .O(N__61639),
            .I(N__61619));
    LocalMux I__14964 (
            .O(N__61636),
            .I(N__61614));
    LocalMux I__14963 (
            .O(N__61633),
            .I(N__61614));
    CascadeMux I__14962 (
            .O(N__61632),
            .I(N__61610));
    InMux I__14961 (
            .O(N__61631),
            .I(N__61607));
    LocalMux I__14960 (
            .O(N__61628),
            .I(N__61604));
    Span4Mux_v I__14959 (
            .O(N__61625),
            .I(N__61599));
    LocalMux I__14958 (
            .O(N__61622),
            .I(N__61599));
    LocalMux I__14957 (
            .O(N__61619),
            .I(N__61596));
    Span4Mux_v I__14956 (
            .O(N__61614),
            .I(N__61593));
    InMux I__14955 (
            .O(N__61613),
            .I(N__61590));
    InMux I__14954 (
            .O(N__61610),
            .I(N__61587));
    LocalMux I__14953 (
            .O(N__61607),
            .I(N__61580));
    Span4Mux_v I__14952 (
            .O(N__61604),
            .I(N__61580));
    Span4Mux_v I__14951 (
            .O(N__61599),
            .I(N__61580));
    Span4Mux_v I__14950 (
            .O(N__61596),
            .I(N__61575));
    Span4Mux_h I__14949 (
            .O(N__61593),
            .I(N__61575));
    LocalMux I__14948 (
            .O(N__61590),
            .I(N__61572));
    LocalMux I__14947 (
            .O(N__61587),
            .I(N__61569));
    Span4Mux_h I__14946 (
            .O(N__61580),
            .I(N__61566));
    Span4Mux_h I__14945 (
            .O(N__61575),
            .I(N__61559));
    Span4Mux_v I__14944 (
            .O(N__61572),
            .I(N__61559));
    Span4Mux_v I__14943 (
            .O(N__61569),
            .I(N__61559));
    Sp12to4 I__14942 (
            .O(N__61566),
            .I(N__61554));
    Sp12to4 I__14941 (
            .O(N__61559),
            .I(N__61554));
    Odrv12 I__14940 (
            .O(N__61554),
            .I(I2C_top_level_inst1_s_data_oreg_19));
    InMux I__14939 (
            .O(N__61551),
            .I(N__61548));
    LocalMux I__14938 (
            .O(N__61548),
            .I(N__61541));
    InMux I__14937 (
            .O(N__61547),
            .I(N__61538));
    InMux I__14936 (
            .O(N__61546),
            .I(N__61535));
    InMux I__14935 (
            .O(N__61545),
            .I(N__61532));
    InMux I__14934 (
            .O(N__61544),
            .I(N__61527));
    Span4Mux_v I__14933 (
            .O(N__61541),
            .I(N__61522));
    LocalMux I__14932 (
            .O(N__61538),
            .I(N__61517));
    LocalMux I__14931 (
            .O(N__61535),
            .I(N__61517));
    LocalMux I__14930 (
            .O(N__61532),
            .I(N__61514));
    InMux I__14929 (
            .O(N__61531),
            .I(N__61511));
    InMux I__14928 (
            .O(N__61530),
            .I(N__61508));
    LocalMux I__14927 (
            .O(N__61527),
            .I(N__61505));
    InMux I__14926 (
            .O(N__61526),
            .I(N__61502));
    InMux I__14925 (
            .O(N__61525),
            .I(N__61499));
    Span4Mux_h I__14924 (
            .O(N__61522),
            .I(N__61494));
    Span4Mux_v I__14923 (
            .O(N__61517),
            .I(N__61494));
    Span4Mux_v I__14922 (
            .O(N__61514),
            .I(N__61491));
    LocalMux I__14921 (
            .O(N__61511),
            .I(N__61486));
    LocalMux I__14920 (
            .O(N__61508),
            .I(N__61486));
    Span4Mux_v I__14919 (
            .O(N__61505),
            .I(N__61483));
    LocalMux I__14918 (
            .O(N__61502),
            .I(N__61478));
    LocalMux I__14917 (
            .O(N__61499),
            .I(N__61478));
    Sp12to4 I__14916 (
            .O(N__61494),
            .I(N__61473));
    Sp12to4 I__14915 (
            .O(N__61491),
            .I(N__61473));
    Span4Mux_v I__14914 (
            .O(N__61486),
            .I(N__61468));
    Span4Mux_h I__14913 (
            .O(N__61483),
            .I(N__61468));
    Odrv4 I__14912 (
            .O(N__61478),
            .I(I2C_top_level_inst1_s_data_oreg_20));
    Odrv12 I__14911 (
            .O(N__61473),
            .I(I2C_top_level_inst1_s_data_oreg_20));
    Odrv4 I__14910 (
            .O(N__61468),
            .I(I2C_top_level_inst1_s_data_oreg_20));
    InMux I__14909 (
            .O(N__61461),
            .I(N__61458));
    LocalMux I__14908 (
            .O(N__61458),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_19 ));
    InMux I__14907 (
            .O(N__61455),
            .I(N__61452));
    LocalMux I__14906 (
            .O(N__61452),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_20 ));
    InMux I__14905 (
            .O(N__61449),
            .I(N__61444));
    CascadeMux I__14904 (
            .O(N__61448),
            .I(N__61441));
    InMux I__14903 (
            .O(N__61447),
            .I(N__61438));
    LocalMux I__14902 (
            .O(N__61444),
            .I(N__61431));
    InMux I__14901 (
            .O(N__61441),
            .I(N__61428));
    LocalMux I__14900 (
            .O(N__61438),
            .I(N__61425));
    InMux I__14899 (
            .O(N__61437),
            .I(N__61422));
    InMux I__14898 (
            .O(N__61436),
            .I(N__61418));
    InMux I__14897 (
            .O(N__61435),
            .I(N__61415));
    InMux I__14896 (
            .O(N__61434),
            .I(N__61412));
    Span4Mux_v I__14895 (
            .O(N__61431),
            .I(N__61407));
    LocalMux I__14894 (
            .O(N__61428),
            .I(N__61407));
    Span4Mux_h I__14893 (
            .O(N__61425),
            .I(N__61401));
    LocalMux I__14892 (
            .O(N__61422),
            .I(N__61401));
    InMux I__14891 (
            .O(N__61421),
            .I(N__61398));
    LocalMux I__14890 (
            .O(N__61418),
            .I(N__61395));
    LocalMux I__14889 (
            .O(N__61415),
            .I(N__61390));
    LocalMux I__14888 (
            .O(N__61412),
            .I(N__61390));
    Span4Mux_h I__14887 (
            .O(N__61407),
            .I(N__61387));
    InMux I__14886 (
            .O(N__61406),
            .I(N__61384));
    Span4Mux_h I__14885 (
            .O(N__61401),
            .I(N__61381));
    LocalMux I__14884 (
            .O(N__61398),
            .I(N__61376));
    Span4Mux_h I__14883 (
            .O(N__61395),
            .I(N__61376));
    Span4Mux_v I__14882 (
            .O(N__61390),
            .I(N__61371));
    Span4Mux_h I__14881 (
            .O(N__61387),
            .I(N__61371));
    LocalMux I__14880 (
            .O(N__61384),
            .I(I2C_top_level_inst1_s_data_oreg_21));
    Odrv4 I__14879 (
            .O(N__61381),
            .I(I2C_top_level_inst1_s_data_oreg_21));
    Odrv4 I__14878 (
            .O(N__61376),
            .I(I2C_top_level_inst1_s_data_oreg_21));
    Odrv4 I__14877 (
            .O(N__61371),
            .I(I2C_top_level_inst1_s_data_oreg_21));
    InMux I__14876 (
            .O(N__61362),
            .I(N__61359));
    LocalMux I__14875 (
            .O(N__61359),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_21 ));
    InMux I__14874 (
            .O(N__61356),
            .I(N__61349));
    InMux I__14873 (
            .O(N__61355),
            .I(N__61345));
    InMux I__14872 (
            .O(N__61354),
            .I(N__61342));
    InMux I__14871 (
            .O(N__61353),
            .I(N__61339));
    InMux I__14870 (
            .O(N__61352),
            .I(N__61336));
    LocalMux I__14869 (
            .O(N__61349),
            .I(N__61333));
    InMux I__14868 (
            .O(N__61348),
            .I(N__61330));
    LocalMux I__14867 (
            .O(N__61345),
            .I(N__61327));
    LocalMux I__14866 (
            .O(N__61342),
            .I(N__61320));
    LocalMux I__14865 (
            .O(N__61339),
            .I(N__61320));
    LocalMux I__14864 (
            .O(N__61336),
            .I(N__61320));
    Span4Mux_v I__14863 (
            .O(N__61333),
            .I(N__61311));
    LocalMux I__14862 (
            .O(N__61330),
            .I(N__61311));
    Span4Mux_v I__14861 (
            .O(N__61327),
            .I(N__61311));
    Span4Mux_v I__14860 (
            .O(N__61320),
            .I(N__61307));
    InMux I__14859 (
            .O(N__61319),
            .I(N__61304));
    InMux I__14858 (
            .O(N__61318),
            .I(N__61301));
    Span4Mux_h I__14857 (
            .O(N__61311),
            .I(N__61298));
    InMux I__14856 (
            .O(N__61310),
            .I(N__61295));
    Span4Mux_h I__14855 (
            .O(N__61307),
            .I(N__61290));
    LocalMux I__14854 (
            .O(N__61304),
            .I(N__61290));
    LocalMux I__14853 (
            .O(N__61301),
            .I(N__61287));
    Span4Mux_h I__14852 (
            .O(N__61298),
            .I(N__61284));
    LocalMux I__14851 (
            .O(N__61295),
            .I(N__61281));
    Span4Mux_v I__14850 (
            .O(N__61290),
            .I(N__61276));
    Span4Mux_h I__14849 (
            .O(N__61287),
            .I(N__61276));
    Span4Mux_v I__14848 (
            .O(N__61284),
            .I(N__61273));
    Span4Mux_h I__14847 (
            .O(N__61281),
            .I(N__61270));
    Span4Mux_v I__14846 (
            .O(N__61276),
            .I(N__61267));
    Odrv4 I__14845 (
            .O(N__61273),
            .I(I2C_top_level_inst1_s_data_oreg_22));
    Odrv4 I__14844 (
            .O(N__61270),
            .I(I2C_top_level_inst1_s_data_oreg_22));
    Odrv4 I__14843 (
            .O(N__61267),
            .I(I2C_top_level_inst1_s_data_oreg_22));
    InMux I__14842 (
            .O(N__61260),
            .I(N__61257));
    LocalMux I__14841 (
            .O(N__61257),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_22 ));
    InMux I__14840 (
            .O(N__61254),
            .I(N__61249));
    InMux I__14839 (
            .O(N__61253),
            .I(N__61243));
    CascadeMux I__14838 (
            .O(N__61252),
            .I(N__61239));
    LocalMux I__14837 (
            .O(N__61249),
            .I(N__61236));
    InMux I__14836 (
            .O(N__61248),
            .I(N__61233));
    InMux I__14835 (
            .O(N__61247),
            .I(N__61230));
    InMux I__14834 (
            .O(N__61246),
            .I(N__61226));
    LocalMux I__14833 (
            .O(N__61243),
            .I(N__61223));
    InMux I__14832 (
            .O(N__61242),
            .I(N__61220));
    InMux I__14831 (
            .O(N__61239),
            .I(N__61217));
    Span4Mux_v I__14830 (
            .O(N__61236),
            .I(N__61212));
    LocalMux I__14829 (
            .O(N__61233),
            .I(N__61212));
    LocalMux I__14828 (
            .O(N__61230),
            .I(N__61209));
    InMux I__14827 (
            .O(N__61229),
            .I(N__61206));
    LocalMux I__14826 (
            .O(N__61226),
            .I(N__61203));
    Span4Mux_v I__14825 (
            .O(N__61223),
            .I(N__61200));
    LocalMux I__14824 (
            .O(N__61220),
            .I(N__61197));
    LocalMux I__14823 (
            .O(N__61217),
            .I(N__61194));
    Span4Mux_v I__14822 (
            .O(N__61212),
            .I(N__61188));
    Span4Mux_v I__14821 (
            .O(N__61209),
            .I(N__61188));
    LocalMux I__14820 (
            .O(N__61206),
            .I(N__61185));
    Span4Mux_v I__14819 (
            .O(N__61203),
            .I(N__61182));
    Span4Mux_h I__14818 (
            .O(N__61200),
            .I(N__61177));
    Span4Mux_v I__14817 (
            .O(N__61197),
            .I(N__61177));
    Span4Mux_v I__14816 (
            .O(N__61194),
            .I(N__61174));
    InMux I__14815 (
            .O(N__61193),
            .I(N__61171));
    Span4Mux_h I__14814 (
            .O(N__61188),
            .I(N__61166));
    Span4Mux_v I__14813 (
            .O(N__61185),
            .I(N__61166));
    Span4Mux_h I__14812 (
            .O(N__61182),
            .I(N__61163));
    Span4Mux_h I__14811 (
            .O(N__61177),
            .I(N__61158));
    Span4Mux_h I__14810 (
            .O(N__61174),
            .I(N__61158));
    LocalMux I__14809 (
            .O(N__61171),
            .I(N__61155));
    Sp12to4 I__14808 (
            .O(N__61166),
            .I(N__61152));
    Span4Mux_h I__14807 (
            .O(N__61163),
            .I(N__61149));
    Span4Mux_h I__14806 (
            .O(N__61158),
            .I(N__61146));
    Odrv12 I__14805 (
            .O(N__61155),
            .I(I2C_top_level_inst1_s_data_oreg_23));
    Odrv12 I__14804 (
            .O(N__61152),
            .I(I2C_top_level_inst1_s_data_oreg_23));
    Odrv4 I__14803 (
            .O(N__61149),
            .I(I2C_top_level_inst1_s_data_oreg_23));
    Odrv4 I__14802 (
            .O(N__61146),
            .I(I2C_top_level_inst1_s_data_oreg_23));
    InMux I__14801 (
            .O(N__61137),
            .I(N__61134));
    LocalMux I__14800 (
            .O(N__61134),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_23 ));
    InMux I__14799 (
            .O(N__61131),
            .I(N__61127));
    InMux I__14798 (
            .O(N__61130),
            .I(N__61121));
    LocalMux I__14797 (
            .O(N__61127),
            .I(N__61118));
    InMux I__14796 (
            .O(N__61126),
            .I(N__61114));
    InMux I__14795 (
            .O(N__61125),
            .I(N__61110));
    InMux I__14794 (
            .O(N__61124),
            .I(N__61107));
    LocalMux I__14793 (
            .O(N__61121),
            .I(N__61104));
    Span4Mux_v I__14792 (
            .O(N__61118),
            .I(N__61100));
    InMux I__14791 (
            .O(N__61117),
            .I(N__61097));
    LocalMux I__14790 (
            .O(N__61114),
            .I(N__61094));
    InMux I__14789 (
            .O(N__61113),
            .I(N__61091));
    LocalMux I__14788 (
            .O(N__61110),
            .I(N__61088));
    LocalMux I__14787 (
            .O(N__61107),
            .I(N__61085));
    Span4Mux_h I__14786 (
            .O(N__61104),
            .I(N__61082));
    InMux I__14785 (
            .O(N__61103),
            .I(N__61079));
    Span4Mux_h I__14784 (
            .O(N__61100),
            .I(N__61076));
    LocalMux I__14783 (
            .O(N__61097),
            .I(N__61073));
    Span4Mux_v I__14782 (
            .O(N__61094),
            .I(N__61070));
    LocalMux I__14781 (
            .O(N__61091),
            .I(N__61063));
    Span4Mux_v I__14780 (
            .O(N__61088),
            .I(N__61063));
    Span4Mux_v I__14779 (
            .O(N__61085),
            .I(N__61063));
    Span4Mux_h I__14778 (
            .O(N__61082),
            .I(N__61060));
    LocalMux I__14777 (
            .O(N__61079),
            .I(N__61057));
    Sp12to4 I__14776 (
            .O(N__61076),
            .I(N__61054));
    Span4Mux_v I__14775 (
            .O(N__61073),
            .I(N__61051));
    Span4Mux_h I__14774 (
            .O(N__61070),
            .I(N__61048));
    Span4Mux_h I__14773 (
            .O(N__61063),
            .I(N__61045));
    Sp12to4 I__14772 (
            .O(N__61060),
            .I(N__61038));
    Sp12to4 I__14771 (
            .O(N__61057),
            .I(N__61038));
    Span12Mux_v I__14770 (
            .O(N__61054),
            .I(N__61038));
    Span4Mux_v I__14769 (
            .O(N__61051),
            .I(N__61033));
    Span4Mux_h I__14768 (
            .O(N__61048),
            .I(N__61033));
    Odrv4 I__14767 (
            .O(N__61045),
            .I(I2C_top_level_inst1_s_data_oreg_24));
    Odrv12 I__14766 (
            .O(N__61038),
            .I(I2C_top_level_inst1_s_data_oreg_24));
    Odrv4 I__14765 (
            .O(N__61033),
            .I(I2C_top_level_inst1_s_data_oreg_24));
    InMux I__14764 (
            .O(N__61026),
            .I(N__61023));
    LocalMux I__14763 (
            .O(N__61023),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_24 ));
    CascadeMux I__14762 (
            .O(N__61020),
            .I(N__61015));
    InMux I__14761 (
            .O(N__61019),
            .I(N__61010));
    InMux I__14760 (
            .O(N__61018),
            .I(N__61007));
    InMux I__14759 (
            .O(N__61015),
            .I(N__61004));
    InMux I__14758 (
            .O(N__61014),
            .I(N__61001));
    InMux I__14757 (
            .O(N__61013),
            .I(N__60997));
    LocalMux I__14756 (
            .O(N__61010),
            .I(N__60994));
    LocalMux I__14755 (
            .O(N__61007),
            .I(N__60991));
    LocalMux I__14754 (
            .O(N__61004),
            .I(N__60988));
    LocalMux I__14753 (
            .O(N__61001),
            .I(N__60985));
    InMux I__14752 (
            .O(N__61000),
            .I(N__60982));
    LocalMux I__14751 (
            .O(N__60997),
            .I(N__60977));
    Span4Mux_v I__14750 (
            .O(N__60994),
            .I(N__60972));
    Span4Mux_v I__14749 (
            .O(N__60991),
            .I(N__60972));
    Span4Mux_v I__14748 (
            .O(N__60988),
            .I(N__60967));
    Span4Mux_v I__14747 (
            .O(N__60985),
            .I(N__60967));
    LocalMux I__14746 (
            .O(N__60982),
            .I(N__60964));
    InMux I__14745 (
            .O(N__60981),
            .I(N__60961));
    InMux I__14744 (
            .O(N__60980),
            .I(N__60958));
    Span4Mux_h I__14743 (
            .O(N__60977),
            .I(N__60955));
    Span4Mux_h I__14742 (
            .O(N__60972),
            .I(N__60952));
    Sp12to4 I__14741 (
            .O(N__60967),
            .I(N__60949));
    Span4Mux_v I__14740 (
            .O(N__60964),
            .I(N__60946));
    LocalMux I__14739 (
            .O(N__60961),
            .I(N__60939));
    LocalMux I__14738 (
            .O(N__60958),
            .I(N__60939));
    Span4Mux_v I__14737 (
            .O(N__60955),
            .I(N__60939));
    Sp12to4 I__14736 (
            .O(N__60952),
            .I(N__60934));
    Span12Mux_h I__14735 (
            .O(N__60949),
            .I(N__60934));
    Odrv4 I__14734 (
            .O(N__60946),
            .I(I2C_top_level_inst1_s_data_oreg_25));
    Odrv4 I__14733 (
            .O(N__60939),
            .I(I2C_top_level_inst1_s_data_oreg_25));
    Odrv12 I__14732 (
            .O(N__60934),
            .I(I2C_top_level_inst1_s_data_oreg_25));
    InMux I__14731 (
            .O(N__60927),
            .I(N__60924));
    LocalMux I__14730 (
            .O(N__60924),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_25 ));
    InMux I__14729 (
            .O(N__60921),
            .I(N__60918));
    LocalMux I__14728 (
            .O(N__60918),
            .I(N__60915));
    Span4Mux_h I__14727 (
            .O(N__60915),
            .I(N__60909));
    InMux I__14726 (
            .O(N__60914),
            .I(N__60906));
    InMux I__14725 (
            .O(N__60913),
            .I(N__60902));
    InMux I__14724 (
            .O(N__60912),
            .I(N__60898));
    Span4Mux_h I__14723 (
            .O(N__60909),
            .I(N__60892));
    LocalMux I__14722 (
            .O(N__60906),
            .I(N__60892));
    InMux I__14721 (
            .O(N__60905),
            .I(N__60889));
    LocalMux I__14720 (
            .O(N__60902),
            .I(N__60886));
    InMux I__14719 (
            .O(N__60901),
            .I(N__60883));
    LocalMux I__14718 (
            .O(N__60898),
            .I(N__60880));
    InMux I__14717 (
            .O(N__60897),
            .I(N__60877));
    Span4Mux_v I__14716 (
            .O(N__60892),
            .I(N__60872));
    LocalMux I__14715 (
            .O(N__60889),
            .I(N__60872));
    Span4Mux_h I__14714 (
            .O(N__60886),
            .I(N__60869));
    LocalMux I__14713 (
            .O(N__60883),
            .I(N__60866));
    Span4Mux_v I__14712 (
            .O(N__60880),
            .I(N__60863));
    LocalMux I__14711 (
            .O(N__60877),
            .I(N__60860));
    Span4Mux_h I__14710 (
            .O(N__60872),
            .I(N__60857));
    Span4Mux_v I__14709 (
            .O(N__60869),
            .I(N__60850));
    Span4Mux_v I__14708 (
            .O(N__60866),
            .I(N__60850));
    Span4Mux_v I__14707 (
            .O(N__60863),
            .I(N__60850));
    Span4Mux_h I__14706 (
            .O(N__60860),
            .I(N__60846));
    Sp12to4 I__14705 (
            .O(N__60857),
            .I(N__60843));
    Sp12to4 I__14704 (
            .O(N__60850),
            .I(N__60840));
    InMux I__14703 (
            .O(N__60849),
            .I(N__60837));
    Span4Mux_v I__14702 (
            .O(N__60846),
            .I(N__60834));
    Span12Mux_v I__14701 (
            .O(N__60843),
            .I(N__60829));
    Span12Mux_h I__14700 (
            .O(N__60840),
            .I(N__60829));
    LocalMux I__14699 (
            .O(N__60837),
            .I(I2C_top_level_inst1_s_data_oreg_26));
    Odrv4 I__14698 (
            .O(N__60834),
            .I(I2C_top_level_inst1_s_data_oreg_26));
    Odrv12 I__14697 (
            .O(N__60829),
            .I(I2C_top_level_inst1_s_data_oreg_26));
    InMux I__14696 (
            .O(N__60822),
            .I(N__60819));
    LocalMux I__14695 (
            .O(N__60819),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_26 ));
    CascadeMux I__14694 (
            .O(N__60816),
            .I(N__60813));
    InMux I__14693 (
            .O(N__60813),
            .I(N__60810));
    LocalMux I__14692 (
            .O(N__60810),
            .I(N__60807));
    Span4Mux_v I__14691 (
            .O(N__60807),
            .I(N__60802));
    InMux I__14690 (
            .O(N__60806),
            .I(N__60799));
    InMux I__14689 (
            .O(N__60805),
            .I(N__60794));
    Span4Mux_h I__14688 (
            .O(N__60802),
            .I(N__60791));
    LocalMux I__14687 (
            .O(N__60799),
            .I(N__60788));
    InMux I__14686 (
            .O(N__60798),
            .I(N__60783));
    InMux I__14685 (
            .O(N__60797),
            .I(N__60780));
    LocalMux I__14684 (
            .O(N__60794),
            .I(N__60777));
    Span4Mux_v I__14683 (
            .O(N__60791),
            .I(N__60771));
    Span4Mux_h I__14682 (
            .O(N__60788),
            .I(N__60771));
    InMux I__14681 (
            .O(N__60787),
            .I(N__60768));
    InMux I__14680 (
            .O(N__60786),
            .I(N__60765));
    LocalMux I__14679 (
            .O(N__60783),
            .I(N__60762));
    LocalMux I__14678 (
            .O(N__60780),
            .I(N__60759));
    Span4Mux_v I__14677 (
            .O(N__60777),
            .I(N__60756));
    InMux I__14676 (
            .O(N__60776),
            .I(N__60753));
    Span4Mux_v I__14675 (
            .O(N__60771),
            .I(N__60746));
    LocalMux I__14674 (
            .O(N__60768),
            .I(N__60746));
    LocalMux I__14673 (
            .O(N__60765),
            .I(N__60746));
    Span4Mux_h I__14672 (
            .O(N__60762),
            .I(N__60743));
    Span4Mux_v I__14671 (
            .O(N__60759),
            .I(N__60740));
    Span4Mux_h I__14670 (
            .O(N__60756),
            .I(N__60737));
    LocalMux I__14669 (
            .O(N__60753),
            .I(N__60734));
    Span4Mux_h I__14668 (
            .O(N__60746),
            .I(N__60731));
    Span4Mux_v I__14667 (
            .O(N__60743),
            .I(N__60728));
    Span4Mux_v I__14666 (
            .O(N__60740),
            .I(N__60723));
    Span4Mux_h I__14665 (
            .O(N__60737),
            .I(N__60723));
    Odrv4 I__14664 (
            .O(N__60734),
            .I(I2C_top_level_inst1_s_data_oreg_27));
    Odrv4 I__14663 (
            .O(N__60731),
            .I(I2C_top_level_inst1_s_data_oreg_27));
    Odrv4 I__14662 (
            .O(N__60728),
            .I(I2C_top_level_inst1_s_data_oreg_27));
    Odrv4 I__14661 (
            .O(N__60723),
            .I(I2C_top_level_inst1_s_data_oreg_27));
    InMux I__14660 (
            .O(N__60714),
            .I(N__60711));
    LocalMux I__14659 (
            .O(N__60711),
            .I(N__60706));
    InMux I__14658 (
            .O(N__60710),
            .I(N__60703));
    CascadeMux I__14657 (
            .O(N__60709),
            .I(N__60700));
    Span4Mux_h I__14656 (
            .O(N__60706),
            .I(N__60697));
    LocalMux I__14655 (
            .O(N__60703),
            .I(N__60694));
    InMux I__14654 (
            .O(N__60700),
            .I(N__60691));
    Span4Mux_h I__14653 (
            .O(N__60697),
            .I(N__60688));
    Span4Mux_h I__14652 (
            .O(N__60694),
            .I(N__60683));
    LocalMux I__14651 (
            .O(N__60691),
            .I(N__60683));
    Odrv4 I__14650 (
            .O(N__60688),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_1));
    Odrv4 I__14649 (
            .O(N__60683),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_1));
    CascadeMux I__14648 (
            .O(N__60678),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_1_cascade_ ));
    InMux I__14647 (
            .O(N__60675),
            .I(N__60672));
    LocalMux I__14646 (
            .O(N__60672),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_1 ));
    CascadeMux I__14645 (
            .O(N__60669),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2QZ0Z5_cascade_ ));
    InMux I__14644 (
            .O(N__60666),
            .I(N__60663));
    LocalMux I__14643 (
            .O(N__60663),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1 ));
    CascadeMux I__14642 (
            .O(N__60660),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_cascade_ ));
    InMux I__14641 (
            .O(N__60657),
            .I(N__60654));
    LocalMux I__14640 (
            .O(N__60654),
            .I(N__60651));
    Span4Mux_h I__14639 (
            .O(N__60651),
            .I(N__60648));
    Odrv4 I__14638 (
            .O(N__60648),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_1 ));
    InMux I__14637 (
            .O(N__60645),
            .I(N__60642));
    LocalMux I__14636 (
            .O(N__60642),
            .I(N__60637));
    InMux I__14635 (
            .O(N__60641),
            .I(N__60634));
    InMux I__14634 (
            .O(N__60640),
            .I(N__60631));
    Span4Mux_v I__14633 (
            .O(N__60637),
            .I(N__60626));
    LocalMux I__14632 (
            .O(N__60634),
            .I(N__60626));
    LocalMux I__14631 (
            .O(N__60631),
            .I(N__60623));
    Odrv4 I__14630 (
            .O(N__60626),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_0));
    Odrv4 I__14629 (
            .O(N__60623),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_0));
    InMux I__14628 (
            .O(N__60618),
            .I(N__60609));
    InMux I__14627 (
            .O(N__60617),
            .I(N__60606));
    InMux I__14626 (
            .O(N__60616),
            .I(N__60599));
    InMux I__14625 (
            .O(N__60615),
            .I(N__60599));
    InMux I__14624 (
            .O(N__60614),
            .I(N__60592));
    InMux I__14623 (
            .O(N__60613),
            .I(N__60592));
    InMux I__14622 (
            .O(N__60612),
            .I(N__60586));
    LocalMux I__14621 (
            .O(N__60609),
            .I(N__60581));
    LocalMux I__14620 (
            .O(N__60606),
            .I(N__60581));
    InMux I__14619 (
            .O(N__60605),
            .I(N__60578));
    InMux I__14618 (
            .O(N__60604),
            .I(N__60575));
    LocalMux I__14617 (
            .O(N__60599),
            .I(N__60572));
    InMux I__14616 (
            .O(N__60598),
            .I(N__60569));
    InMux I__14615 (
            .O(N__60597),
            .I(N__60566));
    LocalMux I__14614 (
            .O(N__60592),
            .I(N__60562));
    InMux I__14613 (
            .O(N__60591),
            .I(N__60559));
    InMux I__14612 (
            .O(N__60590),
            .I(N__60552));
    InMux I__14611 (
            .O(N__60589),
            .I(N__60552));
    LocalMux I__14610 (
            .O(N__60586),
            .I(N__60549));
    Span4Mux_h I__14609 (
            .O(N__60581),
            .I(N__60544));
    LocalMux I__14608 (
            .O(N__60578),
            .I(N__60544));
    LocalMux I__14607 (
            .O(N__60575),
            .I(N__60541));
    Span4Mux_v I__14606 (
            .O(N__60572),
            .I(N__60535));
    LocalMux I__14605 (
            .O(N__60569),
            .I(N__60535));
    LocalMux I__14604 (
            .O(N__60566),
            .I(N__60532));
    InMux I__14603 (
            .O(N__60565),
            .I(N__60529));
    Span4Mux_h I__14602 (
            .O(N__60562),
            .I(N__60524));
    LocalMux I__14601 (
            .O(N__60559),
            .I(N__60524));
    InMux I__14600 (
            .O(N__60558),
            .I(N__60521));
    InMux I__14599 (
            .O(N__60557),
            .I(N__60518));
    LocalMux I__14598 (
            .O(N__60552),
            .I(N__60512));
    Span4Mux_v I__14597 (
            .O(N__60549),
            .I(N__60507));
    Span4Mux_v I__14596 (
            .O(N__60544),
            .I(N__60507));
    Span4Mux_h I__14595 (
            .O(N__60541),
            .I(N__60504));
    InMux I__14594 (
            .O(N__60540),
            .I(N__60501));
    Span4Mux_h I__14593 (
            .O(N__60535),
            .I(N__60496));
    Span4Mux_v I__14592 (
            .O(N__60532),
            .I(N__60496));
    LocalMux I__14591 (
            .O(N__60529),
            .I(N__60489));
    Span4Mux_h I__14590 (
            .O(N__60524),
            .I(N__60489));
    LocalMux I__14589 (
            .O(N__60521),
            .I(N__60489));
    LocalMux I__14588 (
            .O(N__60518),
            .I(N__60486));
    InMux I__14587 (
            .O(N__60517),
            .I(N__60483));
    InMux I__14586 (
            .O(N__60516),
            .I(N__60478));
    InMux I__14585 (
            .O(N__60515),
            .I(N__60478));
    Span4Mux_v I__14584 (
            .O(N__60512),
            .I(N__60475));
    Span4Mux_h I__14583 (
            .O(N__60507),
            .I(N__60469));
    Span4Mux_h I__14582 (
            .O(N__60504),
            .I(N__60464));
    LocalMux I__14581 (
            .O(N__60501),
            .I(N__60464));
    Span4Mux_h I__14580 (
            .O(N__60496),
            .I(N__60461));
    Span4Mux_v I__14579 (
            .O(N__60489),
            .I(N__60456));
    Span4Mux_h I__14578 (
            .O(N__60486),
            .I(N__60456));
    LocalMux I__14577 (
            .O(N__60483),
            .I(N__60451));
    LocalMux I__14576 (
            .O(N__60478),
            .I(N__60451));
    Sp12to4 I__14575 (
            .O(N__60475),
            .I(N__60448));
    InMux I__14574 (
            .O(N__60474),
            .I(N__60445));
    InMux I__14573 (
            .O(N__60473),
            .I(N__60440));
    InMux I__14572 (
            .O(N__60472),
            .I(N__60440));
    Span4Mux_h I__14571 (
            .O(N__60469),
            .I(N__60435));
    Span4Mux_v I__14570 (
            .O(N__60464),
            .I(N__60435));
    Span4Mux_h I__14569 (
            .O(N__60461),
            .I(N__60430));
    Span4Mux_h I__14568 (
            .O(N__60456),
            .I(N__60430));
    Span12Mux_v I__14567 (
            .O(N__60451),
            .I(N__60427));
    Span12Mux_h I__14566 (
            .O(N__60448),
            .I(N__60420));
    LocalMux I__14565 (
            .O(N__60445),
            .I(N__60420));
    LocalMux I__14564 (
            .O(N__60440),
            .I(N__60420));
    Odrv4 I__14563 (
            .O(N__60435),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340 ));
    Odrv4 I__14562 (
            .O(N__60430),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340 ));
    Odrv12 I__14561 (
            .O(N__60427),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340 ));
    Odrv12 I__14560 (
            .O(N__60420),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340 ));
    CascadeMux I__14559 (
            .O(N__60411),
            .I(N__60408));
    InMux I__14558 (
            .O(N__60408),
            .I(N__60405));
    LocalMux I__14557 (
            .O(N__60405),
            .I(N__60402));
    Span4Mux_v I__14556 (
            .O(N__60402),
            .I(N__60399));
    Span4Mux_h I__14555 (
            .O(N__60399),
            .I(N__60396));
    Odrv4 I__14554 (
            .O(N__60396),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_0 ));
    InMux I__14553 (
            .O(N__60393),
            .I(N__60390));
    LocalMux I__14552 (
            .O(N__60390),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_0 ));
    InMux I__14551 (
            .O(N__60387),
            .I(N__60369));
    InMux I__14550 (
            .O(N__60386),
            .I(N__60369));
    InMux I__14549 (
            .O(N__60385),
            .I(N__60364));
    InMux I__14548 (
            .O(N__60384),
            .I(N__60364));
    InMux I__14547 (
            .O(N__60383),
            .I(N__60359));
    InMux I__14546 (
            .O(N__60382),
            .I(N__60359));
    InMux I__14545 (
            .O(N__60381),
            .I(N__60350));
    InMux I__14544 (
            .O(N__60380),
            .I(N__60347));
    InMux I__14543 (
            .O(N__60379),
            .I(N__60340));
    InMux I__14542 (
            .O(N__60378),
            .I(N__60340));
    InMux I__14541 (
            .O(N__60377),
            .I(N__60335));
    InMux I__14540 (
            .O(N__60376),
            .I(N__60335));
    InMux I__14539 (
            .O(N__60375),
            .I(N__60330));
    InMux I__14538 (
            .O(N__60374),
            .I(N__60330));
    LocalMux I__14537 (
            .O(N__60369),
            .I(N__60325));
    LocalMux I__14536 (
            .O(N__60364),
            .I(N__60320));
    LocalMux I__14535 (
            .O(N__60359),
            .I(N__60320));
    InMux I__14534 (
            .O(N__60358),
            .I(N__60317));
    InMux I__14533 (
            .O(N__60357),
            .I(N__60312));
    InMux I__14532 (
            .O(N__60356),
            .I(N__60312));
    InMux I__14531 (
            .O(N__60355),
            .I(N__60307));
    InMux I__14530 (
            .O(N__60354),
            .I(N__60307));
    InMux I__14529 (
            .O(N__60353),
            .I(N__60304));
    LocalMux I__14528 (
            .O(N__60350),
            .I(N__60299));
    LocalMux I__14527 (
            .O(N__60347),
            .I(N__60299));
    InMux I__14526 (
            .O(N__60346),
            .I(N__60294));
    InMux I__14525 (
            .O(N__60345),
            .I(N__60294));
    LocalMux I__14524 (
            .O(N__60340),
            .I(N__60287));
    LocalMux I__14523 (
            .O(N__60335),
            .I(N__60287));
    LocalMux I__14522 (
            .O(N__60330),
            .I(N__60287));
    InMux I__14521 (
            .O(N__60329),
            .I(N__60282));
    InMux I__14520 (
            .O(N__60328),
            .I(N__60282));
    Span4Mux_h I__14519 (
            .O(N__60325),
            .I(N__60277));
    Span4Mux_v I__14518 (
            .O(N__60320),
            .I(N__60277));
    LocalMux I__14517 (
            .O(N__60317),
            .I(N__60272));
    LocalMux I__14516 (
            .O(N__60312),
            .I(N__60272));
    LocalMux I__14515 (
            .O(N__60307),
            .I(N__60269));
    LocalMux I__14514 (
            .O(N__60304),
            .I(N__60266));
    Span4Mux_v I__14513 (
            .O(N__60299),
            .I(N__60263));
    LocalMux I__14512 (
            .O(N__60294),
            .I(N__60260));
    Span4Mux_v I__14511 (
            .O(N__60287),
            .I(N__60257));
    LocalMux I__14510 (
            .O(N__60282),
            .I(N__60254));
    Span4Mux_h I__14509 (
            .O(N__60277),
            .I(N__60249));
    Span4Mux_v I__14508 (
            .O(N__60272),
            .I(N__60249));
    Sp12to4 I__14507 (
            .O(N__60269),
            .I(N__60246));
    Span12Mux_v I__14506 (
            .O(N__60266),
            .I(N__60243));
    Span4Mux_v I__14505 (
            .O(N__60263),
            .I(N__60240));
    Sp12to4 I__14504 (
            .O(N__60260),
            .I(N__60235));
    Sp12to4 I__14503 (
            .O(N__60257),
            .I(N__60235));
    Span4Mux_h I__14502 (
            .O(N__60254),
            .I(N__60230));
    Span4Mux_h I__14501 (
            .O(N__60249),
            .I(N__60230));
    Odrv12 I__14500 (
            .O(N__60246),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ));
    Odrv12 I__14499 (
            .O(N__60243),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ));
    Odrv4 I__14498 (
            .O(N__60240),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ));
    Odrv12 I__14497 (
            .O(N__60235),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ));
    Odrv4 I__14496 (
            .O(N__60230),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ));
    CascadeMux I__14495 (
            .O(N__60219),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2QZ0Z5_cascade_ ));
    InMux I__14494 (
            .O(N__60216),
            .I(N__60213));
    LocalMux I__14493 (
            .O(N__60213),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0 ));
    CascadeMux I__14492 (
            .O(N__60210),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0_cascade_ ));
    InMux I__14491 (
            .O(N__60207),
            .I(N__60197));
    InMux I__14490 (
            .O(N__60206),
            .I(N__60197));
    InMux I__14489 (
            .O(N__60205),
            .I(N__60188));
    InMux I__14488 (
            .O(N__60204),
            .I(N__60188));
    InMux I__14487 (
            .O(N__60203),
            .I(N__60181));
    InMux I__14486 (
            .O(N__60202),
            .I(N__60181));
    LocalMux I__14485 (
            .O(N__60197),
            .I(N__60178));
    InMux I__14484 (
            .O(N__60196),
            .I(N__60173));
    InMux I__14483 (
            .O(N__60195),
            .I(N__60173));
    InMux I__14482 (
            .O(N__60194),
            .I(N__60168));
    InMux I__14481 (
            .O(N__60193),
            .I(N__60168));
    LocalMux I__14480 (
            .O(N__60188),
            .I(N__60159));
    InMux I__14479 (
            .O(N__60187),
            .I(N__60152));
    InMux I__14478 (
            .O(N__60186),
            .I(N__60152));
    LocalMux I__14477 (
            .O(N__60181),
            .I(N__60145));
    Span4Mux_v I__14476 (
            .O(N__60178),
            .I(N__60138));
    LocalMux I__14475 (
            .O(N__60173),
            .I(N__60138));
    LocalMux I__14474 (
            .O(N__60168),
            .I(N__60138));
    InMux I__14473 (
            .O(N__60167),
            .I(N__60133));
    InMux I__14472 (
            .O(N__60166),
            .I(N__60133));
    InMux I__14471 (
            .O(N__60165),
            .I(N__60128));
    InMux I__14470 (
            .O(N__60164),
            .I(N__60128));
    InMux I__14469 (
            .O(N__60163),
            .I(N__60122));
    InMux I__14468 (
            .O(N__60162),
            .I(N__60122));
    Span4Mux_v I__14467 (
            .O(N__60159),
            .I(N__60119));
    InMux I__14466 (
            .O(N__60158),
            .I(N__60114));
    InMux I__14465 (
            .O(N__60157),
            .I(N__60114));
    LocalMux I__14464 (
            .O(N__60152),
            .I(N__60111));
    InMux I__14463 (
            .O(N__60151),
            .I(N__60106));
    InMux I__14462 (
            .O(N__60150),
            .I(N__60106));
    InMux I__14461 (
            .O(N__60149),
            .I(N__60101));
    InMux I__14460 (
            .O(N__60148),
            .I(N__60101));
    Span4Mux_v I__14459 (
            .O(N__60145),
            .I(N__60098));
    Span4Mux_v I__14458 (
            .O(N__60138),
            .I(N__60093));
    LocalMux I__14457 (
            .O(N__60133),
            .I(N__60093));
    LocalMux I__14456 (
            .O(N__60128),
            .I(N__60090));
    InMux I__14455 (
            .O(N__60127),
            .I(N__60087));
    LocalMux I__14454 (
            .O(N__60122),
            .I(N__60084));
    Span4Mux_h I__14453 (
            .O(N__60119),
            .I(N__60081));
    LocalMux I__14452 (
            .O(N__60114),
            .I(N__60078));
    Span4Mux_h I__14451 (
            .O(N__60111),
            .I(N__60073));
    LocalMux I__14450 (
            .O(N__60106),
            .I(N__60073));
    LocalMux I__14449 (
            .O(N__60101),
            .I(N__60070));
    Span4Mux_v I__14448 (
            .O(N__60098),
            .I(N__60063));
    Span4Mux_h I__14447 (
            .O(N__60093),
            .I(N__60063));
    Span4Mux_v I__14446 (
            .O(N__60090),
            .I(N__60063));
    LocalMux I__14445 (
            .O(N__60087),
            .I(N__60060));
    Span12Mux_v I__14444 (
            .O(N__60084),
            .I(N__60057));
    Span4Mux_h I__14443 (
            .O(N__60081),
            .I(N__60054));
    Span4Mux_v I__14442 (
            .O(N__60078),
            .I(N__60051));
    Span4Mux_v I__14441 (
            .O(N__60073),
            .I(N__60046));
    Span4Mux_h I__14440 (
            .O(N__60070),
            .I(N__60046));
    Span4Mux_h I__14439 (
            .O(N__60063),
            .I(N__60041));
    Span4Mux_h I__14438 (
            .O(N__60060),
            .I(N__60041));
    Odrv12 I__14437 (
            .O(N__60057),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ));
    Odrv4 I__14436 (
            .O(N__60054),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ));
    Odrv4 I__14435 (
            .O(N__60051),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ));
    Odrv4 I__14434 (
            .O(N__60046),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ));
    Odrv4 I__14433 (
            .O(N__60041),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ));
    InMux I__14432 (
            .O(N__60030),
            .I(N__60027));
    LocalMux I__14431 (
            .O(N__60027),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_0 ));
    CEMux I__14430 (
            .O(N__60024),
            .I(N__60019));
    CEMux I__14429 (
            .O(N__60023),
            .I(N__60013));
    CEMux I__14428 (
            .O(N__60022),
            .I(N__60010));
    LocalMux I__14427 (
            .O(N__60019),
            .I(N__60006));
    CEMux I__14426 (
            .O(N__60018),
            .I(N__60001));
    CEMux I__14425 (
            .O(N__60017),
            .I(N__59998));
    CEMux I__14424 (
            .O(N__60016),
            .I(N__59995));
    LocalMux I__14423 (
            .O(N__60013),
            .I(N__59991));
    LocalMux I__14422 (
            .O(N__60010),
            .I(N__59988));
    CEMux I__14421 (
            .O(N__60009),
            .I(N__59985));
    Span4Mux_h I__14420 (
            .O(N__60006),
            .I(N__59981));
    CEMux I__14419 (
            .O(N__60005),
            .I(N__59978));
    CEMux I__14418 (
            .O(N__60004),
            .I(N__59975));
    LocalMux I__14417 (
            .O(N__60001),
            .I(N__59972));
    LocalMux I__14416 (
            .O(N__59998),
            .I(N__59969));
    LocalMux I__14415 (
            .O(N__59995),
            .I(N__59966));
    CEMux I__14414 (
            .O(N__59994),
            .I(N__59963));
    Span4Mux_v I__14413 (
            .O(N__59991),
            .I(N__59958));
    Span4Mux_v I__14412 (
            .O(N__59988),
            .I(N__59958));
    LocalMux I__14411 (
            .O(N__59985),
            .I(N__59955));
    CEMux I__14410 (
            .O(N__59984),
            .I(N__59952));
    Span4Mux_h I__14409 (
            .O(N__59981),
            .I(N__59947));
    LocalMux I__14408 (
            .O(N__59978),
            .I(N__59947));
    LocalMux I__14407 (
            .O(N__59975),
            .I(N__59944));
    Span4Mux_h I__14406 (
            .O(N__59972),
            .I(N__59941));
    Span4Mux_v I__14405 (
            .O(N__59969),
            .I(N__59935));
    Span4Mux_v I__14404 (
            .O(N__59966),
            .I(N__59935));
    LocalMux I__14403 (
            .O(N__59963),
            .I(N__59932));
    Span4Mux_h I__14402 (
            .O(N__59958),
            .I(N__59929));
    Span4Mux_v I__14401 (
            .O(N__59955),
            .I(N__59926));
    LocalMux I__14400 (
            .O(N__59952),
            .I(N__59923));
    Span4Mux_h I__14399 (
            .O(N__59947),
            .I(N__59920));
    Span4Mux_v I__14398 (
            .O(N__59944),
            .I(N__59917));
    Span4Mux_h I__14397 (
            .O(N__59941),
            .I(N__59914));
    CEMux I__14396 (
            .O(N__59940),
            .I(N__59911));
    Sp12to4 I__14395 (
            .O(N__59935),
            .I(N__59906));
    Sp12to4 I__14394 (
            .O(N__59932),
            .I(N__59906));
    Span4Mux_h I__14393 (
            .O(N__59929),
            .I(N__59901));
    Span4Mux_v I__14392 (
            .O(N__59926),
            .I(N__59901));
    Span4Mux_h I__14391 (
            .O(N__59923),
            .I(N__59896));
    Span4Mux_v I__14390 (
            .O(N__59920),
            .I(N__59896));
    Span4Mux_h I__14389 (
            .O(N__59917),
            .I(N__59893));
    Span4Mux_h I__14388 (
            .O(N__59914),
            .I(N__59888));
    LocalMux I__14387 (
            .O(N__59911),
            .I(N__59888));
    Span12Mux_h I__14386 (
            .O(N__59906),
            .I(N__59885));
    Span4Mux_h I__14385 (
            .O(N__59901),
            .I(N__59882));
    Span4Mux_h I__14384 (
            .O(N__59896),
            .I(N__59879));
    Span4Mux_v I__14383 (
            .O(N__59893),
            .I(N__59874));
    Span4Mux_v I__14382 (
            .O(N__59888),
            .I(N__59874));
    Odrv12 I__14381 (
            .O(N__59885),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i ));
    Odrv4 I__14380 (
            .O(N__59882),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i ));
    Odrv4 I__14379 (
            .O(N__59879),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i ));
    Odrv4 I__14378 (
            .O(N__59874),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i ));
    InMux I__14377 (
            .O(N__59865),
            .I(N__59860));
    InMux I__14376 (
            .O(N__59864),
            .I(N__59857));
    InMux I__14375 (
            .O(N__59863),
            .I(N__59854));
    LocalMux I__14374 (
            .O(N__59860),
            .I(N__59845));
    LocalMux I__14373 (
            .O(N__59857),
            .I(N__59845));
    LocalMux I__14372 (
            .O(N__59854),
            .I(N__59841));
    InMux I__14371 (
            .O(N__59853),
            .I(N__59838));
    InMux I__14370 (
            .O(N__59852),
            .I(N__59835));
    InMux I__14369 (
            .O(N__59851),
            .I(N__59831));
    InMux I__14368 (
            .O(N__59850),
            .I(N__59828));
    Span4Mux_v I__14367 (
            .O(N__59845),
            .I(N__59825));
    InMux I__14366 (
            .O(N__59844),
            .I(N__59822));
    Span4Mux_h I__14365 (
            .O(N__59841),
            .I(N__59817));
    LocalMux I__14364 (
            .O(N__59838),
            .I(N__59817));
    LocalMux I__14363 (
            .O(N__59835),
            .I(N__59814));
    InMux I__14362 (
            .O(N__59834),
            .I(N__59811));
    LocalMux I__14361 (
            .O(N__59831),
            .I(N__59808));
    LocalMux I__14360 (
            .O(N__59828),
            .I(N__59805));
    Span4Mux_h I__14359 (
            .O(N__59825),
            .I(N__59802));
    LocalMux I__14358 (
            .O(N__59822),
            .I(N__59797));
    Span4Mux_v I__14357 (
            .O(N__59817),
            .I(N__59797));
    Span4Mux_h I__14356 (
            .O(N__59814),
            .I(N__59794));
    LocalMux I__14355 (
            .O(N__59811),
            .I(N__59791));
    Span4Mux_v I__14354 (
            .O(N__59808),
            .I(N__59788));
    Span4Mux_v I__14353 (
            .O(N__59805),
            .I(N__59783));
    Span4Mux_h I__14352 (
            .O(N__59802),
            .I(N__59783));
    Span4Mux_h I__14351 (
            .O(N__59797),
            .I(N__59780));
    Span4Mux_h I__14350 (
            .O(N__59794),
            .I(N__59775));
    Span4Mux_h I__14349 (
            .O(N__59791),
            .I(N__59775));
    Span4Mux_h I__14348 (
            .O(N__59788),
            .I(N__59772));
    Odrv4 I__14347 (
            .O(N__59783),
            .I(I2C_top_level_inst1_s_data_oreg_18));
    Odrv4 I__14346 (
            .O(N__59780),
            .I(I2C_top_level_inst1_s_data_oreg_18));
    Odrv4 I__14345 (
            .O(N__59775),
            .I(I2C_top_level_inst1_s_data_oreg_18));
    Odrv4 I__14344 (
            .O(N__59772),
            .I(I2C_top_level_inst1_s_data_oreg_18));
    InMux I__14343 (
            .O(N__59763),
            .I(N__59760));
    LocalMux I__14342 (
            .O(N__59760),
            .I(N__59757));
    Odrv12 I__14341 (
            .O(N__59757),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_17 ));
    InMux I__14340 (
            .O(N__59754),
            .I(N__59751));
    LocalMux I__14339 (
            .O(N__59751),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_18 ));
    CascadeMux I__14338 (
            .O(N__59748),
            .I(N__59745));
    InMux I__14337 (
            .O(N__59745),
            .I(N__59742));
    LocalMux I__14336 (
            .O(N__59742),
            .I(N__59739));
    Span4Mux_h I__14335 (
            .O(N__59739),
            .I(N__59736));
    Span4Mux_h I__14334 (
            .O(N__59736),
            .I(N__59733));
    Odrv4 I__14333 (
            .O(N__59733),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_29));
    CascadeMux I__14332 (
            .O(N__59730),
            .I(N__59723));
    CascadeMux I__14331 (
            .O(N__59729),
            .I(N__59720));
    CascadeMux I__14330 (
            .O(N__59728),
            .I(N__59699));
    InMux I__14329 (
            .O(N__59727),
            .I(N__59690));
    InMux I__14328 (
            .O(N__59726),
            .I(N__59690));
    InMux I__14327 (
            .O(N__59723),
            .I(N__59677));
    InMux I__14326 (
            .O(N__59720),
            .I(N__59677));
    InMux I__14325 (
            .O(N__59719),
            .I(N__59677));
    InMux I__14324 (
            .O(N__59718),
            .I(N__59677));
    InMux I__14323 (
            .O(N__59717),
            .I(N__59677));
    InMux I__14322 (
            .O(N__59716),
            .I(N__59677));
    InMux I__14321 (
            .O(N__59715),
            .I(N__59654));
    InMux I__14320 (
            .O(N__59714),
            .I(N__59654));
    InMux I__14319 (
            .O(N__59713),
            .I(N__59654));
    InMux I__14318 (
            .O(N__59712),
            .I(N__59654));
    InMux I__14317 (
            .O(N__59711),
            .I(N__59654));
    InMux I__14316 (
            .O(N__59710),
            .I(N__59654));
    InMux I__14315 (
            .O(N__59709),
            .I(N__59654));
    InMux I__14314 (
            .O(N__59708),
            .I(N__59654));
    InMux I__14313 (
            .O(N__59707),
            .I(N__59625));
    InMux I__14312 (
            .O(N__59706),
            .I(N__59625));
    InMux I__14311 (
            .O(N__59705),
            .I(N__59625));
    InMux I__14310 (
            .O(N__59704),
            .I(N__59608));
    InMux I__14309 (
            .O(N__59703),
            .I(N__59608));
    InMux I__14308 (
            .O(N__59702),
            .I(N__59608));
    InMux I__14307 (
            .O(N__59699),
            .I(N__59608));
    InMux I__14306 (
            .O(N__59698),
            .I(N__59608));
    InMux I__14305 (
            .O(N__59697),
            .I(N__59608));
    InMux I__14304 (
            .O(N__59696),
            .I(N__59608));
    InMux I__14303 (
            .O(N__59695),
            .I(N__59608));
    LocalMux I__14302 (
            .O(N__59690),
            .I(N__59582));
    LocalMux I__14301 (
            .O(N__59677),
            .I(N__59582));
    InMux I__14300 (
            .O(N__59676),
            .I(N__59569));
    InMux I__14299 (
            .O(N__59675),
            .I(N__59569));
    InMux I__14298 (
            .O(N__59674),
            .I(N__59569));
    InMux I__14297 (
            .O(N__59673),
            .I(N__59569));
    InMux I__14296 (
            .O(N__59672),
            .I(N__59569));
    InMux I__14295 (
            .O(N__59671),
            .I(N__59569));
    LocalMux I__14294 (
            .O(N__59654),
            .I(N__59566));
    InMux I__14293 (
            .O(N__59653),
            .I(N__59559));
    InMux I__14292 (
            .O(N__59652),
            .I(N__59559));
    InMux I__14291 (
            .O(N__59651),
            .I(N__59559));
    InMux I__14290 (
            .O(N__59650),
            .I(N__59524));
    InMux I__14289 (
            .O(N__59649),
            .I(N__59524));
    InMux I__14288 (
            .O(N__59648),
            .I(N__59524));
    InMux I__14287 (
            .O(N__59647),
            .I(N__59524));
    InMux I__14286 (
            .O(N__59646),
            .I(N__59524));
    InMux I__14285 (
            .O(N__59645),
            .I(N__59524));
    InMux I__14284 (
            .O(N__59644),
            .I(N__59524));
    InMux I__14283 (
            .O(N__59643),
            .I(N__59524));
    InMux I__14282 (
            .O(N__59642),
            .I(N__59517));
    InMux I__14281 (
            .O(N__59641),
            .I(N__59517));
    InMux I__14280 (
            .O(N__59640),
            .I(N__59517));
    InMux I__14279 (
            .O(N__59639),
            .I(N__59487));
    InMux I__14278 (
            .O(N__59638),
            .I(N__59487));
    InMux I__14277 (
            .O(N__59637),
            .I(N__59487));
    InMux I__14276 (
            .O(N__59636),
            .I(N__59487));
    InMux I__14275 (
            .O(N__59635),
            .I(N__59487));
    InMux I__14274 (
            .O(N__59634),
            .I(N__59487));
    InMux I__14273 (
            .O(N__59633),
            .I(N__59487));
    InMux I__14272 (
            .O(N__59632),
            .I(N__59487));
    LocalMux I__14271 (
            .O(N__59625),
            .I(N__59482));
    LocalMux I__14270 (
            .O(N__59608),
            .I(N__59482));
    InMux I__14269 (
            .O(N__59607),
            .I(N__59465));
    InMux I__14268 (
            .O(N__59606),
            .I(N__59465));
    InMux I__14267 (
            .O(N__59605),
            .I(N__59465));
    InMux I__14266 (
            .O(N__59604),
            .I(N__59465));
    InMux I__14265 (
            .O(N__59603),
            .I(N__59465));
    InMux I__14264 (
            .O(N__59602),
            .I(N__59465));
    InMux I__14263 (
            .O(N__59601),
            .I(N__59465));
    InMux I__14262 (
            .O(N__59600),
            .I(N__59465));
    InMux I__14261 (
            .O(N__59599),
            .I(N__59460));
    InMux I__14260 (
            .O(N__59598),
            .I(N__59460));
    InMux I__14259 (
            .O(N__59597),
            .I(N__59449));
    InMux I__14258 (
            .O(N__59596),
            .I(N__59449));
    InMux I__14257 (
            .O(N__59595),
            .I(N__59449));
    InMux I__14256 (
            .O(N__59594),
            .I(N__59449));
    InMux I__14255 (
            .O(N__59593),
            .I(N__59449));
    InMux I__14254 (
            .O(N__59592),
            .I(N__59399));
    InMux I__14253 (
            .O(N__59591),
            .I(N__59399));
    InMux I__14252 (
            .O(N__59590),
            .I(N__59399));
    InMux I__14251 (
            .O(N__59589),
            .I(N__59399));
    InMux I__14250 (
            .O(N__59588),
            .I(N__59399));
    InMux I__14249 (
            .O(N__59587),
            .I(N__59399));
    Span4Mux_v I__14248 (
            .O(N__59582),
            .I(N__59394));
    LocalMux I__14247 (
            .O(N__59569),
            .I(N__59394));
    Span4Mux_h I__14246 (
            .O(N__59566),
            .I(N__59389));
    LocalMux I__14245 (
            .O(N__59559),
            .I(N__59389));
    InMux I__14244 (
            .O(N__59558),
            .I(N__59374));
    InMux I__14243 (
            .O(N__59557),
            .I(N__59374));
    InMux I__14242 (
            .O(N__59556),
            .I(N__59374));
    InMux I__14241 (
            .O(N__59555),
            .I(N__59371));
    InMux I__14240 (
            .O(N__59554),
            .I(N__59368));
    InMux I__14239 (
            .O(N__59553),
            .I(N__59365));
    InMux I__14238 (
            .O(N__59552),
            .I(N__59348));
    InMux I__14237 (
            .O(N__59551),
            .I(N__59348));
    InMux I__14236 (
            .O(N__59550),
            .I(N__59348));
    InMux I__14235 (
            .O(N__59549),
            .I(N__59348));
    InMux I__14234 (
            .O(N__59548),
            .I(N__59348));
    InMux I__14233 (
            .O(N__59547),
            .I(N__59348));
    InMux I__14232 (
            .O(N__59546),
            .I(N__59348));
    InMux I__14231 (
            .O(N__59545),
            .I(N__59348));
    CascadeMux I__14230 (
            .O(N__59544),
            .I(N__59345));
    CascadeMux I__14229 (
            .O(N__59543),
            .I(N__59342));
    CascadeMux I__14228 (
            .O(N__59542),
            .I(N__59339));
    CascadeMux I__14227 (
            .O(N__59541),
            .I(N__59336));
    LocalMux I__14226 (
            .O(N__59524),
            .I(N__59328));
    LocalMux I__14225 (
            .O(N__59517),
            .I(N__59328));
    InMux I__14224 (
            .O(N__59516),
            .I(N__59311));
    InMux I__14223 (
            .O(N__59515),
            .I(N__59311));
    InMux I__14222 (
            .O(N__59514),
            .I(N__59311));
    InMux I__14221 (
            .O(N__59513),
            .I(N__59311));
    InMux I__14220 (
            .O(N__59512),
            .I(N__59311));
    InMux I__14219 (
            .O(N__59511),
            .I(N__59311));
    InMux I__14218 (
            .O(N__59510),
            .I(N__59311));
    InMux I__14217 (
            .O(N__59509),
            .I(N__59311));
    InMux I__14216 (
            .O(N__59508),
            .I(N__59308));
    InMux I__14215 (
            .O(N__59507),
            .I(N__59299));
    InMux I__14214 (
            .O(N__59506),
            .I(N__59299));
    InMux I__14213 (
            .O(N__59505),
            .I(N__59299));
    InMux I__14212 (
            .O(N__59504),
            .I(N__59299));
    LocalMux I__14211 (
            .O(N__59487),
            .I(N__59294));
    Span4Mux_v I__14210 (
            .O(N__59482),
            .I(N__59294));
    LocalMux I__14209 (
            .O(N__59465),
            .I(N__59287));
    LocalMux I__14208 (
            .O(N__59460),
            .I(N__59287));
    LocalMux I__14207 (
            .O(N__59449),
            .I(N__59287));
    CascadeMux I__14206 (
            .O(N__59448),
            .I(N__59284));
    CascadeMux I__14205 (
            .O(N__59447),
            .I(N__59281));
    CascadeMux I__14204 (
            .O(N__59446),
            .I(N__59278));
    CascadeMux I__14203 (
            .O(N__59445),
            .I(N__59272));
    InMux I__14202 (
            .O(N__59444),
            .I(N__59269));
    InMux I__14201 (
            .O(N__59443),
            .I(N__59262));
    InMux I__14200 (
            .O(N__59442),
            .I(N__59262));
    InMux I__14199 (
            .O(N__59441),
            .I(N__59262));
    InMux I__14198 (
            .O(N__59440),
            .I(N__59245));
    InMux I__14197 (
            .O(N__59439),
            .I(N__59245));
    InMux I__14196 (
            .O(N__59438),
            .I(N__59245));
    InMux I__14195 (
            .O(N__59437),
            .I(N__59245));
    InMux I__14194 (
            .O(N__59436),
            .I(N__59245));
    InMux I__14193 (
            .O(N__59435),
            .I(N__59245));
    InMux I__14192 (
            .O(N__59434),
            .I(N__59245));
    InMux I__14191 (
            .O(N__59433),
            .I(N__59245));
    InMux I__14190 (
            .O(N__59432),
            .I(N__59240));
    InMux I__14189 (
            .O(N__59431),
            .I(N__59240));
    InMux I__14188 (
            .O(N__59430),
            .I(N__59223));
    InMux I__14187 (
            .O(N__59429),
            .I(N__59223));
    InMux I__14186 (
            .O(N__59428),
            .I(N__59223));
    InMux I__14185 (
            .O(N__59427),
            .I(N__59223));
    InMux I__14184 (
            .O(N__59426),
            .I(N__59223));
    InMux I__14183 (
            .O(N__59425),
            .I(N__59223));
    InMux I__14182 (
            .O(N__59424),
            .I(N__59223));
    InMux I__14181 (
            .O(N__59423),
            .I(N__59223));
    InMux I__14180 (
            .O(N__59422),
            .I(N__59216));
    InMux I__14179 (
            .O(N__59421),
            .I(N__59216));
    InMux I__14178 (
            .O(N__59420),
            .I(N__59216));
    InMux I__14177 (
            .O(N__59419),
            .I(N__59199));
    InMux I__14176 (
            .O(N__59418),
            .I(N__59199));
    InMux I__14175 (
            .O(N__59417),
            .I(N__59199));
    InMux I__14174 (
            .O(N__59416),
            .I(N__59199));
    InMux I__14173 (
            .O(N__59415),
            .I(N__59199));
    InMux I__14172 (
            .O(N__59414),
            .I(N__59199));
    InMux I__14171 (
            .O(N__59413),
            .I(N__59199));
    InMux I__14170 (
            .O(N__59412),
            .I(N__59199));
    LocalMux I__14169 (
            .O(N__59399),
            .I(N__59194));
    Span4Mux_h I__14168 (
            .O(N__59394),
            .I(N__59194));
    Span4Mux_v I__14167 (
            .O(N__59389),
            .I(N__59191));
    InMux I__14166 (
            .O(N__59388),
            .I(N__59180));
    InMux I__14165 (
            .O(N__59387),
            .I(N__59171));
    InMux I__14164 (
            .O(N__59386),
            .I(N__59171));
    InMux I__14163 (
            .O(N__59385),
            .I(N__59171));
    InMux I__14162 (
            .O(N__59384),
            .I(N__59171));
    InMux I__14161 (
            .O(N__59383),
            .I(N__59166));
    InMux I__14160 (
            .O(N__59382),
            .I(N__59166));
    InMux I__14159 (
            .O(N__59381),
            .I(N__59157));
    LocalMux I__14158 (
            .O(N__59374),
            .I(N__59150));
    LocalMux I__14157 (
            .O(N__59371),
            .I(N__59150));
    LocalMux I__14156 (
            .O(N__59368),
            .I(N__59150));
    LocalMux I__14155 (
            .O(N__59365),
            .I(N__59134));
    LocalMux I__14154 (
            .O(N__59348),
            .I(N__59134));
    InMux I__14153 (
            .O(N__59345),
            .I(N__59119));
    InMux I__14152 (
            .O(N__59342),
            .I(N__59119));
    InMux I__14151 (
            .O(N__59339),
            .I(N__59119));
    InMux I__14150 (
            .O(N__59336),
            .I(N__59119));
    InMux I__14149 (
            .O(N__59335),
            .I(N__59119));
    InMux I__14148 (
            .O(N__59334),
            .I(N__59119));
    InMux I__14147 (
            .O(N__59333),
            .I(N__59119));
    Span4Mux_v I__14146 (
            .O(N__59328),
            .I(N__59106));
    LocalMux I__14145 (
            .O(N__59311),
            .I(N__59106));
    LocalMux I__14144 (
            .O(N__59308),
            .I(N__59106));
    LocalMux I__14143 (
            .O(N__59299),
            .I(N__59106));
    Span4Mux_h I__14142 (
            .O(N__59294),
            .I(N__59106));
    Span4Mux_v I__14141 (
            .O(N__59287),
            .I(N__59106));
    InMux I__14140 (
            .O(N__59284),
            .I(N__59093));
    InMux I__14139 (
            .O(N__59281),
            .I(N__59093));
    InMux I__14138 (
            .O(N__59278),
            .I(N__59093));
    InMux I__14137 (
            .O(N__59277),
            .I(N__59093));
    InMux I__14136 (
            .O(N__59276),
            .I(N__59093));
    InMux I__14135 (
            .O(N__59275),
            .I(N__59093));
    InMux I__14134 (
            .O(N__59272),
            .I(N__59090));
    LocalMux I__14133 (
            .O(N__59269),
            .I(N__59085));
    LocalMux I__14132 (
            .O(N__59262),
            .I(N__59085));
    LocalMux I__14131 (
            .O(N__59245),
            .I(N__59082));
    LocalMux I__14130 (
            .O(N__59240),
            .I(N__59071));
    LocalMux I__14129 (
            .O(N__59223),
            .I(N__59071));
    LocalMux I__14128 (
            .O(N__59216),
            .I(N__59071));
    LocalMux I__14127 (
            .O(N__59199),
            .I(N__59071));
    Span4Mux_v I__14126 (
            .O(N__59194),
            .I(N__59071));
    Span4Mux_v I__14125 (
            .O(N__59191),
            .I(N__59068));
    InMux I__14124 (
            .O(N__59190),
            .I(N__59051));
    InMux I__14123 (
            .O(N__59189),
            .I(N__59051));
    InMux I__14122 (
            .O(N__59188),
            .I(N__59051));
    InMux I__14121 (
            .O(N__59187),
            .I(N__59051));
    InMux I__14120 (
            .O(N__59186),
            .I(N__59051));
    InMux I__14119 (
            .O(N__59185),
            .I(N__59051));
    InMux I__14118 (
            .O(N__59184),
            .I(N__59051));
    InMux I__14117 (
            .O(N__59183),
            .I(N__59051));
    LocalMux I__14116 (
            .O(N__59180),
            .I(N__59046));
    LocalMux I__14115 (
            .O(N__59171),
            .I(N__59046));
    LocalMux I__14114 (
            .O(N__59166),
            .I(N__59043));
    InMux I__14113 (
            .O(N__59165),
            .I(N__59038));
    InMux I__14112 (
            .O(N__59164),
            .I(N__59038));
    CascadeMux I__14111 (
            .O(N__59163),
            .I(N__59035));
    CascadeMux I__14110 (
            .O(N__59162),
            .I(N__59032));
    CascadeMux I__14109 (
            .O(N__59161),
            .I(N__59029));
    CascadeMux I__14108 (
            .O(N__59160),
            .I(N__59026));
    LocalMux I__14107 (
            .O(N__59157),
            .I(N__59020));
    Span4Mux_v I__14106 (
            .O(N__59150),
            .I(N__59017));
    InMux I__14105 (
            .O(N__59149),
            .I(N__58993));
    InMux I__14104 (
            .O(N__59148),
            .I(N__58993));
    InMux I__14103 (
            .O(N__59147),
            .I(N__58993));
    InMux I__14102 (
            .O(N__59146),
            .I(N__58993));
    InMux I__14101 (
            .O(N__59145),
            .I(N__58993));
    InMux I__14100 (
            .O(N__59144),
            .I(N__58993));
    InMux I__14099 (
            .O(N__59143),
            .I(N__58993));
    InMux I__14098 (
            .O(N__59142),
            .I(N__58993));
    InMux I__14097 (
            .O(N__59141),
            .I(N__58988));
    InMux I__14096 (
            .O(N__59140),
            .I(N__58988));
    InMux I__14095 (
            .O(N__59139),
            .I(N__58985));
    Span4Mux_v I__14094 (
            .O(N__59134),
            .I(N__58978));
    LocalMux I__14093 (
            .O(N__59119),
            .I(N__58978));
    Span4Mux_h I__14092 (
            .O(N__59106),
            .I(N__58978));
    LocalMux I__14091 (
            .O(N__59093),
            .I(N__58971));
    LocalMux I__14090 (
            .O(N__59090),
            .I(N__58971));
    Span4Mux_v I__14089 (
            .O(N__59085),
            .I(N__58971));
    Span4Mux_v I__14088 (
            .O(N__59082),
            .I(N__58964));
    Span4Mux_v I__14087 (
            .O(N__59071),
            .I(N__58964));
    Span4Mux_h I__14086 (
            .O(N__59068),
            .I(N__58964));
    LocalMux I__14085 (
            .O(N__59051),
            .I(N__58955));
    Span4Mux_v I__14084 (
            .O(N__59046),
            .I(N__58955));
    Span4Mux_h I__14083 (
            .O(N__59043),
            .I(N__58955));
    LocalMux I__14082 (
            .O(N__59038),
            .I(N__58955));
    InMux I__14081 (
            .O(N__59035),
            .I(N__58940));
    InMux I__14080 (
            .O(N__59032),
            .I(N__58940));
    InMux I__14079 (
            .O(N__59029),
            .I(N__58940));
    InMux I__14078 (
            .O(N__59026),
            .I(N__58940));
    InMux I__14077 (
            .O(N__59025),
            .I(N__58940));
    InMux I__14076 (
            .O(N__59024),
            .I(N__58940));
    InMux I__14075 (
            .O(N__59023),
            .I(N__58940));
    Span4Mux_v I__14074 (
            .O(N__59020),
            .I(N__58935));
    Span4Mux_v I__14073 (
            .O(N__59017),
            .I(N__58935));
    InMux I__14072 (
            .O(N__59016),
            .I(N__58926));
    InMux I__14071 (
            .O(N__59015),
            .I(N__58926));
    InMux I__14070 (
            .O(N__59014),
            .I(N__58926));
    InMux I__14069 (
            .O(N__59013),
            .I(N__58926));
    InMux I__14068 (
            .O(N__59012),
            .I(N__58919));
    InMux I__14067 (
            .O(N__59011),
            .I(N__58919));
    InMux I__14066 (
            .O(N__59010),
            .I(N__58919));
    LocalMux I__14065 (
            .O(N__58993),
            .I(N__58916));
    LocalMux I__14064 (
            .O(N__58988),
            .I(N__58909));
    LocalMux I__14063 (
            .O(N__58985),
            .I(N__58909));
    Span4Mux_h I__14062 (
            .O(N__58978),
            .I(N__58909));
    Span4Mux_v I__14061 (
            .O(N__58971),
            .I(N__58902));
    Span4Mux_h I__14060 (
            .O(N__58964),
            .I(N__58902));
    Span4Mux_v I__14059 (
            .O(N__58955),
            .I(N__58902));
    LocalMux I__14058 (
            .O(N__58940),
            .I(N__58897));
    Span4Mux_h I__14057 (
            .O(N__58935),
            .I(N__58897));
    LocalMux I__14056 (
            .O(N__58926),
            .I(N_1592_0));
    LocalMux I__14055 (
            .O(N__58919),
            .I(N_1592_0));
    Odrv12 I__14054 (
            .O(N__58916),
            .I(N_1592_0));
    Odrv4 I__14053 (
            .O(N__58909),
            .I(N_1592_0));
    Odrv4 I__14052 (
            .O(N__58902),
            .I(N_1592_0));
    Odrv4 I__14051 (
            .O(N__58897),
            .I(N_1592_0));
    CEMux I__14050 (
            .O(N__58884),
            .I(N__58881));
    LocalMux I__14049 (
            .O(N__58881),
            .I(N__58876));
    CEMux I__14048 (
            .O(N__58880),
            .I(N__58873));
    CEMux I__14047 (
            .O(N__58879),
            .I(N__58870));
    Span4Mux_h I__14046 (
            .O(N__58876),
            .I(N__58862));
    LocalMux I__14045 (
            .O(N__58873),
            .I(N__58862));
    LocalMux I__14044 (
            .O(N__58870),
            .I(N__58859));
    CEMux I__14043 (
            .O(N__58869),
            .I(N__58856));
    CEMux I__14042 (
            .O(N__58868),
            .I(N__58853));
    CEMux I__14041 (
            .O(N__58867),
            .I(N__58850));
    Span4Mux_h I__14040 (
            .O(N__58862),
            .I(N__58843));
    Span4Mux_h I__14039 (
            .O(N__58859),
            .I(N__58843));
    LocalMux I__14038 (
            .O(N__58856),
            .I(N__58843));
    LocalMux I__14037 (
            .O(N__58853),
            .I(N__58840));
    LocalMux I__14036 (
            .O(N__58850),
            .I(N__58837));
    Span4Mux_v I__14035 (
            .O(N__58843),
            .I(N__58834));
    Span12Mux_v I__14034 (
            .O(N__58840),
            .I(N__58831));
    Span4Mux_v I__14033 (
            .O(N__58837),
            .I(N__58828));
    Span4Mux_h I__14032 (
            .O(N__58834),
            .I(N__58825));
    Odrv12 I__14031 (
            .O(N__58831),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0 ));
    Odrv4 I__14030 (
            .O(N__58828),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0 ));
    Odrv4 I__14029 (
            .O(N__58825),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0 ));
    InMux I__14028 (
            .O(N__58818),
            .I(N__58815));
    LocalMux I__14027 (
            .O(N__58815),
            .I(N__58812));
    Span4Mux_v I__14026 (
            .O(N__58812),
            .I(N__58809));
    Span4Mux_h I__14025 (
            .O(N__58809),
            .I(N__58806));
    Sp12to4 I__14024 (
            .O(N__58806),
            .I(N__58803));
    Span12Mux_h I__14023 (
            .O(N__58803),
            .I(N__58800));
    Odrv12 I__14022 (
            .O(N__58800),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_9 ));
    InMux I__14021 (
            .O(N__58797),
            .I(N__58792));
    InMux I__14020 (
            .O(N__58796),
            .I(N__58789));
    InMux I__14019 (
            .O(N__58795),
            .I(N__58784));
    LocalMux I__14018 (
            .O(N__58792),
            .I(N__58780));
    LocalMux I__14017 (
            .O(N__58789),
            .I(N__58776));
    InMux I__14016 (
            .O(N__58788),
            .I(N__58773));
    InMux I__14015 (
            .O(N__58787),
            .I(N__58770));
    LocalMux I__14014 (
            .O(N__58784),
            .I(N__58767));
    InMux I__14013 (
            .O(N__58783),
            .I(N__58763));
    Span4Mux_h I__14012 (
            .O(N__58780),
            .I(N__58760));
    InMux I__14011 (
            .O(N__58779),
            .I(N__58757));
    Span4Mux_h I__14010 (
            .O(N__58776),
            .I(N__58750));
    LocalMux I__14009 (
            .O(N__58773),
            .I(N__58750));
    LocalMux I__14008 (
            .O(N__58770),
            .I(N__58750));
    Span4Mux_v I__14007 (
            .O(N__58767),
            .I(N__58746));
    CascadeMux I__14006 (
            .O(N__58766),
            .I(N__58743));
    LocalMux I__14005 (
            .O(N__58763),
            .I(N__58738));
    Span4Mux_h I__14004 (
            .O(N__58760),
            .I(N__58738));
    LocalMux I__14003 (
            .O(N__58757),
            .I(N__58733));
    Sp12to4 I__14002 (
            .O(N__58750),
            .I(N__58733));
    InMux I__14001 (
            .O(N__58749),
            .I(N__58730));
    Sp12to4 I__14000 (
            .O(N__58746),
            .I(N__58727));
    InMux I__13999 (
            .O(N__58743),
            .I(N__58724));
    Span4Mux_v I__13998 (
            .O(N__58738),
            .I(N__58721));
    Span12Mux_v I__13997 (
            .O(N__58733),
            .I(N__58716));
    LocalMux I__13996 (
            .O(N__58730),
            .I(N__58716));
    Odrv12 I__13995 (
            .O(N__58727),
            .I(I2C_top_level_inst1_s_data_oreg_10));
    LocalMux I__13994 (
            .O(N__58724),
            .I(I2C_top_level_inst1_s_data_oreg_10));
    Odrv4 I__13993 (
            .O(N__58721),
            .I(I2C_top_level_inst1_s_data_oreg_10));
    Odrv12 I__13992 (
            .O(N__58716),
            .I(I2C_top_level_inst1_s_data_oreg_10));
    InMux I__13991 (
            .O(N__58707),
            .I(N__58704));
    LocalMux I__13990 (
            .O(N__58704),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_10 ));
    InMux I__13989 (
            .O(N__58701),
            .I(N__58697));
    InMux I__13988 (
            .O(N__58700),
            .I(N__58693));
    LocalMux I__13987 (
            .O(N__58697),
            .I(N__58688));
    InMux I__13986 (
            .O(N__58696),
            .I(N__58685));
    LocalMux I__13985 (
            .O(N__58693),
            .I(N__58681));
    InMux I__13984 (
            .O(N__58692),
            .I(N__58678));
    InMux I__13983 (
            .O(N__58691),
            .I(N__58675));
    Span4Mux_v I__13982 (
            .O(N__58688),
            .I(N__58670));
    LocalMux I__13981 (
            .O(N__58685),
            .I(N__58670));
    InMux I__13980 (
            .O(N__58684),
            .I(N__58667));
    Span4Mux_h I__13979 (
            .O(N__58681),
            .I(N__58661));
    LocalMux I__13978 (
            .O(N__58678),
            .I(N__58661));
    LocalMux I__13977 (
            .O(N__58675),
            .I(N__58657));
    Span4Mux_h I__13976 (
            .O(N__58670),
            .I(N__58652));
    LocalMux I__13975 (
            .O(N__58667),
            .I(N__58652));
    InMux I__13974 (
            .O(N__58666),
            .I(N__58649));
    Span4Mux_v I__13973 (
            .O(N__58661),
            .I(N__58646));
    InMux I__13972 (
            .O(N__58660),
            .I(N__58643));
    Span4Mux_v I__13971 (
            .O(N__58657),
            .I(N__58638));
    Span4Mux_v I__13970 (
            .O(N__58652),
            .I(N__58638));
    LocalMux I__13969 (
            .O(N__58649),
            .I(N__58635));
    Span4Mux_h I__13968 (
            .O(N__58646),
            .I(N__58629));
    LocalMux I__13967 (
            .O(N__58643),
            .I(N__58629));
    Sp12to4 I__13966 (
            .O(N__58638),
            .I(N__58626));
    Span4Mux_v I__13965 (
            .O(N__58635),
            .I(N__58623));
    CascadeMux I__13964 (
            .O(N__58634),
            .I(N__58620));
    Span4Mux_v I__13963 (
            .O(N__58629),
            .I(N__58617));
    Span12Mux_h I__13962 (
            .O(N__58626),
            .I(N__58612));
    Sp12to4 I__13961 (
            .O(N__58623),
            .I(N__58612));
    InMux I__13960 (
            .O(N__58620),
            .I(N__58609));
    Odrv4 I__13959 (
            .O(N__58617),
            .I(I2C_top_level_inst1_s_data_oreg_11));
    Odrv12 I__13958 (
            .O(N__58612),
            .I(I2C_top_level_inst1_s_data_oreg_11));
    LocalMux I__13957 (
            .O(N__58609),
            .I(I2C_top_level_inst1_s_data_oreg_11));
    InMux I__13956 (
            .O(N__58602),
            .I(N__58599));
    LocalMux I__13955 (
            .O(N__58599),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_11 ));
    InMux I__13954 (
            .O(N__58596),
            .I(N__58586));
    InMux I__13953 (
            .O(N__58595),
            .I(N__58583));
    InMux I__13952 (
            .O(N__58594),
            .I(N__58580));
    CascadeMux I__13951 (
            .O(N__58593),
            .I(N__58577));
    InMux I__13950 (
            .O(N__58592),
            .I(N__58574));
    InMux I__13949 (
            .O(N__58591),
            .I(N__58571));
    InMux I__13948 (
            .O(N__58590),
            .I(N__58568));
    InMux I__13947 (
            .O(N__58589),
            .I(N__58565));
    LocalMux I__13946 (
            .O(N__58586),
            .I(N__58562));
    LocalMux I__13945 (
            .O(N__58583),
            .I(N__58556));
    LocalMux I__13944 (
            .O(N__58580),
            .I(N__58556));
    InMux I__13943 (
            .O(N__58577),
            .I(N__58553));
    LocalMux I__13942 (
            .O(N__58574),
            .I(N__58550));
    LocalMux I__13941 (
            .O(N__58571),
            .I(N__58545));
    LocalMux I__13940 (
            .O(N__58568),
            .I(N__58545));
    LocalMux I__13939 (
            .O(N__58565),
            .I(N__58540));
    Span4Mux_h I__13938 (
            .O(N__58562),
            .I(N__58540));
    InMux I__13937 (
            .O(N__58561),
            .I(N__58537));
    Span4Mux_v I__13936 (
            .O(N__58556),
            .I(N__58534));
    LocalMux I__13935 (
            .O(N__58553),
            .I(N__58531));
    Span4Mux_h I__13934 (
            .O(N__58550),
            .I(N__58524));
    Span4Mux_v I__13933 (
            .O(N__58545),
            .I(N__58524));
    Span4Mux_v I__13932 (
            .O(N__58540),
            .I(N__58524));
    LocalMux I__13931 (
            .O(N__58537),
            .I(N__58521));
    Span4Mux_h I__13930 (
            .O(N__58534),
            .I(N__58518));
    Span4Mux_v I__13929 (
            .O(N__58531),
            .I(N__58515));
    Span4Mux_h I__13928 (
            .O(N__58524),
            .I(N__58512));
    Span12Mux_s8_v I__13927 (
            .O(N__58521),
            .I(N__58509));
    Odrv4 I__13926 (
            .O(N__58518),
            .I(I2C_top_level_inst1_s_data_oreg_12));
    Odrv4 I__13925 (
            .O(N__58515),
            .I(I2C_top_level_inst1_s_data_oreg_12));
    Odrv4 I__13924 (
            .O(N__58512),
            .I(I2C_top_level_inst1_s_data_oreg_12));
    Odrv12 I__13923 (
            .O(N__58509),
            .I(I2C_top_level_inst1_s_data_oreg_12));
    InMux I__13922 (
            .O(N__58500),
            .I(N__58493));
    InMux I__13921 (
            .O(N__58499),
            .I(N__58490));
    InMux I__13920 (
            .O(N__58498),
            .I(N__58486));
    InMux I__13919 (
            .O(N__58497),
            .I(N__58483));
    InMux I__13918 (
            .O(N__58496),
            .I(N__58480));
    LocalMux I__13917 (
            .O(N__58493),
            .I(N__58477));
    LocalMux I__13916 (
            .O(N__58490),
            .I(N__58474));
    InMux I__13915 (
            .O(N__58489),
            .I(N__58470));
    LocalMux I__13914 (
            .O(N__58486),
            .I(N__58465));
    LocalMux I__13913 (
            .O(N__58483),
            .I(N__58465));
    LocalMux I__13912 (
            .O(N__58480),
            .I(N__58462));
    Span4Mux_v I__13911 (
            .O(N__58477),
            .I(N__58459));
    Span4Mux_v I__13910 (
            .O(N__58474),
            .I(N__58456));
    InMux I__13909 (
            .O(N__58473),
            .I(N__58452));
    LocalMux I__13908 (
            .O(N__58470),
            .I(N__58449));
    Span4Mux_h I__13907 (
            .O(N__58465),
            .I(N__58444));
    Span4Mux_v I__13906 (
            .O(N__58462),
            .I(N__58444));
    Span4Mux_h I__13905 (
            .O(N__58459),
            .I(N__58441));
    Span4Mux_h I__13904 (
            .O(N__58456),
            .I(N__58437));
    InMux I__13903 (
            .O(N__58455),
            .I(N__58434));
    LocalMux I__13902 (
            .O(N__58452),
            .I(N__58431));
    Span4Mux_v I__13901 (
            .O(N__58449),
            .I(N__58428));
    Span4Mux_v I__13900 (
            .O(N__58444),
            .I(N__58425));
    Span4Mux_h I__13899 (
            .O(N__58441),
            .I(N__58422));
    CascadeMux I__13898 (
            .O(N__58440),
            .I(N__58419));
    Span4Mux_v I__13897 (
            .O(N__58437),
            .I(N__58416));
    LocalMux I__13896 (
            .O(N__58434),
            .I(N__58413));
    Span12Mux_v I__13895 (
            .O(N__58431),
            .I(N__58406));
    Sp12to4 I__13894 (
            .O(N__58428),
            .I(N__58406));
    Sp12to4 I__13893 (
            .O(N__58425),
            .I(N__58406));
    Span4Mux_v I__13892 (
            .O(N__58422),
            .I(N__58403));
    InMux I__13891 (
            .O(N__58419),
            .I(N__58400));
    Span4Mux_h I__13890 (
            .O(N__58416),
            .I(N__58395));
    Span4Mux_h I__13889 (
            .O(N__58413),
            .I(N__58395));
    Odrv12 I__13888 (
            .O(N__58406),
            .I(I2C_top_level_inst1_s_data_oreg_14));
    Odrv4 I__13887 (
            .O(N__58403),
            .I(I2C_top_level_inst1_s_data_oreg_14));
    LocalMux I__13886 (
            .O(N__58400),
            .I(I2C_top_level_inst1_s_data_oreg_14));
    Odrv4 I__13885 (
            .O(N__58395),
            .I(I2C_top_level_inst1_s_data_oreg_14));
    InMux I__13884 (
            .O(N__58386),
            .I(N__58383));
    LocalMux I__13883 (
            .O(N__58383),
            .I(N__58380));
    Odrv4 I__13882 (
            .O(N__58380),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_14 ));
    InMux I__13881 (
            .O(N__58377),
            .I(N__58373));
    InMux I__13880 (
            .O(N__58376),
            .I(N__58370));
    LocalMux I__13879 (
            .O(N__58373),
            .I(N__58365));
    LocalMux I__13878 (
            .O(N__58370),
            .I(N__58365));
    Span4Mux_h I__13877 (
            .O(N__58365),
            .I(N__58361));
    InMux I__13876 (
            .O(N__58364),
            .I(N__58358));
    Span4Mux_v I__13875 (
            .O(N__58361),
            .I(N__58352));
    LocalMux I__13874 (
            .O(N__58358),
            .I(N__58352));
    CascadeMux I__13873 (
            .O(N__58357),
            .I(N__58345));
    Span4Mux_v I__13872 (
            .O(N__58352),
            .I(N__58342));
    InMux I__13871 (
            .O(N__58351),
            .I(N__58339));
    InMux I__13870 (
            .O(N__58350),
            .I(N__58336));
    InMux I__13869 (
            .O(N__58349),
            .I(N__58333));
    InMux I__13868 (
            .O(N__58348),
            .I(N__58329));
    InMux I__13867 (
            .O(N__58345),
            .I(N__58326));
    Span4Mux_v I__13866 (
            .O(N__58342),
            .I(N__58323));
    LocalMux I__13865 (
            .O(N__58339),
            .I(N__58316));
    LocalMux I__13864 (
            .O(N__58336),
            .I(N__58316));
    LocalMux I__13863 (
            .O(N__58333),
            .I(N__58316));
    InMux I__13862 (
            .O(N__58332),
            .I(N__58313));
    LocalMux I__13861 (
            .O(N__58329),
            .I(N__58310));
    LocalMux I__13860 (
            .O(N__58326),
            .I(N__58307));
    Span4Mux_h I__13859 (
            .O(N__58323),
            .I(N__58302));
    Span4Mux_v I__13858 (
            .O(N__58316),
            .I(N__58302));
    LocalMux I__13857 (
            .O(N__58313),
            .I(N__58299));
    Span4Mux_v I__13856 (
            .O(N__58310),
            .I(N__58296));
    Span4Mux_v I__13855 (
            .O(N__58307),
            .I(N__58293));
    Span4Mux_v I__13854 (
            .O(N__58302),
            .I(N__58290));
    Span4Mux_h I__13853 (
            .O(N__58299),
            .I(N__58287));
    Sp12to4 I__13852 (
            .O(N__58296),
            .I(N__58284));
    Span4Mux_v I__13851 (
            .O(N__58293),
            .I(N__58281));
    Span4Mux_h I__13850 (
            .O(N__58290),
            .I(N__58276));
    Span4Mux_h I__13849 (
            .O(N__58287),
            .I(N__58276));
    Odrv12 I__13848 (
            .O(N__58284),
            .I(I2C_top_level_inst1_s_data_oreg_13));
    Odrv4 I__13847 (
            .O(N__58281),
            .I(I2C_top_level_inst1_s_data_oreg_13));
    Odrv4 I__13846 (
            .O(N__58276),
            .I(I2C_top_level_inst1_s_data_oreg_13));
    InMux I__13845 (
            .O(N__58269),
            .I(N__58266));
    LocalMux I__13844 (
            .O(N__58266),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_12 ));
    InMux I__13843 (
            .O(N__58263),
            .I(N__58260));
    LocalMux I__13842 (
            .O(N__58260),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_13 ));
    CascadeMux I__13841 (
            .O(N__58257),
            .I(N__58253));
    InMux I__13840 (
            .O(N__58256),
            .I(N__58250));
    InMux I__13839 (
            .O(N__58253),
            .I(N__58247));
    LocalMux I__13838 (
            .O(N__58250),
            .I(N__58243));
    LocalMux I__13837 (
            .O(N__58247),
            .I(N__58240));
    InMux I__13836 (
            .O(N__58246),
            .I(N__58237));
    Span4Mux_v I__13835 (
            .O(N__58243),
            .I(N__58232));
    Span4Mux_v I__13834 (
            .O(N__58240),
            .I(N__58232));
    LocalMux I__13833 (
            .O(N__58237),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_0));
    Odrv4 I__13832 (
            .O(N__58232),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_0));
    InMux I__13831 (
            .O(N__58227),
            .I(N__58224));
    LocalMux I__13830 (
            .O(N__58224),
            .I(N__58220));
    InMux I__13829 (
            .O(N__58223),
            .I(N__58217));
    Span4Mux_v I__13828 (
            .O(N__58220),
            .I(N__58212));
    LocalMux I__13827 (
            .O(N__58217),
            .I(N__58212));
    Span4Mux_v I__13826 (
            .O(N__58212),
            .I(N__58208));
    InMux I__13825 (
            .O(N__58211),
            .I(N__58205));
    Odrv4 I__13824 (
            .O(N__58208),
            .I(cemf_module_64ch_ctrl_inst1_data_config_0));
    LocalMux I__13823 (
            .O(N__58205),
            .I(cemf_module_64ch_ctrl_inst1_data_config_0));
    InMux I__13822 (
            .O(N__58200),
            .I(N__58191));
    InMux I__13821 (
            .O(N__58199),
            .I(N__58191));
    CascadeMux I__13820 (
            .O(N__58198),
            .I(N__58187));
    InMux I__13819 (
            .O(N__58197),
            .I(N__58174));
    InMux I__13818 (
            .O(N__58196),
            .I(N__58174));
    LocalMux I__13817 (
            .O(N__58191),
            .I(N__58171));
    InMux I__13816 (
            .O(N__58190),
            .I(N__58166));
    InMux I__13815 (
            .O(N__58187),
            .I(N__58166));
    InMux I__13814 (
            .O(N__58186),
            .I(N__58160));
    InMux I__13813 (
            .O(N__58185),
            .I(N__58160));
    InMux I__13812 (
            .O(N__58184),
            .I(N__58153));
    InMux I__13811 (
            .O(N__58183),
            .I(N__58148));
    InMux I__13810 (
            .O(N__58182),
            .I(N__58148));
    InMux I__13809 (
            .O(N__58181),
            .I(N__58143));
    InMux I__13808 (
            .O(N__58180),
            .I(N__58143));
    InMux I__13807 (
            .O(N__58179),
            .I(N__58140));
    LocalMux I__13806 (
            .O(N__58174),
            .I(N__58135));
    Span4Mux_v I__13805 (
            .O(N__58171),
            .I(N__58135));
    LocalMux I__13804 (
            .O(N__58166),
            .I(N__58132));
    InMux I__13803 (
            .O(N__58165),
            .I(N__58129));
    LocalMux I__13802 (
            .O(N__58160),
            .I(N__58126));
    InMux I__13801 (
            .O(N__58159),
            .I(N__58121));
    InMux I__13800 (
            .O(N__58158),
            .I(N__58121));
    InMux I__13799 (
            .O(N__58157),
            .I(N__58117));
    InMux I__13798 (
            .O(N__58156),
            .I(N__58114));
    LocalMux I__13797 (
            .O(N__58153),
            .I(N__58105));
    LocalMux I__13796 (
            .O(N__58148),
            .I(N__58105));
    LocalMux I__13795 (
            .O(N__58143),
            .I(N__58102));
    LocalMux I__13794 (
            .O(N__58140),
            .I(N__58099));
    Span4Mux_h I__13793 (
            .O(N__58135),
            .I(N__58094));
    Span4Mux_h I__13792 (
            .O(N__58132),
            .I(N__58094));
    LocalMux I__13791 (
            .O(N__58129),
            .I(N__58089));
    Span4Mux_h I__13790 (
            .O(N__58126),
            .I(N__58089));
    LocalMux I__13789 (
            .O(N__58121),
            .I(N__58086));
    InMux I__13788 (
            .O(N__58120),
            .I(N__58083));
    LocalMux I__13787 (
            .O(N__58117),
            .I(N__58078));
    LocalMux I__13786 (
            .O(N__58114),
            .I(N__58078));
    InMux I__13785 (
            .O(N__58113),
            .I(N__58073));
    InMux I__13784 (
            .O(N__58112),
            .I(N__58073));
    InMux I__13783 (
            .O(N__58111),
            .I(N__58068));
    InMux I__13782 (
            .O(N__58110),
            .I(N__58068));
    Span4Mux_v I__13781 (
            .O(N__58105),
            .I(N__58065));
    Span4Mux_v I__13780 (
            .O(N__58102),
            .I(N__58060));
    Span4Mux_v I__13779 (
            .O(N__58099),
            .I(N__58060));
    Span4Mux_v I__13778 (
            .O(N__58094),
            .I(N__58057));
    Span4Mux_v I__13777 (
            .O(N__58089),
            .I(N__58050));
    Span4Mux_v I__13776 (
            .O(N__58086),
            .I(N__58050));
    LocalMux I__13775 (
            .O(N__58083),
            .I(N__58050));
    Span4Mux_v I__13774 (
            .O(N__58078),
            .I(N__58045));
    LocalMux I__13773 (
            .O(N__58073),
            .I(N__58045));
    LocalMux I__13772 (
            .O(N__58068),
            .I(N__58038));
    Sp12to4 I__13771 (
            .O(N__58065),
            .I(N__58038));
    Sp12to4 I__13770 (
            .O(N__58060),
            .I(N__58038));
    Sp12to4 I__13769 (
            .O(N__58057),
            .I(N__58035));
    Span4Mux_h I__13768 (
            .O(N__58050),
            .I(N__58032));
    Sp12to4 I__13767 (
            .O(N__58045),
            .I(N__58027));
    Span12Mux_h I__13766 (
            .O(N__58038),
            .I(N__58027));
    Span12Mux_v I__13765 (
            .O(N__58035),
            .I(N__58024));
    Odrv4 I__13764 (
            .O(N__58032),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0 ));
    Odrv12 I__13763 (
            .O(N__58027),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0 ));
    Odrv12 I__13762 (
            .O(N__58024),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0 ));
    InMux I__13761 (
            .O(N__58017),
            .I(N__58008));
    InMux I__13760 (
            .O(N__58016),
            .I(N__58008));
    InMux I__13759 (
            .O(N__58015),
            .I(N__58001));
    InMux I__13758 (
            .O(N__58014),
            .I(N__57996));
    InMux I__13757 (
            .O(N__58013),
            .I(N__57996));
    LocalMux I__13756 (
            .O(N__58008),
            .I(N__57993));
    InMux I__13755 (
            .O(N__58007),
            .I(N__57982));
    InMux I__13754 (
            .O(N__58006),
            .I(N__57982));
    InMux I__13753 (
            .O(N__58005),
            .I(N__57973));
    InMux I__13752 (
            .O(N__58004),
            .I(N__57973));
    LocalMux I__13751 (
            .O(N__58001),
            .I(N__57970));
    LocalMux I__13750 (
            .O(N__57996),
            .I(N__57967));
    Span4Mux_v I__13749 (
            .O(N__57993),
            .I(N__57964));
    InMux I__13748 (
            .O(N__57992),
            .I(N__57959));
    InMux I__13747 (
            .O(N__57991),
            .I(N__57959));
    InMux I__13746 (
            .O(N__57990),
            .I(N__57954));
    InMux I__13745 (
            .O(N__57989),
            .I(N__57954));
    InMux I__13744 (
            .O(N__57988),
            .I(N__57949));
    InMux I__13743 (
            .O(N__57987),
            .I(N__57949));
    LocalMux I__13742 (
            .O(N__57982),
            .I(N__57946));
    InMux I__13741 (
            .O(N__57981),
            .I(N__57943));
    InMux I__13740 (
            .O(N__57980),
            .I(N__57936));
    InMux I__13739 (
            .O(N__57979),
            .I(N__57936));
    InMux I__13738 (
            .O(N__57978),
            .I(N__57932));
    LocalMux I__13737 (
            .O(N__57973),
            .I(N__57927));
    Span4Mux_v I__13736 (
            .O(N__57970),
            .I(N__57927));
    Span4Mux_v I__13735 (
            .O(N__57967),
            .I(N__57923));
    Span4Mux_h I__13734 (
            .O(N__57964),
            .I(N__57918));
    LocalMux I__13733 (
            .O(N__57959),
            .I(N__57918));
    LocalMux I__13732 (
            .O(N__57954),
            .I(N__57915));
    LocalMux I__13731 (
            .O(N__57949),
            .I(N__57911));
    Span4Mux_h I__13730 (
            .O(N__57946),
            .I(N__57906));
    LocalMux I__13729 (
            .O(N__57943),
            .I(N__57906));
    InMux I__13728 (
            .O(N__57942),
            .I(N__57901));
    InMux I__13727 (
            .O(N__57941),
            .I(N__57901));
    LocalMux I__13726 (
            .O(N__57936),
            .I(N__57898));
    InMux I__13725 (
            .O(N__57935),
            .I(N__57895));
    LocalMux I__13724 (
            .O(N__57932),
            .I(N__57890));
    Span4Mux_h I__13723 (
            .O(N__57927),
            .I(N__57890));
    InMux I__13722 (
            .O(N__57926),
            .I(N__57887));
    Span4Mux_h I__13721 (
            .O(N__57923),
            .I(N__57880));
    Span4Mux_v I__13720 (
            .O(N__57918),
            .I(N__57880));
    Span4Mux_v I__13719 (
            .O(N__57915),
            .I(N__57880));
    InMux I__13718 (
            .O(N__57914),
            .I(N__57877));
    Span4Mux_v I__13717 (
            .O(N__57911),
            .I(N__57872));
    Span4Mux_v I__13716 (
            .O(N__57906),
            .I(N__57872));
    LocalMux I__13715 (
            .O(N__57901),
            .I(N__57869));
    Span4Mux_h I__13714 (
            .O(N__57898),
            .I(N__57866));
    LocalMux I__13713 (
            .O(N__57895),
            .I(N__57861));
    Span4Mux_h I__13712 (
            .O(N__57890),
            .I(N__57861));
    LocalMux I__13711 (
            .O(N__57887),
            .I(N__57852));
    Sp12to4 I__13710 (
            .O(N__57880),
            .I(N__57852));
    LocalMux I__13709 (
            .O(N__57877),
            .I(N__57852));
    Sp12to4 I__13708 (
            .O(N__57872),
            .I(N__57852));
    Span4Mux_v I__13707 (
            .O(N__57869),
            .I(N__57849));
    Span4Mux_h I__13706 (
            .O(N__57866),
            .I(N__57846));
    Sp12to4 I__13705 (
            .O(N__57861),
            .I(N__57841));
    Span12Mux_h I__13704 (
            .O(N__57852),
            .I(N__57841));
    Odrv4 I__13703 (
            .O(N__57849),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273 ));
    Odrv4 I__13702 (
            .O(N__57846),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273 ));
    Odrv12 I__13701 (
            .O(N__57841),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273 ));
    InMux I__13700 (
            .O(N__57834),
            .I(N__57830));
    CascadeMux I__13699 (
            .O(N__57833),
            .I(N__57827));
    LocalMux I__13698 (
            .O(N__57830),
            .I(N__57823));
    InMux I__13697 (
            .O(N__57827),
            .I(N__57820));
    InMux I__13696 (
            .O(N__57826),
            .I(N__57817));
    Span12Mux_h I__13695 (
            .O(N__57823),
            .I(N__57814));
    LocalMux I__13694 (
            .O(N__57820),
            .I(N__57811));
    LocalMux I__13693 (
            .O(N__57817),
            .I(N__57808));
    Odrv12 I__13692 (
            .O(N__57814),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_1));
    Odrv12 I__13691 (
            .O(N__57811),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_1));
    Odrv4 I__13690 (
            .O(N__57808),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_1));
    InMux I__13689 (
            .O(N__57801),
            .I(N__57796));
    InMux I__13688 (
            .O(N__57800),
            .I(N__57793));
    InMux I__13687 (
            .O(N__57799),
            .I(N__57790));
    LocalMux I__13686 (
            .O(N__57796),
            .I(N__57787));
    LocalMux I__13685 (
            .O(N__57793),
            .I(N__57784));
    LocalMux I__13684 (
            .O(N__57790),
            .I(N__57781));
    Span4Mux_v I__13683 (
            .O(N__57787),
            .I(N__57778));
    Span4Mux_v I__13682 (
            .O(N__57784),
            .I(N__57775));
    Span4Mux_h I__13681 (
            .O(N__57781),
            .I(N__57772));
    Span4Mux_h I__13680 (
            .O(N__57778),
            .I(N__57769));
    Span4Mux_h I__13679 (
            .O(N__57775),
            .I(N__57764));
    Span4Mux_h I__13678 (
            .O(N__57772),
            .I(N__57764));
    Span4Mux_h I__13677 (
            .O(N__57769),
            .I(N__57761));
    Span4Mux_h I__13676 (
            .O(N__57764),
            .I(N__57758));
    Odrv4 I__13675 (
            .O(N__57761),
            .I(cemf_module_64ch_ctrl_inst1_data_config_1));
    Odrv4 I__13674 (
            .O(N__57758),
            .I(cemf_module_64ch_ctrl_inst1_data_config_1));
    InMux I__13673 (
            .O(N__57753),
            .I(N__57750));
    LocalMux I__13672 (
            .O(N__57750),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1776 ));
    CascadeMux I__13671 (
            .O(N__57747),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0_cascade_ ));
    InMux I__13670 (
            .O(N__57744),
            .I(N__57740));
    InMux I__13669 (
            .O(N__57743),
            .I(N__57737));
    LocalMux I__13668 (
            .O(N__57740),
            .I(N__57731));
    LocalMux I__13667 (
            .O(N__57737),
            .I(N__57731));
    InMux I__13666 (
            .O(N__57736),
            .I(N__57728));
    Span4Mux_v I__13665 (
            .O(N__57731),
            .I(N__57723));
    LocalMux I__13664 (
            .O(N__57728),
            .I(N__57723));
    Span4Mux_v I__13663 (
            .O(N__57723),
            .I(N__57720));
    Sp12to4 I__13662 (
            .O(N__57720),
            .I(N__57715));
    InMux I__13661 (
            .O(N__57719),
            .I(N__57710));
    InMux I__13660 (
            .O(N__57718),
            .I(N__57710));
    Odrv12 I__13659 (
            .O(N__57715),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11 ));
    LocalMux I__13658 (
            .O(N__57710),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11 ));
    InMux I__13657 (
            .O(N__57705),
            .I(N__57702));
    LocalMux I__13656 (
            .O(N__57702),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_209 ));
    IoInMux I__13655 (
            .O(N__57699),
            .I(N__57696));
    LocalMux I__13654 (
            .O(N__57696),
            .I(N__57693));
    IoSpan4Mux I__13653 (
            .O(N__57693),
            .I(N__57690));
    Span4Mux_s1_h I__13652 (
            .O(N__57690),
            .I(N__57687));
    Span4Mux_h I__13651 (
            .O(N__57687),
            .I(N__57682));
    InMux I__13650 (
            .O(N__57686),
            .I(N__57679));
    InMux I__13649 (
            .O(N__57685),
            .I(N__57676));
    Span4Mux_h I__13648 (
            .O(N__57682),
            .I(N__57671));
    LocalMux I__13647 (
            .O(N__57679),
            .I(N__57671));
    LocalMux I__13646 (
            .O(N__57676),
            .I(N__57668));
    Span4Mux_v I__13645 (
            .O(N__57671),
            .I(N__57665));
    Span4Mux_v I__13644 (
            .O(N__57668),
            .I(N__57662));
    Span4Mux_v I__13643 (
            .O(N__57665),
            .I(N__57659));
    Span4Mux_h I__13642 (
            .O(N__57662),
            .I(N__57656));
    Sp12to4 I__13641 (
            .O(N__57659),
            .I(N__57653));
    Sp12to4 I__13640 (
            .O(N__57656),
            .I(N__57650));
    Span12Mux_h I__13639 (
            .O(N__57653),
            .I(N__57645));
    Span12Mux_v I__13638 (
            .O(N__57650),
            .I(N__57645));
    Odrv12 I__13637 (
            .O(N__57645),
            .I(s_sda_i));
    InMux I__13636 (
            .O(N__57642),
            .I(N__57639));
    LocalMux I__13635 (
            .O(N__57639),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_0 ));
    InMux I__13634 (
            .O(N__57636),
            .I(N__57633));
    LocalMux I__13633 (
            .O(N__57633),
            .I(N__57629));
    InMux I__13632 (
            .O(N__57632),
            .I(N__57624));
    Span4Mux_v I__13631 (
            .O(N__57629),
            .I(N__57621));
    InMux I__13630 (
            .O(N__57628),
            .I(N__57615));
    InMux I__13629 (
            .O(N__57627),
            .I(N__57612));
    LocalMux I__13628 (
            .O(N__57624),
            .I(N__57609));
    Span4Mux_h I__13627 (
            .O(N__57621),
            .I(N__57605));
    InMux I__13626 (
            .O(N__57620),
            .I(N__57602));
    InMux I__13625 (
            .O(N__57619),
            .I(N__57598));
    InMux I__13624 (
            .O(N__57618),
            .I(N__57595));
    LocalMux I__13623 (
            .O(N__57615),
            .I(N__57592));
    LocalMux I__13622 (
            .O(N__57612),
            .I(N__57589));
    Span4Mux_h I__13621 (
            .O(N__57609),
            .I(N__57586));
    CascadeMux I__13620 (
            .O(N__57608),
            .I(N__57583));
    Span4Mux_h I__13619 (
            .O(N__57605),
            .I(N__57580));
    LocalMux I__13618 (
            .O(N__57602),
            .I(N__57577));
    InMux I__13617 (
            .O(N__57601),
            .I(N__57574));
    LocalMux I__13616 (
            .O(N__57598),
            .I(N__57571));
    LocalMux I__13615 (
            .O(N__57595),
            .I(N__57568));
    Span4Mux_h I__13614 (
            .O(N__57592),
            .I(N__57561));
    Span4Mux_h I__13613 (
            .O(N__57589),
            .I(N__57561));
    Span4Mux_h I__13612 (
            .O(N__57586),
            .I(N__57561));
    InMux I__13611 (
            .O(N__57583),
            .I(N__57558));
    Span4Mux_h I__13610 (
            .O(N__57580),
            .I(N__57555));
    Odrv12 I__13609 (
            .O(N__57577),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    LocalMux I__13608 (
            .O(N__57574),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    Odrv4 I__13607 (
            .O(N__57571),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    Odrv12 I__13606 (
            .O(N__57568),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    Odrv4 I__13605 (
            .O(N__57561),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    LocalMux I__13604 (
            .O(N__57558),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    Odrv4 I__13603 (
            .O(N__57555),
            .I(I2C_top_level_inst1_s_data_oreg_16));
    InMux I__13602 (
            .O(N__57540),
            .I(N__57537));
    LocalMux I__13601 (
            .O(N__57537),
            .I(N__57531));
    InMux I__13600 (
            .O(N__57536),
            .I(N__57528));
    InMux I__13599 (
            .O(N__57535),
            .I(N__57525));
    InMux I__13598 (
            .O(N__57534),
            .I(N__57521));
    Span4Mux_v I__13597 (
            .O(N__57531),
            .I(N__57513));
    LocalMux I__13596 (
            .O(N__57528),
            .I(N__57513));
    LocalMux I__13595 (
            .O(N__57525),
            .I(N__57513));
    InMux I__13594 (
            .O(N__57524),
            .I(N__57510));
    LocalMux I__13593 (
            .O(N__57521),
            .I(N__57506));
    InMux I__13592 (
            .O(N__57520),
            .I(N__57503));
    Span4Mux_h I__13591 (
            .O(N__57513),
            .I(N__57500));
    LocalMux I__13590 (
            .O(N__57510),
            .I(N__57497));
    InMux I__13589 (
            .O(N__57509),
            .I(N__57493));
    Span4Mux_v I__13588 (
            .O(N__57506),
            .I(N__57490));
    LocalMux I__13587 (
            .O(N__57503),
            .I(N__57487));
    Span4Mux_v I__13586 (
            .O(N__57500),
            .I(N__57482));
    Span4Mux_v I__13585 (
            .O(N__57497),
            .I(N__57482));
    InMux I__13584 (
            .O(N__57496),
            .I(N__57479));
    LocalMux I__13583 (
            .O(N__57493),
            .I(N__57476));
    Span4Mux_h I__13582 (
            .O(N__57490),
            .I(N__57472));
    Span4Mux_v I__13581 (
            .O(N__57487),
            .I(N__57469));
    Sp12to4 I__13580 (
            .O(N__57482),
            .I(N__57464));
    LocalMux I__13579 (
            .O(N__57479),
            .I(N__57464));
    Span4Mux_v I__13578 (
            .O(N__57476),
            .I(N__57461));
    CascadeMux I__13577 (
            .O(N__57475),
            .I(N__57458));
    Span4Mux_h I__13576 (
            .O(N__57472),
            .I(N__57453));
    Span4Mux_v I__13575 (
            .O(N__57469),
            .I(N__57453));
    Span12Mux_h I__13574 (
            .O(N__57464),
            .I(N__57450));
    Span4Mux_h I__13573 (
            .O(N__57461),
            .I(N__57447));
    InMux I__13572 (
            .O(N__57458),
            .I(N__57444));
    Odrv4 I__13571 (
            .O(N__57453),
            .I(I2C_top_level_inst1_s_data_oreg_15));
    Odrv12 I__13570 (
            .O(N__57450),
            .I(I2C_top_level_inst1_s_data_oreg_15));
    Odrv4 I__13569 (
            .O(N__57447),
            .I(I2C_top_level_inst1_s_data_oreg_15));
    LocalMux I__13568 (
            .O(N__57444),
            .I(I2C_top_level_inst1_s_data_oreg_15));
    InMux I__13567 (
            .O(N__57435),
            .I(N__57432));
    LocalMux I__13566 (
            .O(N__57432),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_15 ));
    InMux I__13565 (
            .O(N__57429),
            .I(N__57426));
    LocalMux I__13564 (
            .O(N__57426),
            .I(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_16 ));
    InMux I__13563 (
            .O(N__57423),
            .I(N__57420));
    LocalMux I__13562 (
            .O(N__57420),
            .I(N__57415));
    InMux I__13561 (
            .O(N__57419),
            .I(N__57409));
    InMux I__13560 (
            .O(N__57418),
            .I(N__57406));
    Span4Mux_v I__13559 (
            .O(N__57415),
            .I(N__57403));
    InMux I__13558 (
            .O(N__57414),
            .I(N__57400));
    InMux I__13557 (
            .O(N__57413),
            .I(N__57397));
    InMux I__13556 (
            .O(N__57412),
            .I(N__57394));
    LocalMux I__13555 (
            .O(N__57409),
            .I(N__57389));
    LocalMux I__13554 (
            .O(N__57406),
            .I(N__57386));
    Span4Mux_h I__13553 (
            .O(N__57403),
            .I(N__57383));
    LocalMux I__13552 (
            .O(N__57400),
            .I(N__57380));
    LocalMux I__13551 (
            .O(N__57397),
            .I(N__57375));
    LocalMux I__13550 (
            .O(N__57394),
            .I(N__57375));
    InMux I__13549 (
            .O(N__57393),
            .I(N__57371));
    InMux I__13548 (
            .O(N__57392),
            .I(N__57368));
    Span4Mux_v I__13547 (
            .O(N__57389),
            .I(N__57361));
    Span4Mux_v I__13546 (
            .O(N__57386),
            .I(N__57361));
    Span4Mux_v I__13545 (
            .O(N__57383),
            .I(N__57361));
    Span4Mux_v I__13544 (
            .O(N__57380),
            .I(N__57356));
    Span4Mux_v I__13543 (
            .O(N__57375),
            .I(N__57356));
    CascadeMux I__13542 (
            .O(N__57374),
            .I(N__57353));
    LocalMux I__13541 (
            .O(N__57371),
            .I(N__57350));
    LocalMux I__13540 (
            .O(N__57368),
            .I(N__57343));
    Sp12to4 I__13539 (
            .O(N__57361),
            .I(N__57343));
    Sp12to4 I__13538 (
            .O(N__57356),
            .I(N__57343));
    InMux I__13537 (
            .O(N__57353),
            .I(N__57340));
    Span4Mux_h I__13536 (
            .O(N__57350),
            .I(N__57337));
    Odrv12 I__13535 (
            .O(N__57343),
            .I(I2C_top_level_inst1_s_data_oreg_17));
    LocalMux I__13534 (
            .O(N__57340),
            .I(I2C_top_level_inst1_s_data_oreg_17));
    Odrv4 I__13533 (
            .O(N__57337),
            .I(I2C_top_level_inst1_s_data_oreg_17));
    InMux I__13532 (
            .O(N__57330),
            .I(N__57327));
    LocalMux I__13531 (
            .O(N__57327),
            .I(N__57324));
    Span4Mux_h I__13530 (
            .O(N__57324),
            .I(N__57320));
    InMux I__13529 (
            .O(N__57323),
            .I(N__57316));
    Span4Mux_h I__13528 (
            .O(N__57320),
            .I(N__57313));
    InMux I__13527 (
            .O(N__57319),
            .I(N__57310));
    LocalMux I__13526 (
            .O(N__57316),
            .I(N__57307));
    Odrv4 I__13525 (
            .O(N__57313),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_19));
    LocalMux I__13524 (
            .O(N__57310),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_19));
    Odrv12 I__13523 (
            .O(N__57307),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_19));
    InMux I__13522 (
            .O(N__57300),
            .I(N__57297));
    LocalMux I__13521 (
            .O(N__57297),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_211 ));
    CascadeMux I__13520 (
            .O(N__57294),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1653_cascade_ ));
    CascadeMux I__13519 (
            .O(N__57291),
            .I(N__57288));
    InMux I__13518 (
            .O(N__57288),
            .I(N__57284));
    InMux I__13517 (
            .O(N__57287),
            .I(N__57281));
    LocalMux I__13516 (
            .O(N__57284),
            .I(N__57278));
    LocalMux I__13515 (
            .O(N__57281),
            .I(N__57275));
    Span4Mux_v I__13514 (
            .O(N__57278),
            .I(N__57272));
    Odrv4 I__13513 (
            .O(N__57275),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0 ));
    Odrv4 I__13512 (
            .O(N__57272),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0 ));
    CascadeMux I__13511 (
            .O(N__57267),
            .I(N__57264));
    InMux I__13510 (
            .O(N__57264),
            .I(N__57261));
    LocalMux I__13509 (
            .O(N__57261),
            .I(N__57258));
    Odrv4 I__13508 (
            .O(N__57258),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_122_0 ));
    InMux I__13507 (
            .O(N__57255),
            .I(N__57252));
    LocalMux I__13506 (
            .O(N__57252),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_208 ));
    InMux I__13505 (
            .O(N__57249),
            .I(N__57243));
    InMux I__13504 (
            .O(N__57248),
            .I(N__57243));
    LocalMux I__13503 (
            .O(N__57243),
            .I(N__57239));
    InMux I__13502 (
            .O(N__57242),
            .I(N__57234));
    Span4Mux_h I__13501 (
            .O(N__57239),
            .I(N__57231));
    InMux I__13500 (
            .O(N__57238),
            .I(N__57228));
    InMux I__13499 (
            .O(N__57237),
            .I(N__57224));
    LocalMux I__13498 (
            .O(N__57234),
            .I(N__57220));
    Span4Mux_h I__13497 (
            .O(N__57231),
            .I(N__57217));
    LocalMux I__13496 (
            .O(N__57228),
            .I(N__57213));
    CascadeMux I__13495 (
            .O(N__57227),
            .I(N__57210));
    LocalMux I__13494 (
            .O(N__57224),
            .I(N__57205));
    InMux I__13493 (
            .O(N__57223),
            .I(N__57202));
    Span4Mux_h I__13492 (
            .O(N__57220),
            .I(N__57197));
    Span4Mux_v I__13491 (
            .O(N__57217),
            .I(N__57197));
    CascadeMux I__13490 (
            .O(N__57216),
            .I(N__57194));
    Span4Mux_h I__13489 (
            .O(N__57213),
            .I(N__57191));
    InMux I__13488 (
            .O(N__57210),
            .I(N__57188));
    InMux I__13487 (
            .O(N__57209),
            .I(N__57185));
    InMux I__13486 (
            .O(N__57208),
            .I(N__57182));
    Span4Mux_v I__13485 (
            .O(N__57205),
            .I(N__57179));
    LocalMux I__13484 (
            .O(N__57202),
            .I(N__57176));
    Span4Mux_h I__13483 (
            .O(N__57197),
            .I(N__57173));
    InMux I__13482 (
            .O(N__57194),
            .I(N__57170));
    Span4Mux_h I__13481 (
            .O(N__57191),
            .I(N__57167));
    LocalMux I__13480 (
            .O(N__57188),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    LocalMux I__13479 (
            .O(N__57185),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    LocalMux I__13478 (
            .O(N__57182),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    Odrv4 I__13477 (
            .O(N__57179),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    Odrv12 I__13476 (
            .O(N__57176),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    Odrv4 I__13475 (
            .O(N__57173),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    LocalMux I__13474 (
            .O(N__57170),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    Odrv4 I__13473 (
            .O(N__57167),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ));
    CascadeMux I__13472 (
            .O(N__57150),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0_cascade_ ));
    CascadeMux I__13471 (
            .O(N__57147),
            .I(N__57143));
    InMux I__13470 (
            .O(N__57146),
            .I(N__57138));
    InMux I__13469 (
            .O(N__57143),
            .I(N__57138));
    LocalMux I__13468 (
            .O(N__57138),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_239 ));
    CascadeMux I__13467 (
            .O(N__57135),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_239_cascade_ ));
    InMux I__13466 (
            .O(N__57132),
            .I(N__57128));
    InMux I__13465 (
            .O(N__57131),
            .I(N__57125));
    LocalMux I__13464 (
            .O(N__57128),
            .I(N__57120));
    LocalMux I__13463 (
            .O(N__57125),
            .I(N__57117));
    InMux I__13462 (
            .O(N__57124),
            .I(N__57114));
    InMux I__13461 (
            .O(N__57123),
            .I(N__57111));
    Span4Mux_h I__13460 (
            .O(N__57120),
            .I(N__57104));
    Span4Mux_h I__13459 (
            .O(N__57117),
            .I(N__57104));
    LocalMux I__13458 (
            .O(N__57114),
            .I(N__57104));
    LocalMux I__13457 (
            .O(N__57111),
            .I(N__57101));
    Span4Mux_v I__13456 (
            .O(N__57104),
            .I(N__57098));
    Odrv4 I__13455 (
            .O(N__57101),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_294 ));
    Odrv4 I__13454 (
            .O(N__57098),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_294 ));
    CascadeMux I__13453 (
            .O(N__57093),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_1_0_0_cascade_ ));
    InMux I__13452 (
            .O(N__57090),
            .I(N__57086));
    InMux I__13451 (
            .O(N__57089),
            .I(N__57083));
    LocalMux I__13450 (
            .O(N__57086),
            .I(N__57079));
    LocalMux I__13449 (
            .O(N__57083),
            .I(N__57076));
    InMux I__13448 (
            .O(N__57082),
            .I(N__57073));
    Odrv4 I__13447 (
            .O(N__57079),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2 ));
    Odrv12 I__13446 (
            .O(N__57076),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2 ));
    LocalMux I__13445 (
            .O(N__57073),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2 ));
    InMux I__13444 (
            .O(N__57066),
            .I(N__57063));
    LocalMux I__13443 (
            .O(N__57063),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_0_0 ));
    CascadeMux I__13442 (
            .O(N__57060),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1446_cascade_ ));
    CascadeMux I__13441 (
            .O(N__57057),
            .I(N__57053));
    InMux I__13440 (
            .O(N__57056),
            .I(N__57050));
    InMux I__13439 (
            .O(N__57053),
            .I(N__57047));
    LocalMux I__13438 (
            .O(N__57050),
            .I(N__57044));
    LocalMux I__13437 (
            .O(N__57047),
            .I(N__57041));
    Span4Mux_v I__13436 (
            .O(N__57044),
            .I(N__57036));
    Span4Mux_v I__13435 (
            .O(N__57041),
            .I(N__57036));
    Span4Mux_h I__13434 (
            .O(N__57036),
            .I(N__57033));
    Odrv4 I__13433 (
            .O(N__57033),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_291 ));
    InMux I__13432 (
            .O(N__57030),
            .I(N__57023));
    InMux I__13431 (
            .O(N__57029),
            .I(N__57023));
    InMux I__13430 (
            .O(N__57028),
            .I(N__57020));
    LocalMux I__13429 (
            .O(N__57023),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24 ));
    LocalMux I__13428 (
            .O(N__57020),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24 ));
    CascadeMux I__13427 (
            .O(N__57015),
            .I(N__57009));
    CascadeMux I__13426 (
            .O(N__57014),
            .I(N__57006));
    CascadeMux I__13425 (
            .O(N__57013),
            .I(N__57003));
    InMux I__13424 (
            .O(N__57012),
            .I(N__56999));
    InMux I__13423 (
            .O(N__57009),
            .I(N__56996));
    InMux I__13422 (
            .O(N__57006),
            .I(N__56990));
    InMux I__13421 (
            .O(N__57003),
            .I(N__56985));
    InMux I__13420 (
            .O(N__57002),
            .I(N__56985));
    LocalMux I__13419 (
            .O(N__56999),
            .I(N__56980));
    LocalMux I__13418 (
            .O(N__56996),
            .I(N__56980));
    InMux I__13417 (
            .O(N__56995),
            .I(N__56973));
    InMux I__13416 (
            .O(N__56994),
            .I(N__56973));
    InMux I__13415 (
            .O(N__56993),
            .I(N__56973));
    LocalMux I__13414 (
            .O(N__56990),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25 ));
    LocalMux I__13413 (
            .O(N__56985),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25 ));
    Odrv4 I__13412 (
            .O(N__56980),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25 ));
    LocalMux I__13411 (
            .O(N__56973),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25 ));
    InMux I__13410 (
            .O(N__56964),
            .I(N__56961));
    LocalMux I__13409 (
            .O(N__56961),
            .I(N__56958));
    Odrv4 I__13408 (
            .O(N__56958),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_0_1 ));
    CascadeMux I__13407 (
            .O(N__56955),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_232_cascade_ ));
    CascadeMux I__13406 (
            .O(N__56952),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_2_1_cascade_ ));
    InMux I__13405 (
            .O(N__56949),
            .I(N__56943));
    InMux I__13404 (
            .O(N__56948),
            .I(N__56940));
    InMux I__13403 (
            .O(N__56947),
            .I(N__56935));
    InMux I__13402 (
            .O(N__56946),
            .I(N__56935));
    LocalMux I__13401 (
            .O(N__56943),
            .I(N__56932));
    LocalMux I__13400 (
            .O(N__56940),
            .I(N__56929));
    LocalMux I__13399 (
            .O(N__56935),
            .I(N__56926));
    Span4Mux_h I__13398 (
            .O(N__56932),
            .I(N__56921));
    Span4Mux_h I__13397 (
            .O(N__56929),
            .I(N__56921));
    Odrv12 I__13396 (
            .O(N__56926),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4));
    Odrv4 I__13395 (
            .O(N__56921),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4));
    InMux I__13394 (
            .O(N__56916),
            .I(N__56910));
    InMux I__13393 (
            .O(N__56915),
            .I(N__56910));
    LocalMux I__13392 (
            .O(N__56910),
            .I(N__56905));
    InMux I__13391 (
            .O(N__56909),
            .I(N__56902));
    InMux I__13390 (
            .O(N__56908),
            .I(N__56899));
    Span4Mux_h I__13389 (
            .O(N__56905),
            .I(N__56896));
    LocalMux I__13388 (
            .O(N__56902),
            .I(N__56889));
    LocalMux I__13387 (
            .O(N__56899),
            .I(N__56889));
    Span4Mux_v I__13386 (
            .O(N__56896),
            .I(N__56889));
    Odrv4 I__13385 (
            .O(N__56889),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_20));
    InMux I__13384 (
            .O(N__56886),
            .I(N__56882));
    InMux I__13383 (
            .O(N__56885),
            .I(N__56879));
    LocalMux I__13382 (
            .O(N__56882),
            .I(N__56873));
    LocalMux I__13381 (
            .O(N__56879),
            .I(N__56873));
    InMux I__13380 (
            .O(N__56878),
            .I(N__56870));
    Span12Mux_h I__13379 (
            .O(N__56873),
            .I(N__56863));
    LocalMux I__13378 (
            .O(N__56870),
            .I(N__56863));
    InMux I__13377 (
            .O(N__56869),
            .I(N__56858));
    InMux I__13376 (
            .O(N__56868),
            .I(N__56858));
    Odrv12 I__13375 (
            .O(N__56863),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12));
    LocalMux I__13374 (
            .O(N__56858),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12));
    InMux I__13373 (
            .O(N__56853),
            .I(N__56850));
    LocalMux I__13372 (
            .O(N__56850),
            .I(N__56847));
    Odrv4 I__13371 (
            .O(N__56847),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_4_0 ));
    CascadeMux I__13370 (
            .O(N__56844),
            .I(N__56840));
    InMux I__13369 (
            .O(N__56843),
            .I(N__56837));
    InMux I__13368 (
            .O(N__56840),
            .I(N__56834));
    LocalMux I__13367 (
            .O(N__56837),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_232 ));
    LocalMux I__13366 (
            .O(N__56834),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_232 ));
    InMux I__13365 (
            .O(N__56829),
            .I(N__56825));
    InMux I__13364 (
            .O(N__56828),
            .I(N__56822));
    LocalMux I__13363 (
            .O(N__56825),
            .I(N__56819));
    LocalMux I__13362 (
            .O(N__56822),
            .I(N__56812));
    Span4Mux_h I__13361 (
            .O(N__56819),
            .I(N__56809));
    InMux I__13360 (
            .O(N__56818),
            .I(N__56806));
    InMux I__13359 (
            .O(N__56817),
            .I(N__56799));
    InMux I__13358 (
            .O(N__56816),
            .I(N__56799));
    InMux I__13357 (
            .O(N__56815),
            .I(N__56799));
    Span4Mux_h I__13356 (
            .O(N__56812),
            .I(N__56796));
    Odrv4 I__13355 (
            .O(N__56809),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22));
    LocalMux I__13354 (
            .O(N__56806),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22));
    LocalMux I__13353 (
            .O(N__56799),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22));
    Odrv4 I__13352 (
            .O(N__56796),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22));
    InMux I__13351 (
            .O(N__56787),
            .I(N__56784));
    LocalMux I__13350 (
            .O(N__56784),
            .I(N__56781));
    Odrv12 I__13349 (
            .O(N__56781),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_1_0 ));
    CascadeMux I__13348 (
            .O(N__56778),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_2_0_cascade_ ));
    InMux I__13347 (
            .O(N__56775),
            .I(N__56772));
    LocalMux I__13346 (
            .O(N__56772),
            .I(N__56767));
    InMux I__13345 (
            .O(N__56771),
            .I(N__56762));
    InMux I__13344 (
            .O(N__56770),
            .I(N__56762));
    Odrv4 I__13343 (
            .O(N__56767),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_231 ));
    LocalMux I__13342 (
            .O(N__56762),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_231 ));
    CascadeMux I__13341 (
            .O(N__56757),
            .I(N__56754));
    InMux I__13340 (
            .O(N__56754),
            .I(N__56751));
    LocalMux I__13339 (
            .O(N__56751),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_212 ));
    InMux I__13338 (
            .O(N__56748),
            .I(N__56745));
    LocalMux I__13337 (
            .O(N__56745),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_288 ));
    CascadeMux I__13336 (
            .O(N__56742),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_288_cascade_ ));
    InMux I__13335 (
            .O(N__56739),
            .I(N__56736));
    LocalMux I__13334 (
            .O(N__56736),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_23 ));
    InMux I__13333 (
            .O(N__56733),
            .I(N__56730));
    LocalMux I__13332 (
            .O(N__56730),
            .I(N__56722));
    InMux I__13331 (
            .O(N__56729),
            .I(N__56719));
    InMux I__13330 (
            .O(N__56728),
            .I(N__56713));
    InMux I__13329 (
            .O(N__56727),
            .I(N__56713));
    InMux I__13328 (
            .O(N__56726),
            .I(N__56708));
    InMux I__13327 (
            .O(N__56725),
            .I(N__56708));
    Span4Mux_v I__13326 (
            .O(N__56722),
            .I(N__56705));
    LocalMux I__13325 (
            .O(N__56719),
            .I(N__56702));
    InMux I__13324 (
            .O(N__56718),
            .I(N__56697));
    LocalMux I__13323 (
            .O(N__56713),
            .I(N__56692));
    LocalMux I__13322 (
            .O(N__56708),
            .I(N__56692));
    Span4Mux_h I__13321 (
            .O(N__56705),
            .I(N__56687));
    Span4Mux_h I__13320 (
            .O(N__56702),
            .I(N__56687));
    InMux I__13319 (
            .O(N__56701),
            .I(N__56684));
    InMux I__13318 (
            .O(N__56700),
            .I(N__56681));
    LocalMux I__13317 (
            .O(N__56697),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ));
    Odrv4 I__13316 (
            .O(N__56692),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ));
    Odrv4 I__13315 (
            .O(N__56687),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ));
    LocalMux I__13314 (
            .O(N__56684),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ));
    LocalMux I__13313 (
            .O(N__56681),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ));
    InMux I__13312 (
            .O(N__56670),
            .I(N__56667));
    LocalMux I__13311 (
            .O(N__56667),
            .I(N__56664));
    Odrv4 I__13310 (
            .O(N__56664),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_115 ));
    InMux I__13309 (
            .O(N__56661),
            .I(N__56657));
    InMux I__13308 (
            .O(N__56660),
            .I(N__56654));
    LocalMux I__13307 (
            .O(N__56657),
            .I(N__56651));
    LocalMux I__13306 (
            .O(N__56654),
            .I(N__56646));
    Span4Mux_h I__13305 (
            .O(N__56651),
            .I(N__56643));
    InMux I__13304 (
            .O(N__56650),
            .I(N__56638));
    InMux I__13303 (
            .O(N__56649),
            .I(N__56638));
    Odrv4 I__13302 (
            .O(N__56646),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16 ));
    Odrv4 I__13301 (
            .O(N__56643),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16 ));
    LocalMux I__13300 (
            .O(N__56638),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16 ));
    CascadeMux I__13299 (
            .O(N__56631),
            .I(N__56628));
    InMux I__13298 (
            .O(N__56628),
            .I(N__56622));
    InMux I__13297 (
            .O(N__56627),
            .I(N__56622));
    LocalMux I__13296 (
            .O(N__56622),
            .I(N__56617));
    InMux I__13295 (
            .O(N__56621),
            .I(N__56612));
    InMux I__13294 (
            .O(N__56620),
            .I(N__56612));
    Odrv4 I__13293 (
            .O(N__56617),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2 ));
    LocalMux I__13292 (
            .O(N__56612),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2 ));
    InMux I__13291 (
            .O(N__56607),
            .I(N__56601));
    InMux I__13290 (
            .O(N__56606),
            .I(N__56601));
    LocalMux I__13289 (
            .O(N__56601),
            .I(N__56598));
    Span4Mux_h I__13288 (
            .O(N__56598),
            .I(N__56595));
    Span4Mux_v I__13287 (
            .O(N__56595),
            .I(N__56588));
    InMux I__13286 (
            .O(N__56594),
            .I(N__56585));
    InMux I__13285 (
            .O(N__56593),
            .I(N__56578));
    InMux I__13284 (
            .O(N__56592),
            .I(N__56578));
    CascadeMux I__13283 (
            .O(N__56591),
            .I(N__56575));
    Span4Mux_v I__13282 (
            .O(N__56588),
            .I(N__56569));
    LocalMux I__13281 (
            .O(N__56585),
            .I(N__56569));
    InMux I__13280 (
            .O(N__56584),
            .I(N__56564));
    InMux I__13279 (
            .O(N__56583),
            .I(N__56564));
    LocalMux I__13278 (
            .O(N__56578),
            .I(N__56561));
    InMux I__13277 (
            .O(N__56575),
            .I(N__56554));
    InMux I__13276 (
            .O(N__56574),
            .I(N__56554));
    Span4Mux_v I__13275 (
            .O(N__56569),
            .I(N__56549));
    LocalMux I__13274 (
            .O(N__56564),
            .I(N__56549));
    Span4Mux_h I__13273 (
            .O(N__56561),
            .I(N__56546));
    InMux I__13272 (
            .O(N__56560),
            .I(N__56543));
    InMux I__13271 (
            .O(N__56559),
            .I(N__56540));
    LocalMux I__13270 (
            .O(N__56554),
            .I(N__56537));
    Span4Mux_h I__13269 (
            .O(N__56549),
            .I(N__56534));
    Span4Mux_h I__13268 (
            .O(N__56546),
            .I(N__56529));
    LocalMux I__13267 (
            .O(N__56543),
            .I(N__56529));
    LocalMux I__13266 (
            .O(N__56540),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1 ));
    Odrv4 I__13265 (
            .O(N__56537),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1 ));
    Odrv4 I__13264 (
            .O(N__56534),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1 ));
    Odrv4 I__13263 (
            .O(N__56529),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1 ));
    CascadeMux I__13262 (
            .O(N__56520),
            .I(N__56517));
    InMux I__13261 (
            .O(N__56517),
            .I(N__56513));
    InMux I__13260 (
            .O(N__56516),
            .I(N__56508));
    LocalMux I__13259 (
            .O(N__56513),
            .I(N__56505));
    InMux I__13258 (
            .O(N__56512),
            .I(N__56500));
    InMux I__13257 (
            .O(N__56511),
            .I(N__56500));
    LocalMux I__13256 (
            .O(N__56508),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_904 ));
    Odrv4 I__13255 (
            .O(N__56505),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_904 ));
    LocalMux I__13254 (
            .O(N__56500),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_904 ));
    CascadeMux I__13253 (
            .O(N__56493),
            .I(N__56490));
    InMux I__13252 (
            .O(N__56490),
            .I(N__56486));
    InMux I__13251 (
            .O(N__56489),
            .I(N__56483));
    LocalMux I__13250 (
            .O(N__56486),
            .I(N__56480));
    LocalMux I__13249 (
            .O(N__56483),
            .I(N__56477));
    Span4Mux_h I__13248 (
            .O(N__56480),
            .I(N__56472));
    Span4Mux_h I__13247 (
            .O(N__56477),
            .I(N__56472));
    Odrv4 I__13246 (
            .O(N__56472),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_2 ));
    InMux I__13245 (
            .O(N__56469),
            .I(N__56465));
    InMux I__13244 (
            .O(N__56468),
            .I(N__56462));
    LocalMux I__13243 (
            .O(N__56465),
            .I(N__56459));
    LocalMux I__13242 (
            .O(N__56462),
            .I(N__56456));
    Span4Mux_v I__13241 (
            .O(N__56459),
            .I(N__56453));
    Odrv4 I__13240 (
            .O(N__56456),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1 ));
    Odrv4 I__13239 (
            .O(N__56453),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1 ));
    InMux I__13238 (
            .O(N__56448),
            .I(N__56443));
    InMux I__13237 (
            .O(N__56447),
            .I(N__56434));
    InMux I__13236 (
            .O(N__56446),
            .I(N__56434));
    LocalMux I__13235 (
            .O(N__56443),
            .I(N__56431));
    InMux I__13234 (
            .O(N__56442),
            .I(N__56428));
    InMux I__13233 (
            .O(N__56441),
            .I(N__56425));
    CascadeMux I__13232 (
            .O(N__56440),
            .I(N__56422));
    InMux I__13231 (
            .O(N__56439),
            .I(N__56419));
    LocalMux I__13230 (
            .O(N__56434),
            .I(N__56416));
    Span4Mux_v I__13229 (
            .O(N__56431),
            .I(N__56411));
    LocalMux I__13228 (
            .O(N__56428),
            .I(N__56411));
    LocalMux I__13227 (
            .O(N__56425),
            .I(N__56408));
    InMux I__13226 (
            .O(N__56422),
            .I(N__56403));
    LocalMux I__13225 (
            .O(N__56419),
            .I(N__56394));
    Span4Mux_v I__13224 (
            .O(N__56416),
            .I(N__56394));
    Span4Mux_v I__13223 (
            .O(N__56411),
            .I(N__56394));
    Span4Mux_h I__13222 (
            .O(N__56408),
            .I(N__56394));
    InMux I__13221 (
            .O(N__56407),
            .I(N__56389));
    InMux I__13220 (
            .O(N__56406),
            .I(N__56389));
    LocalMux I__13219 (
            .O(N__56403),
            .I(N__56384));
    Span4Mux_h I__13218 (
            .O(N__56394),
            .I(N__56384));
    LocalMux I__13217 (
            .O(N__56389),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26 ));
    Odrv4 I__13216 (
            .O(N__56384),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26 ));
    CascadeMux I__13215 (
            .O(N__56379),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un30_i_a2_9_a2_4_a2_0_1_2_cascade_ ));
    InMux I__13214 (
            .O(N__56376),
            .I(N__56373));
    LocalMux I__13213 (
            .O(N__56373),
            .I(N__56370));
    Span12Mux_h I__13212 (
            .O(N__56370),
            .I(N__56367));
    Odrv12 I__13211 (
            .O(N__56367),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1446 ));
    CascadeMux I__13210 (
            .O(N__56364),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0_cascade_ ));
    InMux I__13209 (
            .O(N__56361),
            .I(N__56354));
    InMux I__13208 (
            .O(N__56360),
            .I(N__56347));
    InMux I__13207 (
            .O(N__56359),
            .I(N__56340));
    InMux I__13206 (
            .O(N__56358),
            .I(N__56340));
    InMux I__13205 (
            .O(N__56357),
            .I(N__56340));
    LocalMux I__13204 (
            .O(N__56354),
            .I(N__56337));
    CascadeMux I__13203 (
            .O(N__56353),
            .I(N__56333));
    InMux I__13202 (
            .O(N__56352),
            .I(N__56330));
    InMux I__13201 (
            .O(N__56351),
            .I(N__56327));
    InMux I__13200 (
            .O(N__56350),
            .I(N__56324));
    LocalMux I__13199 (
            .O(N__56347),
            .I(N__56317));
    LocalMux I__13198 (
            .O(N__56340),
            .I(N__56317));
    Span4Mux_h I__13197 (
            .O(N__56337),
            .I(N__56317));
    InMux I__13196 (
            .O(N__56336),
            .I(N__56312));
    InMux I__13195 (
            .O(N__56333),
            .I(N__56312));
    LocalMux I__13194 (
            .O(N__56330),
            .I(N__56309));
    LocalMux I__13193 (
            .O(N__56327),
            .I(N__56299));
    LocalMux I__13192 (
            .O(N__56324),
            .I(N__56299));
    Sp12to4 I__13191 (
            .O(N__56317),
            .I(N__56299));
    LocalMux I__13190 (
            .O(N__56312),
            .I(N__56299));
    Span4Mux_v I__13189 (
            .O(N__56309),
            .I(N__56296));
    InMux I__13188 (
            .O(N__56308),
            .I(N__56293));
    Span12Mux_v I__13187 (
            .O(N__56299),
            .I(N__56290));
    Odrv4 I__13186 (
            .O(N__56296),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15 ));
    LocalMux I__13185 (
            .O(N__56293),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15 ));
    Odrv12 I__13184 (
            .O(N__56290),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15 ));
    CascadeMux I__13183 (
            .O(N__56283),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_5_0_cascade_ ));
    InMux I__13182 (
            .O(N__56280),
            .I(N__56277));
    LocalMux I__13181 (
            .O(N__56277),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_6_0 ));
    InMux I__13180 (
            .O(N__56274),
            .I(N__56271));
    LocalMux I__13179 (
            .O(N__56271),
            .I(N__56268));
    Span4Mux_h I__13178 (
            .O(N__56268),
            .I(N__56265));
    Odrv4 I__13177 (
            .O(N__56265),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_7_0 ));
    InMux I__13176 (
            .O(N__56262),
            .I(N__56259));
    LocalMux I__13175 (
            .O(N__56259),
            .I(N__56256));
    Odrv4 I__13174 (
            .O(N__56256),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_0 ));
    CascadeMux I__13173 (
            .O(N__56253),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_11_0_cascade_ ));
    CascadeMux I__13172 (
            .O(N__56250),
            .I(N__56242));
    InMux I__13171 (
            .O(N__56249),
            .I(N__56239));
    InMux I__13170 (
            .O(N__56248),
            .I(N__56236));
    InMux I__13169 (
            .O(N__56247),
            .I(N__56233));
    InMux I__13168 (
            .O(N__56246),
            .I(N__56229));
    CascadeMux I__13167 (
            .O(N__56245),
            .I(N__56226));
    InMux I__13166 (
            .O(N__56242),
            .I(N__56223));
    LocalMux I__13165 (
            .O(N__56239),
            .I(N__56216));
    LocalMux I__13164 (
            .O(N__56236),
            .I(N__56216));
    LocalMux I__13163 (
            .O(N__56233),
            .I(N__56216));
    InMux I__13162 (
            .O(N__56232),
            .I(N__56213));
    LocalMux I__13161 (
            .O(N__56229),
            .I(N__56210));
    InMux I__13160 (
            .O(N__56226),
            .I(N__56207));
    LocalMux I__13159 (
            .O(N__56223),
            .I(N__56204));
    Span4Mux_v I__13158 (
            .O(N__56216),
            .I(N__56201));
    LocalMux I__13157 (
            .O(N__56213),
            .I(N__56198));
    Span4Mux_h I__13156 (
            .O(N__56210),
            .I(N__56195));
    LocalMux I__13155 (
            .O(N__56207),
            .I(N__56186));
    Span4Mux_v I__13154 (
            .O(N__56204),
            .I(N__56186));
    Span4Mux_h I__13153 (
            .O(N__56201),
            .I(N__56186));
    Span4Mux_v I__13152 (
            .O(N__56198),
            .I(N__56186));
    Odrv4 I__13151 (
            .O(N__56195),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13));
    Odrv4 I__13150 (
            .O(N__56186),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13));
    InMux I__13149 (
            .O(N__56181),
            .I(N__56177));
    InMux I__13148 (
            .O(N__56180),
            .I(N__56174));
    LocalMux I__13147 (
            .O(N__56177),
            .I(N__56170));
    LocalMux I__13146 (
            .O(N__56174),
            .I(N__56167));
    InMux I__13145 (
            .O(N__56173),
            .I(N__56164));
    Span4Mux_v I__13144 (
            .O(N__56170),
            .I(N__56159));
    Span4Mux_v I__13143 (
            .O(N__56167),
            .I(N__56159));
    LocalMux I__13142 (
            .O(N__56164),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6 ));
    Odrv4 I__13141 (
            .O(N__56159),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6 ));
    CascadeMux I__13140 (
            .O(N__56154),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_23_cascade_ ));
    CascadeMux I__13139 (
            .O(N__56151),
            .I(N__56148));
    InMux I__13138 (
            .O(N__56148),
            .I(N__56141));
    InMux I__13137 (
            .O(N__56147),
            .I(N__56138));
    InMux I__13136 (
            .O(N__56146),
            .I(N__56131));
    InMux I__13135 (
            .O(N__56145),
            .I(N__56131));
    InMux I__13134 (
            .O(N__56144),
            .I(N__56131));
    LocalMux I__13133 (
            .O(N__56141),
            .I(N__56124));
    LocalMux I__13132 (
            .O(N__56138),
            .I(N__56119));
    LocalMux I__13131 (
            .O(N__56131),
            .I(N__56116));
    InMux I__13130 (
            .O(N__56130),
            .I(N__56113));
    InMux I__13129 (
            .O(N__56129),
            .I(N__56110));
    InMux I__13128 (
            .O(N__56128),
            .I(N__56105));
    InMux I__13127 (
            .O(N__56127),
            .I(N__56105));
    Span4Mux_h I__13126 (
            .O(N__56124),
            .I(N__56102));
    InMux I__13125 (
            .O(N__56123),
            .I(N__56099));
    InMux I__13124 (
            .O(N__56122),
            .I(N__56096));
    Span4Mux_h I__13123 (
            .O(N__56119),
            .I(N__56093));
    Span4Mux_h I__13122 (
            .O(N__56116),
            .I(N__56088));
    LocalMux I__13121 (
            .O(N__56113),
            .I(N__56088));
    LocalMux I__13120 (
            .O(N__56110),
            .I(N__56081));
    LocalMux I__13119 (
            .O(N__56105),
            .I(N__56081));
    Span4Mux_h I__13118 (
            .O(N__56102),
            .I(N__56081));
    LocalMux I__13117 (
            .O(N__56099),
            .I(s_paddr_I2C_8));
    LocalMux I__13116 (
            .O(N__56096),
            .I(s_paddr_I2C_8));
    Odrv4 I__13115 (
            .O(N__56093),
            .I(s_paddr_I2C_8));
    Odrv4 I__13114 (
            .O(N__56088),
            .I(s_paddr_I2C_8));
    Odrv4 I__13113 (
            .O(N__56081),
            .I(s_paddr_I2C_8));
    InMux I__13112 (
            .O(N__56070),
            .I(N__56066));
    InMux I__13111 (
            .O(N__56069),
            .I(N__56063));
    LocalMux I__13110 (
            .O(N__56066),
            .I(N__56058));
    LocalMux I__13109 (
            .O(N__56063),
            .I(N__56058));
    Span4Mux_h I__13108 (
            .O(N__56058),
            .I(N__56053));
    InMux I__13107 (
            .O(N__56057),
            .I(N__56050));
    InMux I__13106 (
            .O(N__56056),
            .I(N__56047));
    Odrv4 I__13105 (
            .O(N__56053),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0 ));
    LocalMux I__13104 (
            .O(N__56050),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0 ));
    LocalMux I__13103 (
            .O(N__56047),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0 ));
    CascadeMux I__13102 (
            .O(N__56040),
            .I(N__56037));
    InMux I__13101 (
            .O(N__56037),
            .I(N__56031));
    InMux I__13100 (
            .O(N__56036),
            .I(N__56031));
    LocalMux I__13099 (
            .O(N__56031),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_230 ));
    InMux I__13098 (
            .O(N__56028),
            .I(N__56022));
    InMux I__13097 (
            .O(N__56027),
            .I(N__56022));
    LocalMux I__13096 (
            .O(N__56022),
            .I(N__56019));
    Span4Mux_v I__13095 (
            .O(N__56019),
            .I(N__56016));
    Odrv4 I__13094 (
            .O(N__56016),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0 ));
    CascadeMux I__13093 (
            .O(N__56013),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0_cascade_ ));
    InMux I__13092 (
            .O(N__56010),
            .I(N__56007));
    LocalMux I__13091 (
            .O(N__56007),
            .I(N__56004));
    Span4Mux_h I__13090 (
            .O(N__56004),
            .I(N__56001));
    Odrv4 I__13089 (
            .O(N__56001),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_4 ));
    CascadeMux I__13088 (
            .O(N__55998),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_365_0_cascade_ ));
    CascadeMux I__13087 (
            .O(N__55995),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_4_0_a2_2_cascade_ ));
    CascadeMux I__13086 (
            .O(N__55992),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_676_0_cascade_ ));
    InMux I__13085 (
            .O(N__55989),
            .I(N__55983));
    InMux I__13084 (
            .O(N__55988),
            .I(N__55983));
    LocalMux I__13083 (
            .O(N__55983),
            .I(N__55979));
    InMux I__13082 (
            .O(N__55982),
            .I(N__55976));
    Span4Mux_v I__13081 (
            .O(N__55979),
            .I(N__55971));
    LocalMux I__13080 (
            .O(N__55976),
            .I(N__55971));
    Odrv4 I__13079 (
            .O(N__55971),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address ));
    InMux I__13078 (
            .O(N__55968),
            .I(N__55965));
    LocalMux I__13077 (
            .O(N__55965),
            .I(N__55961));
    InMux I__13076 (
            .O(N__55964),
            .I(N__55957));
    Span4Mux_v I__13075 (
            .O(N__55961),
            .I(N__55954));
    InMux I__13074 (
            .O(N__55960),
            .I(N__55951));
    LocalMux I__13073 (
            .O(N__55957),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1 ));
    Odrv4 I__13072 (
            .O(N__55954),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1 ));
    LocalMux I__13071 (
            .O(N__55951),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1 ));
    CascadeMux I__13070 (
            .O(N__55944),
            .I(N__55940));
    InMux I__13069 (
            .O(N__55943),
            .I(N__55937));
    InMux I__13068 (
            .O(N__55940),
            .I(N__55934));
    LocalMux I__13067 (
            .O(N__55937),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3 ));
    LocalMux I__13066 (
            .O(N__55934),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3 ));
    InMux I__13065 (
            .O(N__55929),
            .I(N__55924));
    InMux I__13064 (
            .O(N__55928),
            .I(N__55921));
    InMux I__13063 (
            .O(N__55927),
            .I(N__55917));
    LocalMux I__13062 (
            .O(N__55924),
            .I(N__55913));
    LocalMux I__13061 (
            .O(N__55921),
            .I(N__55910));
    InMux I__13060 (
            .O(N__55920),
            .I(N__55907));
    LocalMux I__13059 (
            .O(N__55917),
            .I(N__55904));
    InMux I__13058 (
            .O(N__55916),
            .I(N__55901));
    Span4Mux_h I__13057 (
            .O(N__55913),
            .I(N__55896));
    Span4Mux_v I__13056 (
            .O(N__55910),
            .I(N__55896));
    LocalMux I__13055 (
            .O(N__55907),
            .I(N__55893));
    Span12Mux_v I__13054 (
            .O(N__55904),
            .I(N__55890));
    LocalMux I__13053 (
            .O(N__55901),
            .I(N__55887));
    Span4Mux_v I__13052 (
            .O(N__55896),
            .I(N__55884));
    Odrv4 I__13051 (
            .O(N__55893),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16 ));
    Odrv12 I__13050 (
            .O(N__55890),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16 ));
    Odrv12 I__13049 (
            .O(N__55887),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16 ));
    Odrv4 I__13048 (
            .O(N__55884),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16 ));
    InMux I__13047 (
            .O(N__55875),
            .I(N__55872));
    LocalMux I__13046 (
            .O(N__55872),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_1 ));
    InMux I__13045 (
            .O(N__55869),
            .I(N__55865));
    InMux I__13044 (
            .O(N__55868),
            .I(N__55858));
    LocalMux I__13043 (
            .O(N__55865),
            .I(N__55850));
    InMux I__13042 (
            .O(N__55864),
            .I(N__55847));
    InMux I__13041 (
            .O(N__55863),
            .I(N__55844));
    InMux I__13040 (
            .O(N__55862),
            .I(N__55841));
    InMux I__13039 (
            .O(N__55861),
            .I(N__55838));
    LocalMux I__13038 (
            .O(N__55858),
            .I(N__55835));
    InMux I__13037 (
            .O(N__55857),
            .I(N__55824));
    InMux I__13036 (
            .O(N__55856),
            .I(N__55824));
    InMux I__13035 (
            .O(N__55855),
            .I(N__55824));
    InMux I__13034 (
            .O(N__55854),
            .I(N__55824));
    InMux I__13033 (
            .O(N__55853),
            .I(N__55824));
    Span4Mux_h I__13032 (
            .O(N__55850),
            .I(N__55817));
    LocalMux I__13031 (
            .O(N__55847),
            .I(N__55817));
    LocalMux I__13030 (
            .O(N__55844),
            .I(N__55817));
    LocalMux I__13029 (
            .O(N__55841),
            .I(N__55808));
    LocalMux I__13028 (
            .O(N__55838),
            .I(N__55808));
    Span4Mux_v I__13027 (
            .O(N__55835),
            .I(N__55808));
    LocalMux I__13026 (
            .O(N__55824),
            .I(N__55808));
    Span4Mux_v I__13025 (
            .O(N__55817),
            .I(N__55805));
    Odrv4 I__13024 (
            .O(N__55808),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0 ));
    Odrv4 I__13023 (
            .O(N__55805),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0 ));
    InMux I__13022 (
            .O(N__55800),
            .I(N__55797));
    LocalMux I__13021 (
            .O(N__55797),
            .I(N__55791));
    InMux I__13020 (
            .O(N__55796),
            .I(N__55788));
    InMux I__13019 (
            .O(N__55795),
            .I(N__55785));
    InMux I__13018 (
            .O(N__55794),
            .I(N__55782));
    Span4Mux_v I__13017 (
            .O(N__55791),
            .I(N__55775));
    LocalMux I__13016 (
            .O(N__55788),
            .I(N__55775));
    LocalMux I__13015 (
            .O(N__55785),
            .I(N__55775));
    LocalMux I__13014 (
            .O(N__55782),
            .I(N__55770));
    Span4Mux_h I__13013 (
            .O(N__55775),
            .I(N__55770));
    Odrv4 I__13012 (
            .O(N__55770),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1606_0 ));
    InMux I__13011 (
            .O(N__55767),
            .I(N__55764));
    LocalMux I__13010 (
            .O(N__55764),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1565_0 ));
    InMux I__13009 (
            .O(N__55761),
            .I(N__55758));
    LocalMux I__13008 (
            .O(N__55758),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0 ));
    CascadeMux I__13007 (
            .O(N__55755),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RLZ0Z7_cascade_ ));
    InMux I__13006 (
            .O(N__55752),
            .I(N__55749));
    LocalMux I__13005 (
            .O(N__55749),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2 ));
    InMux I__13004 (
            .O(N__55746),
            .I(N__55735));
    InMux I__13003 (
            .O(N__55745),
            .I(N__55735));
    InMux I__13002 (
            .O(N__55744),
            .I(N__55728));
    InMux I__13001 (
            .O(N__55743),
            .I(N__55728));
    InMux I__13000 (
            .O(N__55742),
            .I(N__55728));
    InMux I__12999 (
            .O(N__55741),
            .I(N__55717));
    InMux I__12998 (
            .O(N__55740),
            .I(N__55717));
    LocalMux I__12997 (
            .O(N__55735),
            .I(N__55712));
    LocalMux I__12996 (
            .O(N__55728),
            .I(N__55712));
    InMux I__12995 (
            .O(N__55727),
            .I(N__55707));
    InMux I__12994 (
            .O(N__55726),
            .I(N__55707));
    InMux I__12993 (
            .O(N__55725),
            .I(N__55702));
    InMux I__12992 (
            .O(N__55724),
            .I(N__55702));
    InMux I__12991 (
            .O(N__55723),
            .I(N__55697));
    InMux I__12990 (
            .O(N__55722),
            .I(N__55697));
    LocalMux I__12989 (
            .O(N__55717),
            .I(N__55690));
    Span4Mux_v I__12988 (
            .O(N__55712),
            .I(N__55683));
    LocalMux I__12987 (
            .O(N__55707),
            .I(N__55680));
    LocalMux I__12986 (
            .O(N__55702),
            .I(N__55675));
    LocalMux I__12985 (
            .O(N__55697),
            .I(N__55675));
    InMux I__12984 (
            .O(N__55696),
            .I(N__55670));
    InMux I__12983 (
            .O(N__55695),
            .I(N__55670));
    InMux I__12982 (
            .O(N__55694),
            .I(N__55665));
    InMux I__12981 (
            .O(N__55693),
            .I(N__55665));
    Span4Mux_h I__12980 (
            .O(N__55690),
            .I(N__55662));
    InMux I__12979 (
            .O(N__55689),
            .I(N__55653));
    InMux I__12978 (
            .O(N__55688),
            .I(N__55653));
    InMux I__12977 (
            .O(N__55687),
            .I(N__55653));
    InMux I__12976 (
            .O(N__55686),
            .I(N__55653));
    Span4Mux_v I__12975 (
            .O(N__55683),
            .I(N__55645));
    Span4Mux_v I__12974 (
            .O(N__55680),
            .I(N__55645));
    Span4Mux_v I__12973 (
            .O(N__55675),
            .I(N__55640));
    LocalMux I__12972 (
            .O(N__55670),
            .I(N__55640));
    LocalMux I__12971 (
            .O(N__55665),
            .I(N__55637));
    Span4Mux_h I__12970 (
            .O(N__55662),
            .I(N__55632));
    LocalMux I__12969 (
            .O(N__55653),
            .I(N__55632));
    InMux I__12968 (
            .O(N__55652),
            .I(N__55625));
    InMux I__12967 (
            .O(N__55651),
            .I(N__55625));
    InMux I__12966 (
            .O(N__55650),
            .I(N__55625));
    Span4Mux_h I__12965 (
            .O(N__55645),
            .I(N__55622));
    Span4Mux_h I__12964 (
            .O(N__55640),
            .I(N__55619));
    Span4Mux_v I__12963 (
            .O(N__55637),
            .I(N__55612));
    Span4Mux_h I__12962 (
            .O(N__55632),
            .I(N__55612));
    LocalMux I__12961 (
            .O(N__55625),
            .I(N__55612));
    Span4Mux_h I__12960 (
            .O(N__55622),
            .I(N__55609));
    Span4Mux_h I__12959 (
            .O(N__55619),
            .I(N__55606));
    Span4Mux_h I__12958 (
            .O(N__55612),
            .I(N__55603));
    Odrv4 I__12957 (
            .O(N__55609),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3 ));
    Odrv4 I__12956 (
            .O(N__55606),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3 ));
    Odrv4 I__12955 (
            .O(N__55603),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3 ));
    CascadeMux I__12954 (
            .O(N__55596),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2_cascade_ ));
    InMux I__12953 (
            .O(N__55593),
            .I(N__55590));
    LocalMux I__12952 (
            .O(N__55590),
            .I(N__55587));
    Odrv4 I__12951 (
            .O(N__55587),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_1 ));
    InMux I__12950 (
            .O(N__55584),
            .I(N__55581));
    LocalMux I__12949 (
            .O(N__55581),
            .I(N__55578));
    Span12Mux_h I__12948 (
            .O(N__55578),
            .I(N__55575));
    Odrv12 I__12947 (
            .O(N__55575),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_2 ));
    CEMux I__12946 (
            .O(N__55572),
            .I(N__55567));
    CEMux I__12945 (
            .O(N__55571),
            .I(N__55564));
    CEMux I__12944 (
            .O(N__55570),
            .I(N__55560));
    LocalMux I__12943 (
            .O(N__55567),
            .I(N__55555));
    LocalMux I__12942 (
            .O(N__55564),
            .I(N__55552));
    CEMux I__12941 (
            .O(N__55563),
            .I(N__55549));
    LocalMux I__12940 (
            .O(N__55560),
            .I(N__55546));
    CEMux I__12939 (
            .O(N__55559),
            .I(N__55543));
    CEMux I__12938 (
            .O(N__55558),
            .I(N__55540));
    Span4Mux_h I__12937 (
            .O(N__55555),
            .I(N__55531));
    Span4Mux_v I__12936 (
            .O(N__55552),
            .I(N__55531));
    LocalMux I__12935 (
            .O(N__55549),
            .I(N__55531));
    Span4Mux_h I__12934 (
            .O(N__55546),
            .I(N__55526));
    LocalMux I__12933 (
            .O(N__55543),
            .I(N__55526));
    LocalMux I__12932 (
            .O(N__55540),
            .I(N__55523));
    CEMux I__12931 (
            .O(N__55539),
            .I(N__55518));
    CEMux I__12930 (
            .O(N__55538),
            .I(N__55515));
    Span4Mux_h I__12929 (
            .O(N__55531),
            .I(N__55512));
    Span4Mux_h I__12928 (
            .O(N__55526),
            .I(N__55507));
    Span4Mux_h I__12927 (
            .O(N__55523),
            .I(N__55507));
    CEMux I__12926 (
            .O(N__55522),
            .I(N__55504));
    CEMux I__12925 (
            .O(N__55521),
            .I(N__55501));
    LocalMux I__12924 (
            .O(N__55518),
            .I(N__55498));
    LocalMux I__12923 (
            .O(N__55515),
            .I(N__55495));
    Span4Mux_h I__12922 (
            .O(N__55512),
            .I(N__55492));
    Span4Mux_h I__12921 (
            .O(N__55507),
            .I(N__55489));
    LocalMux I__12920 (
            .O(N__55504),
            .I(N__55484));
    LocalMux I__12919 (
            .O(N__55501),
            .I(N__55484));
    Span4Mux_v I__12918 (
            .O(N__55498),
            .I(N__55481));
    Span4Mux_v I__12917 (
            .O(N__55495),
            .I(N__55478));
    Sp12to4 I__12916 (
            .O(N__55492),
            .I(N__55475));
    Sp12to4 I__12915 (
            .O(N__55489),
            .I(N__55472));
    Span4Mux_v I__12914 (
            .O(N__55484),
            .I(N__55467));
    Span4Mux_h I__12913 (
            .O(N__55481),
            .I(N__55467));
    Sp12to4 I__12912 (
            .O(N__55478),
            .I(N__55460));
    Span12Mux_v I__12911 (
            .O(N__55475),
            .I(N__55460));
    Span12Mux_v I__12910 (
            .O(N__55472),
            .I(N__55460));
    Odrv4 I__12909 (
            .O(N__55467),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i ));
    Odrv12 I__12908 (
            .O(N__55460),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i ));
    InMux I__12907 (
            .O(N__55455),
            .I(N__55439));
    InMux I__12906 (
            .O(N__55454),
            .I(N__55439));
    InMux I__12905 (
            .O(N__55453),
            .I(N__55435));
    InMux I__12904 (
            .O(N__55452),
            .I(N__55432));
    CascadeMux I__12903 (
            .O(N__55451),
            .I(N__55424));
    InMux I__12902 (
            .O(N__55450),
            .I(N__55420));
    InMux I__12901 (
            .O(N__55449),
            .I(N__55417));
    InMux I__12900 (
            .O(N__55448),
            .I(N__55410));
    InMux I__12899 (
            .O(N__55447),
            .I(N__55410));
    InMux I__12898 (
            .O(N__55446),
            .I(N__55410));
    InMux I__12897 (
            .O(N__55445),
            .I(N__55406));
    InMux I__12896 (
            .O(N__55444),
            .I(N__55403));
    LocalMux I__12895 (
            .O(N__55439),
            .I(N__55400));
    InMux I__12894 (
            .O(N__55438),
            .I(N__55396));
    LocalMux I__12893 (
            .O(N__55435),
            .I(N__55391));
    LocalMux I__12892 (
            .O(N__55432),
            .I(N__55391));
    InMux I__12891 (
            .O(N__55431),
            .I(N__55388));
    InMux I__12890 (
            .O(N__55430),
            .I(N__55383));
    InMux I__12889 (
            .O(N__55429),
            .I(N__55376));
    InMux I__12888 (
            .O(N__55428),
            .I(N__55376));
    InMux I__12887 (
            .O(N__55427),
            .I(N__55376));
    InMux I__12886 (
            .O(N__55424),
            .I(N__55373));
    InMux I__12885 (
            .O(N__55423),
            .I(N__55370));
    LocalMux I__12884 (
            .O(N__55420),
            .I(N__55367));
    LocalMux I__12883 (
            .O(N__55417),
            .I(N__55362));
    LocalMux I__12882 (
            .O(N__55410),
            .I(N__55362));
    InMux I__12881 (
            .O(N__55409),
            .I(N__55359));
    LocalMux I__12880 (
            .O(N__55406),
            .I(N__55352));
    LocalMux I__12879 (
            .O(N__55403),
            .I(N__55352));
    Span4Mux_h I__12878 (
            .O(N__55400),
            .I(N__55352));
    InMux I__12877 (
            .O(N__55399),
            .I(N__55348));
    LocalMux I__12876 (
            .O(N__55396),
            .I(N__55345));
    Span4Mux_v I__12875 (
            .O(N__55391),
            .I(N__55342));
    LocalMux I__12874 (
            .O(N__55388),
            .I(N__55339));
    InMux I__12873 (
            .O(N__55387),
            .I(N__55336));
    InMux I__12872 (
            .O(N__55386),
            .I(N__55333));
    LocalMux I__12871 (
            .O(N__55383),
            .I(N__55328));
    LocalMux I__12870 (
            .O(N__55376),
            .I(N__55328));
    LocalMux I__12869 (
            .O(N__55373),
            .I(N__55319));
    LocalMux I__12868 (
            .O(N__55370),
            .I(N__55319));
    Span4Mux_h I__12867 (
            .O(N__55367),
            .I(N__55319));
    Span4Mux_h I__12866 (
            .O(N__55362),
            .I(N__55319));
    LocalMux I__12865 (
            .O(N__55359),
            .I(N__55314));
    Span4Mux_v I__12864 (
            .O(N__55352),
            .I(N__55314));
    InMux I__12863 (
            .O(N__55351),
            .I(N__55311));
    LocalMux I__12862 (
            .O(N__55348),
            .I(N__55306));
    Span4Mux_h I__12861 (
            .O(N__55345),
            .I(N__55306));
    Span4Mux_h I__12860 (
            .O(N__55342),
            .I(N__55303));
    Span4Mux_v I__12859 (
            .O(N__55339),
            .I(N__55296));
    LocalMux I__12858 (
            .O(N__55336),
            .I(N__55296));
    LocalMux I__12857 (
            .O(N__55333),
            .I(N__55296));
    Span4Mux_h I__12856 (
            .O(N__55328),
            .I(N__55291));
    Span4Mux_v I__12855 (
            .O(N__55319),
            .I(N__55291));
    Span4Mux_h I__12854 (
            .O(N__55314),
            .I(N__55288));
    LocalMux I__12853 (
            .O(N__55311),
            .I(N__55283));
    Span4Mux_v I__12852 (
            .O(N__55306),
            .I(N__55283));
    Span4Mux_h I__12851 (
            .O(N__55303),
            .I(N__55278));
    Span4Mux_v I__12850 (
            .O(N__55296),
            .I(N__55278));
    Span4Mux_h I__12849 (
            .O(N__55291),
            .I(N__55275));
    Span4Mux_v I__12848 (
            .O(N__55288),
            .I(N__55272));
    Odrv4 I__12847 (
            .O(N__55283),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270 ));
    Odrv4 I__12846 (
            .O(N__55278),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270 ));
    Odrv4 I__12845 (
            .O(N__55275),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270 ));
    Odrv4 I__12844 (
            .O(N__55272),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270 ));
    InMux I__12843 (
            .O(N__55263),
            .I(N__55259));
    InMux I__12842 (
            .O(N__55262),
            .I(N__55251));
    LocalMux I__12841 (
            .O(N__55259),
            .I(N__55246));
    InMux I__12840 (
            .O(N__55258),
            .I(N__55239));
    InMux I__12839 (
            .O(N__55257),
            .I(N__55239));
    InMux I__12838 (
            .O(N__55256),
            .I(N__55239));
    InMux I__12837 (
            .O(N__55255),
            .I(N__55236));
    InMux I__12836 (
            .O(N__55254),
            .I(N__55233));
    LocalMux I__12835 (
            .O(N__55251),
            .I(N__55225));
    InMux I__12834 (
            .O(N__55250),
            .I(N__55222));
    InMux I__12833 (
            .O(N__55249),
            .I(N__55218));
    Span4Mux_h I__12832 (
            .O(N__55246),
            .I(N__55212));
    LocalMux I__12831 (
            .O(N__55239),
            .I(N__55212));
    LocalMux I__12830 (
            .O(N__55236),
            .I(N__55209));
    LocalMux I__12829 (
            .O(N__55233),
            .I(N__55206));
    InMux I__12828 (
            .O(N__55232),
            .I(N__55199));
    InMux I__12827 (
            .O(N__55231),
            .I(N__55199));
    InMux I__12826 (
            .O(N__55230),
            .I(N__55199));
    InMux I__12825 (
            .O(N__55229),
            .I(N__55193));
    InMux I__12824 (
            .O(N__55228),
            .I(N__55193));
    Span4Mux_v I__12823 (
            .O(N__55225),
            .I(N__55187));
    LocalMux I__12822 (
            .O(N__55222),
            .I(N__55187));
    InMux I__12821 (
            .O(N__55221),
            .I(N__55184));
    LocalMux I__12820 (
            .O(N__55218),
            .I(N__55180));
    InMux I__12819 (
            .O(N__55217),
            .I(N__55177));
    Span4Mux_h I__12818 (
            .O(N__55212),
            .I(N__55174));
    Span4Mux_h I__12817 (
            .O(N__55209),
            .I(N__55167));
    Span4Mux_v I__12816 (
            .O(N__55206),
            .I(N__55167));
    LocalMux I__12815 (
            .O(N__55199),
            .I(N__55167));
    InMux I__12814 (
            .O(N__55198),
            .I(N__55164));
    LocalMux I__12813 (
            .O(N__55193),
            .I(N__55160));
    CascadeMux I__12812 (
            .O(N__55192),
            .I(N__55157));
    Span4Mux_h I__12811 (
            .O(N__55187),
            .I(N__55151));
    LocalMux I__12810 (
            .O(N__55184),
            .I(N__55148));
    InMux I__12809 (
            .O(N__55183),
            .I(N__55145));
    Span4Mux_h I__12808 (
            .O(N__55180),
            .I(N__55140));
    LocalMux I__12807 (
            .O(N__55177),
            .I(N__55140));
    Span4Mux_v I__12806 (
            .O(N__55174),
            .I(N__55135));
    Span4Mux_h I__12805 (
            .O(N__55167),
            .I(N__55135));
    LocalMux I__12804 (
            .O(N__55164),
            .I(N__55132));
    InMux I__12803 (
            .O(N__55163),
            .I(N__55129));
    Span4Mux_v I__12802 (
            .O(N__55160),
            .I(N__55126));
    InMux I__12801 (
            .O(N__55157),
            .I(N__55123));
    InMux I__12800 (
            .O(N__55156),
            .I(N__55120));
    InMux I__12799 (
            .O(N__55155),
            .I(N__55117));
    InMux I__12798 (
            .O(N__55154),
            .I(N__55114));
    Span4Mux_h I__12797 (
            .O(N__55151),
            .I(N__55110));
    Span4Mux_h I__12796 (
            .O(N__55148),
            .I(N__55105));
    LocalMux I__12795 (
            .O(N__55145),
            .I(N__55105));
    Span4Mux_h I__12794 (
            .O(N__55140),
            .I(N__55098));
    Span4Mux_h I__12793 (
            .O(N__55135),
            .I(N__55098));
    Span4Mux_v I__12792 (
            .O(N__55132),
            .I(N__55098));
    LocalMux I__12791 (
            .O(N__55129),
            .I(N__55085));
    Sp12to4 I__12790 (
            .O(N__55126),
            .I(N__55085));
    LocalMux I__12789 (
            .O(N__55123),
            .I(N__55085));
    LocalMux I__12788 (
            .O(N__55120),
            .I(N__55085));
    LocalMux I__12787 (
            .O(N__55117),
            .I(N__55085));
    LocalMux I__12786 (
            .O(N__55114),
            .I(N__55085));
    InMux I__12785 (
            .O(N__55113),
            .I(N__55082));
    Span4Mux_v I__12784 (
            .O(N__55110),
            .I(N__55079));
    Span4Mux_v I__12783 (
            .O(N__55105),
            .I(N__55076));
    Sp12to4 I__12782 (
            .O(N__55098),
            .I(N__55069));
    Span12Mux_h I__12781 (
            .O(N__55085),
            .I(N__55069));
    LocalMux I__12780 (
            .O(N__55082),
            .I(N__55069));
    Odrv4 I__12779 (
            .O(N__55079),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274 ));
    Odrv4 I__12778 (
            .O(N__55076),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274 ));
    Odrv12 I__12777 (
            .O(N__55069),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274 ));
    CascadeMux I__12776 (
            .O(N__55062),
            .I(N__55059));
    InMux I__12775 (
            .O(N__55059),
            .I(N__55049));
    InMux I__12774 (
            .O(N__55058),
            .I(N__55046));
    InMux I__12773 (
            .O(N__55057),
            .I(N__55043));
    InMux I__12772 (
            .O(N__55056),
            .I(N__55040));
    InMux I__12771 (
            .O(N__55055),
            .I(N__55037));
    InMux I__12770 (
            .O(N__55054),
            .I(N__55032));
    CascadeMux I__12769 (
            .O(N__55053),
            .I(N__55026));
    CascadeMux I__12768 (
            .O(N__55052),
            .I(N__55023));
    LocalMux I__12767 (
            .O(N__55049),
            .I(N__55014));
    LocalMux I__12766 (
            .O(N__55046),
            .I(N__55014));
    LocalMux I__12765 (
            .O(N__55043),
            .I(N__55011));
    LocalMux I__12764 (
            .O(N__55040),
            .I(N__55005));
    LocalMux I__12763 (
            .O(N__55037),
            .I(N__55005));
    InMux I__12762 (
            .O(N__55036),
            .I(N__55002));
    CascadeMux I__12761 (
            .O(N__55035),
            .I(N__54998));
    LocalMux I__12760 (
            .O(N__55032),
            .I(N__54995));
    InMux I__12759 (
            .O(N__55031),
            .I(N__54992));
    InMux I__12758 (
            .O(N__55030),
            .I(N__54989));
    InMux I__12757 (
            .O(N__55029),
            .I(N__54986));
    InMux I__12756 (
            .O(N__55026),
            .I(N__54979));
    InMux I__12755 (
            .O(N__55023),
            .I(N__54979));
    InMux I__12754 (
            .O(N__55022),
            .I(N__54979));
    InMux I__12753 (
            .O(N__55021),
            .I(N__54976));
    InMux I__12752 (
            .O(N__55020),
            .I(N__54973));
    CascadeMux I__12751 (
            .O(N__55019),
            .I(N__54970));
    Span4Mux_v I__12750 (
            .O(N__55014),
            .I(N__54967));
    Span4Mux_v I__12749 (
            .O(N__55011),
            .I(N__54964));
    InMux I__12748 (
            .O(N__55010),
            .I(N__54960));
    Span4Mux_v I__12747 (
            .O(N__55005),
            .I(N__54955));
    LocalMux I__12746 (
            .O(N__55002),
            .I(N__54955));
    InMux I__12745 (
            .O(N__55001),
            .I(N__54950));
    InMux I__12744 (
            .O(N__54998),
            .I(N__54947));
    Span4Mux_v I__12743 (
            .O(N__54995),
            .I(N__54944));
    LocalMux I__12742 (
            .O(N__54992),
            .I(N__54939));
    LocalMux I__12741 (
            .O(N__54989),
            .I(N__54939));
    LocalMux I__12740 (
            .O(N__54986),
            .I(N__54930));
    LocalMux I__12739 (
            .O(N__54979),
            .I(N__54930));
    LocalMux I__12738 (
            .O(N__54976),
            .I(N__54930));
    LocalMux I__12737 (
            .O(N__54973),
            .I(N__54930));
    InMux I__12736 (
            .O(N__54970),
            .I(N__54925));
    Span4Mux_v I__12735 (
            .O(N__54967),
            .I(N__54920));
    Span4Mux_v I__12734 (
            .O(N__54964),
            .I(N__54920));
    InMux I__12733 (
            .O(N__54963),
            .I(N__54917));
    LocalMux I__12732 (
            .O(N__54960),
            .I(N__54914));
    Span4Mux_v I__12731 (
            .O(N__54955),
            .I(N__54911));
    InMux I__12730 (
            .O(N__54954),
            .I(N__54908));
    InMux I__12729 (
            .O(N__54953),
            .I(N__54905));
    LocalMux I__12728 (
            .O(N__54950),
            .I(N__54902));
    LocalMux I__12727 (
            .O(N__54947),
            .I(N__54893));
    Span4Mux_h I__12726 (
            .O(N__54944),
            .I(N__54893));
    Span4Mux_v I__12725 (
            .O(N__54939),
            .I(N__54893));
    Span4Mux_v I__12724 (
            .O(N__54930),
            .I(N__54893));
    InMux I__12723 (
            .O(N__54929),
            .I(N__54888));
    InMux I__12722 (
            .O(N__54928),
            .I(N__54888));
    LocalMux I__12721 (
            .O(N__54925),
            .I(N__54885));
    Span4Mux_h I__12720 (
            .O(N__54920),
            .I(N__54882));
    LocalMux I__12719 (
            .O(N__54917),
            .I(N__54879));
    Span4Mux_v I__12718 (
            .O(N__54914),
            .I(N__54874));
    Span4Mux_h I__12717 (
            .O(N__54911),
            .I(N__54874));
    LocalMux I__12716 (
            .O(N__54908),
            .I(N__54871));
    LocalMux I__12715 (
            .O(N__54905),
            .I(N__54862));
    Span4Mux_v I__12714 (
            .O(N__54902),
            .I(N__54862));
    Span4Mux_h I__12713 (
            .O(N__54893),
            .I(N__54862));
    LocalMux I__12712 (
            .O(N__54888),
            .I(N__54862));
    Span12Mux_h I__12711 (
            .O(N__54885),
            .I(N__54859));
    Sp12to4 I__12710 (
            .O(N__54882),
            .I(N__54854));
    Span12Mux_v I__12709 (
            .O(N__54879),
            .I(N__54854));
    Span4Mux_h I__12708 (
            .O(N__54874),
            .I(N__54851));
    Span4Mux_v I__12707 (
            .O(N__54871),
            .I(N__54846));
    Span4Mux_h I__12706 (
            .O(N__54862),
            .I(N__54846));
    Odrv12 I__12705 (
            .O(N__54859),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0 ));
    Odrv12 I__12704 (
            .O(N__54854),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0 ));
    Odrv4 I__12703 (
            .O(N__54851),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0 ));
    Odrv4 I__12702 (
            .O(N__54846),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0 ));
    InMux I__12701 (
            .O(N__54837),
            .I(N__54829));
    CascadeMux I__12700 (
            .O(N__54836),
            .I(N__54826));
    CascadeMux I__12699 (
            .O(N__54835),
            .I(N__54822));
    InMux I__12698 (
            .O(N__54834),
            .I(N__54813));
    InMux I__12697 (
            .O(N__54833),
            .I(N__54810));
    InMux I__12696 (
            .O(N__54832),
            .I(N__54807));
    LocalMux I__12695 (
            .O(N__54829),
            .I(N__54803));
    InMux I__12694 (
            .O(N__54826),
            .I(N__54799));
    InMux I__12693 (
            .O(N__54825),
            .I(N__54795));
    InMux I__12692 (
            .O(N__54822),
            .I(N__54792));
    InMux I__12691 (
            .O(N__54821),
            .I(N__54789));
    InMux I__12690 (
            .O(N__54820),
            .I(N__54784));
    InMux I__12689 (
            .O(N__54819),
            .I(N__54784));
    InMux I__12688 (
            .O(N__54818),
            .I(N__54775));
    InMux I__12687 (
            .O(N__54817),
            .I(N__54775));
    InMux I__12686 (
            .O(N__54816),
            .I(N__54772));
    LocalMux I__12685 (
            .O(N__54813),
            .I(N__54769));
    LocalMux I__12684 (
            .O(N__54810),
            .I(N__54764));
    LocalMux I__12683 (
            .O(N__54807),
            .I(N__54764));
    InMux I__12682 (
            .O(N__54806),
            .I(N__54761));
    Span4Mux_h I__12681 (
            .O(N__54803),
            .I(N__54758));
    InMux I__12680 (
            .O(N__54802),
            .I(N__54753));
    LocalMux I__12679 (
            .O(N__54799),
            .I(N__54750));
    InMux I__12678 (
            .O(N__54798),
            .I(N__54747));
    LocalMux I__12677 (
            .O(N__54795),
            .I(N__54744));
    LocalMux I__12676 (
            .O(N__54792),
            .I(N__54737));
    LocalMux I__12675 (
            .O(N__54789),
            .I(N__54737));
    LocalMux I__12674 (
            .O(N__54784),
            .I(N__54737));
    InMux I__12673 (
            .O(N__54783),
            .I(N__54732));
    InMux I__12672 (
            .O(N__54782),
            .I(N__54729));
    InMux I__12671 (
            .O(N__54781),
            .I(N__54724));
    InMux I__12670 (
            .O(N__54780),
            .I(N__54724));
    LocalMux I__12669 (
            .O(N__54775),
            .I(N__54721));
    LocalMux I__12668 (
            .O(N__54772),
            .I(N__54712));
    Span4Mux_v I__12667 (
            .O(N__54769),
            .I(N__54712));
    Span4Mux_h I__12666 (
            .O(N__54764),
            .I(N__54712));
    LocalMux I__12665 (
            .O(N__54761),
            .I(N__54712));
    Span4Mux_v I__12664 (
            .O(N__54758),
            .I(N__54709));
    InMux I__12663 (
            .O(N__54757),
            .I(N__54706));
    InMux I__12662 (
            .O(N__54756),
            .I(N__54703));
    LocalMux I__12661 (
            .O(N__54753),
            .I(N__54698));
    Span4Mux_v I__12660 (
            .O(N__54750),
            .I(N__54698));
    LocalMux I__12659 (
            .O(N__54747),
            .I(N__54691));
    Span4Mux_h I__12658 (
            .O(N__54744),
            .I(N__54691));
    Span4Mux_v I__12657 (
            .O(N__54737),
            .I(N__54691));
    InMux I__12656 (
            .O(N__54736),
            .I(N__54686));
    InMux I__12655 (
            .O(N__54735),
            .I(N__54686));
    LocalMux I__12654 (
            .O(N__54732),
            .I(N__54675));
    LocalMux I__12653 (
            .O(N__54729),
            .I(N__54675));
    LocalMux I__12652 (
            .O(N__54724),
            .I(N__54675));
    Span4Mux_v I__12651 (
            .O(N__54721),
            .I(N__54675));
    Span4Mux_v I__12650 (
            .O(N__54712),
            .I(N__54675));
    Span4Mux_h I__12649 (
            .O(N__54709),
            .I(N__54672));
    LocalMux I__12648 (
            .O(N__54706),
            .I(N__54669));
    LocalMux I__12647 (
            .O(N__54703),
            .I(N__54660));
    Span4Mux_h I__12646 (
            .O(N__54698),
            .I(N__54660));
    Span4Mux_h I__12645 (
            .O(N__54691),
            .I(N__54660));
    LocalMux I__12644 (
            .O(N__54686),
            .I(N__54660));
    Span4Mux_h I__12643 (
            .O(N__54675),
            .I(N__54657));
    Span4Mux_h I__12642 (
            .O(N__54672),
            .I(N__54654));
    Span4Mux_v I__12641 (
            .O(N__54669),
            .I(N__54649));
    Span4Mux_h I__12640 (
            .O(N__54660),
            .I(N__54649));
    Span4Mux_h I__12639 (
            .O(N__54657),
            .I(N__54646));
    Odrv4 I__12638 (
            .O(N__54654),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270 ));
    Odrv4 I__12637 (
            .O(N__54649),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270 ));
    Odrv4 I__12636 (
            .O(N__54646),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270 ));
    InMux I__12635 (
            .O(N__54639),
            .I(N__54635));
    CascadeMux I__12634 (
            .O(N__54638),
            .I(N__54631));
    LocalMux I__12633 (
            .O(N__54635),
            .I(N__54628));
    InMux I__12632 (
            .O(N__54634),
            .I(N__54623));
    InMux I__12631 (
            .O(N__54631),
            .I(N__54623));
    Span4Mux_h I__12630 (
            .O(N__54628),
            .I(N__54620));
    LocalMux I__12629 (
            .O(N__54623),
            .I(N__54617));
    Span4Mux_v I__12628 (
            .O(N__54620),
            .I(N__54614));
    Span4Mux_v I__12627 (
            .O(N__54617),
            .I(N__54611));
    Span4Mux_h I__12626 (
            .O(N__54614),
            .I(N__54606));
    Span4Mux_h I__12625 (
            .O(N__54611),
            .I(N__54606));
    Odrv4 I__12624 (
            .O(N__54606),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_1));
    InMux I__12623 (
            .O(N__54603),
            .I(N__54600));
    LocalMux I__12622 (
            .O(N__54600),
            .I(N__54595));
    InMux I__12621 (
            .O(N__54599),
            .I(N__54592));
    InMux I__12620 (
            .O(N__54598),
            .I(N__54589));
    Span12Mux_h I__12619 (
            .O(N__54595),
            .I(N__54586));
    LocalMux I__12618 (
            .O(N__54592),
            .I(N__54581));
    LocalMux I__12617 (
            .O(N__54589),
            .I(N__54581));
    Odrv12 I__12616 (
            .O(N__54586),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_1));
    Odrv12 I__12615 (
            .O(N__54581),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_1));
    InMux I__12614 (
            .O(N__54576),
            .I(N__54573));
    LocalMux I__12613 (
            .O(N__54573),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_1 ));
    InMux I__12612 (
            .O(N__54570),
            .I(N__54567));
    LocalMux I__12611 (
            .O(N__54567),
            .I(N__54564));
    Span12Mux_h I__12610 (
            .O(N__54564),
            .I(N__54561));
    Odrv12 I__12609 (
            .O(N__54561),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_3_26 ));
    InMux I__12608 (
            .O(N__54558),
            .I(N__54555));
    LocalMux I__12607 (
            .O(N__54555),
            .I(N__54552));
    Span12Mux_v I__12606 (
            .O(N__54552),
            .I(N__54549));
    Odrv12 I__12605 (
            .O(N__54549),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_4093_0 ));
    CascadeMux I__12604 (
            .O(N__54546),
            .I(N__54543));
    InMux I__12603 (
            .O(N__54543),
            .I(N__54540));
    LocalMux I__12602 (
            .O(N__54540),
            .I(N__54537));
    Span4Mux_h I__12601 (
            .O(N__54537),
            .I(N__54534));
    Span4Mux_h I__12600 (
            .O(N__54534),
            .I(N__54531));
    Span4Mux_h I__12599 (
            .O(N__54531),
            .I(N__54528));
    Odrv4 I__12598 (
            .O(N__54528),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_26 ));
    CEMux I__12597 (
            .O(N__54525),
            .I(N__54429));
    CEMux I__12596 (
            .O(N__54524),
            .I(N__54429));
    CEMux I__12595 (
            .O(N__54523),
            .I(N__54429));
    CEMux I__12594 (
            .O(N__54522),
            .I(N__54429));
    CEMux I__12593 (
            .O(N__54521),
            .I(N__54429));
    CEMux I__12592 (
            .O(N__54520),
            .I(N__54429));
    CEMux I__12591 (
            .O(N__54519),
            .I(N__54429));
    CEMux I__12590 (
            .O(N__54518),
            .I(N__54429));
    CEMux I__12589 (
            .O(N__54517),
            .I(N__54429));
    CEMux I__12588 (
            .O(N__54516),
            .I(N__54429));
    CEMux I__12587 (
            .O(N__54515),
            .I(N__54429));
    CEMux I__12586 (
            .O(N__54514),
            .I(N__54429));
    CEMux I__12585 (
            .O(N__54513),
            .I(N__54429));
    CEMux I__12584 (
            .O(N__54512),
            .I(N__54429));
    CEMux I__12583 (
            .O(N__54511),
            .I(N__54429));
    CEMux I__12582 (
            .O(N__54510),
            .I(N__54429));
    CEMux I__12581 (
            .O(N__54509),
            .I(N__54429));
    CEMux I__12580 (
            .O(N__54508),
            .I(N__54429));
    CEMux I__12579 (
            .O(N__54507),
            .I(N__54429));
    CEMux I__12578 (
            .O(N__54506),
            .I(N__54429));
    CEMux I__12577 (
            .O(N__54505),
            .I(N__54429));
    CEMux I__12576 (
            .O(N__54504),
            .I(N__54429));
    CEMux I__12575 (
            .O(N__54503),
            .I(N__54429));
    CEMux I__12574 (
            .O(N__54502),
            .I(N__54429));
    CEMux I__12573 (
            .O(N__54501),
            .I(N__54429));
    CEMux I__12572 (
            .O(N__54500),
            .I(N__54429));
    CEMux I__12571 (
            .O(N__54499),
            .I(N__54429));
    CEMux I__12570 (
            .O(N__54498),
            .I(N__54429));
    CEMux I__12569 (
            .O(N__54497),
            .I(N__54429));
    CEMux I__12568 (
            .O(N__54496),
            .I(N__54429));
    CEMux I__12567 (
            .O(N__54495),
            .I(N__54429));
    CEMux I__12566 (
            .O(N__54494),
            .I(N__54429));
    GlobalMux I__12565 (
            .O(N__54429),
            .I(N__54426));
    gio2CtrlBuf I__12564 (
            .O(N__54426),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_g ));
    InMux I__12563 (
            .O(N__54423),
            .I(N__54420));
    LocalMux I__12562 (
            .O(N__54420),
            .I(N__54416));
    InMux I__12561 (
            .O(N__54419),
            .I(N__54413));
    Span4Mux_v I__12560 (
            .O(N__54416),
            .I(N__54410));
    LocalMux I__12559 (
            .O(N__54413),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i ));
    Odrv4 I__12558 (
            .O(N__54410),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i ));
    CascadeMux I__12557 (
            .O(N__54405),
            .I(N__54399));
    InMux I__12556 (
            .O(N__54404),
            .I(N__54395));
    InMux I__12555 (
            .O(N__54403),
            .I(N__54392));
    InMux I__12554 (
            .O(N__54402),
            .I(N__54389));
    InMux I__12553 (
            .O(N__54399),
            .I(N__54384));
    InMux I__12552 (
            .O(N__54398),
            .I(N__54384));
    LocalMux I__12551 (
            .O(N__54395),
            .I(N__54381));
    LocalMux I__12550 (
            .O(N__54392),
            .I(N__54373));
    LocalMux I__12549 (
            .O(N__54389),
            .I(N__54373));
    LocalMux I__12548 (
            .O(N__54384),
            .I(N__54373));
    Span4Mux_v I__12547 (
            .O(N__54381),
            .I(N__54370));
    InMux I__12546 (
            .O(N__54380),
            .I(N__54367));
    Span4Mux_h I__12545 (
            .O(N__54373),
            .I(N__54364));
    Sp12to4 I__12544 (
            .O(N__54370),
            .I(N__54359));
    LocalMux I__12543 (
            .O(N__54367),
            .I(N__54359));
    Span4Mux_h I__12542 (
            .O(N__54364),
            .I(N__54356));
    Odrv12 I__12541 (
            .O(N__54359),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0 ));
    Odrv4 I__12540 (
            .O(N__54356),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0 ));
    CascadeMux I__12539 (
            .O(N__54351),
            .I(N__54348));
    InMux I__12538 (
            .O(N__54348),
            .I(N__54345));
    LocalMux I__12537 (
            .O(N__54345),
            .I(N__54339));
    InMux I__12536 (
            .O(N__54344),
            .I(N__54331));
    InMux I__12535 (
            .O(N__54343),
            .I(N__54326));
    InMux I__12534 (
            .O(N__54342),
            .I(N__54326));
    Span4Mux_v I__12533 (
            .O(N__54339),
            .I(N__54323));
    InMux I__12532 (
            .O(N__54338),
            .I(N__54320));
    InMux I__12531 (
            .O(N__54337),
            .I(N__54315));
    InMux I__12530 (
            .O(N__54336),
            .I(N__54315));
    InMux I__12529 (
            .O(N__54335),
            .I(N__54312));
    InMux I__12528 (
            .O(N__54334),
            .I(N__54309));
    LocalMux I__12527 (
            .O(N__54331),
            .I(N__54306));
    LocalMux I__12526 (
            .O(N__54326),
            .I(N__54303));
    Span4Mux_h I__12525 (
            .O(N__54323),
            .I(N__54300));
    LocalMux I__12524 (
            .O(N__54320),
            .I(N__54293));
    LocalMux I__12523 (
            .O(N__54315),
            .I(N__54293));
    LocalMux I__12522 (
            .O(N__54312),
            .I(N__54293));
    LocalMux I__12521 (
            .O(N__54309),
            .I(N__54290));
    Span12Mux_v I__12520 (
            .O(N__54306),
            .I(N__54285));
    Span4Mux_v I__12519 (
            .O(N__54303),
            .I(N__54282));
    Span4Mux_h I__12518 (
            .O(N__54300),
            .I(N__54277));
    Span4Mux_v I__12517 (
            .O(N__54293),
            .I(N__54277));
    Span4Mux_h I__12516 (
            .O(N__54290),
            .I(N__54274));
    InMux I__12515 (
            .O(N__54289),
            .I(N__54269));
    InMux I__12514 (
            .O(N__54288),
            .I(N__54269));
    Odrv12 I__12513 (
            .O(N__54285),
            .I(s_paddr_I2C_3));
    Odrv4 I__12512 (
            .O(N__54282),
            .I(s_paddr_I2C_3));
    Odrv4 I__12511 (
            .O(N__54277),
            .I(s_paddr_I2C_3));
    Odrv4 I__12510 (
            .O(N__54274),
            .I(s_paddr_I2C_3));
    LocalMux I__12509 (
            .O(N__54269),
            .I(s_paddr_I2C_3));
    InMux I__12508 (
            .O(N__54258),
            .I(N__54255));
    LocalMux I__12507 (
            .O(N__54255),
            .I(N__54252));
    Span4Mux_v I__12506 (
            .O(N__54252),
            .I(N__54248));
    InMux I__12505 (
            .O(N__54251),
            .I(N__54245));
    Odrv4 I__12504 (
            .O(N__54248),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0 ));
    LocalMux I__12503 (
            .O(N__54245),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0 ));
    CascadeMux I__12502 (
            .O(N__54240),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_230_cascade_ ));
    InMux I__12501 (
            .O(N__54237),
            .I(N__54234));
    LocalMux I__12500 (
            .O(N__54234),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_0_sqmuxa ));
    CascadeMux I__12499 (
            .O(N__54231),
            .I(N__54228));
    InMux I__12498 (
            .O(N__54228),
            .I(N__54225));
    LocalMux I__12497 (
            .O(N__54225),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_2_sqmuxa ));
    InMux I__12496 (
            .O(N__54222),
            .I(N__54219));
    LocalMux I__12495 (
            .O(N__54219),
            .I(N__54216));
    Span4Mux_v I__12494 (
            .O(N__54216),
            .I(N__54213));
    Span4Mux_h I__12493 (
            .O(N__54213),
            .I(N__54210));
    Odrv4 I__12492 (
            .O(N__54210),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_24));
    InMux I__12491 (
            .O(N__54207),
            .I(N__54203));
    InMux I__12490 (
            .O(N__54206),
            .I(N__54200));
    LocalMux I__12489 (
            .O(N__54203),
            .I(N__54197));
    LocalMux I__12488 (
            .O(N__54200),
            .I(N__54194));
    Span4Mux_h I__12487 (
            .O(N__54197),
            .I(N__54190));
    Span4Mux_h I__12486 (
            .O(N__54194),
            .I(N__54187));
    InMux I__12485 (
            .O(N__54193),
            .I(N__54184));
    Odrv4 I__12484 (
            .O(N__54190),
            .I(cemf_module_64ch_ctrl_inst1_data_config_16));
    Odrv4 I__12483 (
            .O(N__54187),
            .I(cemf_module_64ch_ctrl_inst1_data_config_16));
    LocalMux I__12482 (
            .O(N__54184),
            .I(cemf_module_64ch_ctrl_inst1_data_config_16));
    InMux I__12481 (
            .O(N__54177),
            .I(N__54174));
    LocalMux I__12480 (
            .O(N__54174),
            .I(N__54171));
    Span12Mux_v I__12479 (
            .O(N__54171),
            .I(N__54168));
    Odrv12 I__12478 (
            .O(N__54168),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_28));
    CascadeMux I__12477 (
            .O(N__54165),
            .I(N__54162));
    InMux I__12476 (
            .O(N__54162),
            .I(N__54159));
    LocalMux I__12475 (
            .O(N__54159),
            .I(N__54156));
    Span4Mux_v I__12474 (
            .O(N__54156),
            .I(N__54153));
    Span4Mux_h I__12473 (
            .O(N__54153),
            .I(N__54149));
    InMux I__12472 (
            .O(N__54152),
            .I(N__54146));
    Span4Mux_h I__12471 (
            .O(N__54149),
            .I(N__54143));
    LocalMux I__12470 (
            .O(N__54146),
            .I(N__54139));
    Span4Mux_h I__12469 (
            .O(N__54143),
            .I(N__54136));
    InMux I__12468 (
            .O(N__54142),
            .I(N__54133));
    Span4Mux_h I__12467 (
            .O(N__54139),
            .I(N__54130));
    Odrv4 I__12466 (
            .O(N__54136),
            .I(cemf_module_64ch_ctrl_inst1_data_config_17));
    LocalMux I__12465 (
            .O(N__54133),
            .I(cemf_module_64ch_ctrl_inst1_data_config_17));
    Odrv4 I__12464 (
            .O(N__54130),
            .I(cemf_module_64ch_ctrl_inst1_data_config_17));
    CEMux I__12463 (
            .O(N__54123),
            .I(N__54120));
    LocalMux I__12462 (
            .O(N__54120),
            .I(N__54115));
    CEMux I__12461 (
            .O(N__54119),
            .I(N__54109));
    CEMux I__12460 (
            .O(N__54118),
            .I(N__54106));
    Span4Mux_h I__12459 (
            .O(N__54115),
            .I(N__54103));
    CEMux I__12458 (
            .O(N__54114),
            .I(N__54100));
    CEMux I__12457 (
            .O(N__54113),
            .I(N__54097));
    CEMux I__12456 (
            .O(N__54112),
            .I(N__54094));
    LocalMux I__12455 (
            .O(N__54109),
            .I(N__54091));
    LocalMux I__12454 (
            .O(N__54106),
            .I(N__54086));
    Span4Mux_v I__12453 (
            .O(N__54103),
            .I(N__54086));
    LocalMux I__12452 (
            .O(N__54100),
            .I(N__54083));
    LocalMux I__12451 (
            .O(N__54097),
            .I(N__54080));
    LocalMux I__12450 (
            .O(N__54094),
            .I(N__54077));
    Span4Mux_h I__12449 (
            .O(N__54091),
            .I(N__54074));
    Span4Mux_h I__12448 (
            .O(N__54086),
            .I(N__54071));
    Span12Mux_h I__12447 (
            .O(N__54083),
            .I(N__54068));
    Span4Mux_h I__12446 (
            .O(N__54080),
            .I(N__54065));
    Span4Mux_h I__12445 (
            .O(N__54077),
            .I(N__54060));
    Span4Mux_h I__12444 (
            .O(N__54074),
            .I(N__54060));
    Span4Mux_h I__12443 (
            .O(N__54071),
            .I(N__54057));
    Odrv12 I__12442 (
            .O(N__54068),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0 ));
    Odrv4 I__12441 (
            .O(N__54065),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0 ));
    Odrv4 I__12440 (
            .O(N__54060),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0 ));
    Odrv4 I__12439 (
            .O(N__54057),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0 ));
    CascadeMux I__12438 (
            .O(N__54048),
            .I(N__54045));
    InMux I__12437 (
            .O(N__54045),
            .I(N__54042));
    LocalMux I__12436 (
            .O(N__54042),
            .I(N__54039));
    Span4Mux_h I__12435 (
            .O(N__54039),
            .I(N__54036));
    Span4Mux_h I__12434 (
            .O(N__54036),
            .I(N__54033));
    Odrv4 I__12433 (
            .O(N__54033),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_1 ));
    CascadeMux I__12432 (
            .O(N__54030),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RLZ0Z7_cascade_ ));
    InMux I__12431 (
            .O(N__54027),
            .I(N__54024));
    LocalMux I__12430 (
            .O(N__54024),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1 ));
    InMux I__12429 (
            .O(N__54021),
            .I(N__54018));
    LocalMux I__12428 (
            .O(N__54018),
            .I(N__54015));
    Span4Mux_v I__12427 (
            .O(N__54015),
            .I(N__54012));
    Odrv4 I__12426 (
            .O(N__54012),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_0 ));
    CascadeMux I__12425 (
            .O(N__54009),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_cascade_ ));
    InMux I__12424 (
            .O(N__54006),
            .I(N__53998));
    InMux I__12423 (
            .O(N__54005),
            .I(N__53995));
    InMux I__12422 (
            .O(N__54004),
            .I(N__53988));
    InMux I__12421 (
            .O(N__54003),
            .I(N__53985));
    InMux I__12420 (
            .O(N__54002),
            .I(N__53980));
    InMux I__12419 (
            .O(N__54001),
            .I(N__53980));
    LocalMux I__12418 (
            .O(N__53998),
            .I(N__53973));
    LocalMux I__12417 (
            .O(N__53995),
            .I(N__53970));
    CascadeMux I__12416 (
            .O(N__53994),
            .I(N__53963));
    InMux I__12415 (
            .O(N__53993),
            .I(N__53956));
    InMux I__12414 (
            .O(N__53992),
            .I(N__53953));
    InMux I__12413 (
            .O(N__53991),
            .I(N__53950));
    LocalMux I__12412 (
            .O(N__53988),
            .I(N__53945));
    LocalMux I__12411 (
            .O(N__53985),
            .I(N__53942));
    LocalMux I__12410 (
            .O(N__53980),
            .I(N__53939));
    InMux I__12409 (
            .O(N__53979),
            .I(N__53934));
    InMux I__12408 (
            .O(N__53978),
            .I(N__53934));
    InMux I__12407 (
            .O(N__53977),
            .I(N__53931));
    InMux I__12406 (
            .O(N__53976),
            .I(N__53928));
    Span4Mux_v I__12405 (
            .O(N__53973),
            .I(N__53925));
    Span4Mux_h I__12404 (
            .O(N__53970),
            .I(N__53922));
    InMux I__12403 (
            .O(N__53969),
            .I(N__53919));
    InMux I__12402 (
            .O(N__53968),
            .I(N__53914));
    InMux I__12401 (
            .O(N__53967),
            .I(N__53914));
    InMux I__12400 (
            .O(N__53966),
            .I(N__53911));
    InMux I__12399 (
            .O(N__53963),
            .I(N__53908));
    InMux I__12398 (
            .O(N__53962),
            .I(N__53905));
    InMux I__12397 (
            .O(N__53961),
            .I(N__53902));
    InMux I__12396 (
            .O(N__53960),
            .I(N__53899));
    InMux I__12395 (
            .O(N__53959),
            .I(N__53896));
    LocalMux I__12394 (
            .O(N__53956),
            .I(N__53893));
    LocalMux I__12393 (
            .O(N__53953),
            .I(N__53888));
    LocalMux I__12392 (
            .O(N__53950),
            .I(N__53888));
    InMux I__12391 (
            .O(N__53949),
            .I(N__53885));
    InMux I__12390 (
            .O(N__53948),
            .I(N__53882));
    Span4Mux_v I__12389 (
            .O(N__53945),
            .I(N__53879));
    Span4Mux_v I__12388 (
            .O(N__53942),
            .I(N__53874));
    Span4Mux_v I__12387 (
            .O(N__53939),
            .I(N__53874));
    LocalMux I__12386 (
            .O(N__53934),
            .I(N__53871));
    LocalMux I__12385 (
            .O(N__53931),
            .I(N__53868));
    LocalMux I__12384 (
            .O(N__53928),
            .I(N__53865));
    Span4Mux_h I__12383 (
            .O(N__53925),
            .I(N__53858));
    Span4Mux_v I__12382 (
            .O(N__53922),
            .I(N__53858));
    LocalMux I__12381 (
            .O(N__53919),
            .I(N__53858));
    LocalMux I__12380 (
            .O(N__53914),
            .I(N__53853));
    LocalMux I__12379 (
            .O(N__53911),
            .I(N__53853));
    LocalMux I__12378 (
            .O(N__53908),
            .I(N__53832));
    LocalMux I__12377 (
            .O(N__53905),
            .I(N__53832));
    LocalMux I__12376 (
            .O(N__53902),
            .I(N__53832));
    LocalMux I__12375 (
            .O(N__53899),
            .I(N__53832));
    LocalMux I__12374 (
            .O(N__53896),
            .I(N__53832));
    Sp12to4 I__12373 (
            .O(N__53893),
            .I(N__53832));
    Span12Mux_v I__12372 (
            .O(N__53888),
            .I(N__53832));
    LocalMux I__12371 (
            .O(N__53885),
            .I(N__53832));
    LocalMux I__12370 (
            .O(N__53882),
            .I(N__53832));
    Sp12to4 I__12369 (
            .O(N__53879),
            .I(N__53832));
    Span4Mux_h I__12368 (
            .O(N__53874),
            .I(N__53827));
    Span4Mux_v I__12367 (
            .O(N__53871),
            .I(N__53827));
    Span4Mux_h I__12366 (
            .O(N__53868),
            .I(N__53824));
    Span4Mux_v I__12365 (
            .O(N__53865),
            .I(N__53819));
    Span4Mux_h I__12364 (
            .O(N__53858),
            .I(N__53819));
    Sp12to4 I__12363 (
            .O(N__53853),
            .I(N__53816));
    Span12Mux_h I__12362 (
            .O(N__53832),
            .I(N__53813));
    Span4Mux_h I__12361 (
            .O(N__53827),
            .I(N__53810));
    Span4Mux_v I__12360 (
            .O(N__53824),
            .I(N__53805));
    Span4Mux_v I__12359 (
            .O(N__53819),
            .I(N__53805));
    Span12Mux_v I__12358 (
            .O(N__53816),
            .I(N__53802));
    Odrv12 I__12357 (
            .O(N__53813),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273 ));
    Odrv4 I__12356 (
            .O(N__53810),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273 ));
    Odrv4 I__12355 (
            .O(N__53805),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273 ));
    Odrv12 I__12354 (
            .O(N__53802),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273 ));
    CascadeMux I__12353 (
            .O(N__53793),
            .I(N__53789));
    InMux I__12352 (
            .O(N__53792),
            .I(N__53785));
    InMux I__12351 (
            .O(N__53789),
            .I(N__53782));
    InMux I__12350 (
            .O(N__53788),
            .I(N__53779));
    LocalMux I__12349 (
            .O(N__53785),
            .I(N__53776));
    LocalMux I__12348 (
            .O(N__53782),
            .I(N__53773));
    LocalMux I__12347 (
            .O(N__53779),
            .I(N__53770));
    Span4Mux_v I__12346 (
            .O(N__53776),
            .I(N__53767));
    Span4Mux_h I__12345 (
            .O(N__53773),
            .I(N__53764));
    Span4Mux_v I__12344 (
            .O(N__53770),
            .I(N__53761));
    Span4Mux_v I__12343 (
            .O(N__53767),
            .I(N__53756));
    Span4Mux_h I__12342 (
            .O(N__53764),
            .I(N__53756));
    Sp12to4 I__12341 (
            .O(N__53761),
            .I(N__53753));
    Span4Mux_v I__12340 (
            .O(N__53756),
            .I(N__53750));
    Odrv12 I__12339 (
            .O(N__53753),
            .I(cemf_module_64ch_ctrl_inst1_data_config_2));
    Odrv4 I__12338 (
            .O(N__53750),
            .I(cemf_module_64ch_ctrl_inst1_data_config_2));
    CascadeMux I__12337 (
            .O(N__53745),
            .I(N__53742));
    InMux I__12336 (
            .O(N__53742),
            .I(N__53739));
    LocalMux I__12335 (
            .O(N__53739),
            .I(N__53736));
    Span4Mux_h I__12334 (
            .O(N__53736),
            .I(N__53733));
    Odrv4 I__12333 (
            .O(N__53733),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_2 ));
    InMux I__12332 (
            .O(N__53730),
            .I(N__53727));
    LocalMux I__12331 (
            .O(N__53727),
            .I(N__53724));
    Odrv12 I__12330 (
            .O(N__53724),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_2 ));
    InMux I__12329 (
            .O(N__53721),
            .I(N__53709));
    InMux I__12328 (
            .O(N__53720),
            .I(N__53704));
    InMux I__12327 (
            .O(N__53719),
            .I(N__53704));
    InMux I__12326 (
            .O(N__53718),
            .I(N__53701));
    InMux I__12325 (
            .O(N__53717),
            .I(N__53696));
    InMux I__12324 (
            .O(N__53716),
            .I(N__53696));
    InMux I__12323 (
            .O(N__53715),
            .I(N__53684));
    InMux I__12322 (
            .O(N__53714),
            .I(N__53684));
    InMux I__12321 (
            .O(N__53713),
            .I(N__53679));
    InMux I__12320 (
            .O(N__53712),
            .I(N__53679));
    LocalMux I__12319 (
            .O(N__53709),
            .I(N__53676));
    LocalMux I__12318 (
            .O(N__53704),
            .I(N__53666));
    LocalMux I__12317 (
            .O(N__53701),
            .I(N__53661));
    LocalMux I__12316 (
            .O(N__53696),
            .I(N__53661));
    InMux I__12315 (
            .O(N__53695),
            .I(N__53656));
    InMux I__12314 (
            .O(N__53694),
            .I(N__53656));
    InMux I__12313 (
            .O(N__53693),
            .I(N__53651));
    InMux I__12312 (
            .O(N__53692),
            .I(N__53651));
    InMux I__12311 (
            .O(N__53691),
            .I(N__53648));
    InMux I__12310 (
            .O(N__53690),
            .I(N__53643));
    InMux I__12309 (
            .O(N__53689),
            .I(N__53643));
    LocalMux I__12308 (
            .O(N__53684),
            .I(N__53640));
    LocalMux I__12307 (
            .O(N__53679),
            .I(N__53637));
    Span4Mux_v I__12306 (
            .O(N__53676),
            .I(N__53634));
    InMux I__12305 (
            .O(N__53675),
            .I(N__53629));
    InMux I__12304 (
            .O(N__53674),
            .I(N__53629));
    InMux I__12303 (
            .O(N__53673),
            .I(N__53626));
    InMux I__12302 (
            .O(N__53672),
            .I(N__53623));
    InMux I__12301 (
            .O(N__53671),
            .I(N__53620));
    InMux I__12300 (
            .O(N__53670),
            .I(N__53615));
    InMux I__12299 (
            .O(N__53669),
            .I(N__53615));
    Span4Mux_h I__12298 (
            .O(N__53666),
            .I(N__53610));
    Span4Mux_v I__12297 (
            .O(N__53661),
            .I(N__53610));
    LocalMux I__12296 (
            .O(N__53656),
            .I(N__53607));
    LocalMux I__12295 (
            .O(N__53651),
            .I(N__53596));
    LocalMux I__12294 (
            .O(N__53648),
            .I(N__53596));
    LocalMux I__12293 (
            .O(N__53643),
            .I(N__53596));
    Span4Mux_v I__12292 (
            .O(N__53640),
            .I(N__53596));
    Span4Mux_v I__12291 (
            .O(N__53637),
            .I(N__53596));
    Span4Mux_h I__12290 (
            .O(N__53634),
            .I(N__53593));
    LocalMux I__12289 (
            .O(N__53629),
            .I(N__53588));
    LocalMux I__12288 (
            .O(N__53626),
            .I(N__53588));
    LocalMux I__12287 (
            .O(N__53623),
            .I(N__53585));
    LocalMux I__12286 (
            .O(N__53620),
            .I(N__53578));
    LocalMux I__12285 (
            .O(N__53615),
            .I(N__53578));
    Span4Mux_h I__12284 (
            .O(N__53610),
            .I(N__53578));
    Span4Mux_v I__12283 (
            .O(N__53607),
            .I(N__53573));
    Span4Mux_h I__12282 (
            .O(N__53596),
            .I(N__53573));
    Span4Mux_v I__12281 (
            .O(N__53593),
            .I(N__53568));
    Span4Mux_v I__12280 (
            .O(N__53588),
            .I(N__53568));
    Sp12to4 I__12279 (
            .O(N__53585),
            .I(N__53565));
    Span4Mux_h I__12278 (
            .O(N__53578),
            .I(N__53562));
    Span4Mux_v I__12277 (
            .O(N__53573),
            .I(N__53559));
    Span4Mux_h I__12276 (
            .O(N__53568),
            .I(N__53556));
    Odrv12 I__12275 (
            .O(N__53565),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i ));
    Odrv4 I__12274 (
            .O(N__53562),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i ));
    Odrv4 I__12273 (
            .O(N__53559),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i ));
    Odrv4 I__12272 (
            .O(N__53556),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i ));
    CascadeMux I__12271 (
            .O(N__53547),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGHZ0Z5_cascade_ ));
    InMux I__12270 (
            .O(N__53544),
            .I(N__53541));
    LocalMux I__12269 (
            .O(N__53541),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17 ));
    CascadeMux I__12268 (
            .O(N__53538),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17_cascade_ ));
    InMux I__12267 (
            .O(N__53535),
            .I(N__53532));
    LocalMux I__12266 (
            .O(N__53532),
            .I(N__53529));
    Odrv12 I__12265 (
            .O(N__53529),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_17 ));
    InMux I__12264 (
            .O(N__53526),
            .I(N__53521));
    CascadeMux I__12263 (
            .O(N__53525),
            .I(N__53518));
    InMux I__12262 (
            .O(N__53524),
            .I(N__53515));
    LocalMux I__12261 (
            .O(N__53521),
            .I(N__53512));
    InMux I__12260 (
            .O(N__53518),
            .I(N__53509));
    LocalMux I__12259 (
            .O(N__53515),
            .I(N__53504));
    Span4Mux_h I__12258 (
            .O(N__53512),
            .I(N__53504));
    LocalMux I__12257 (
            .O(N__53509),
            .I(N__53501));
    Odrv4 I__12256 (
            .O(N__53504),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_16));
    Odrv4 I__12255 (
            .O(N__53501),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_16));
    CascadeMux I__12254 (
            .O(N__53496),
            .I(N__53493));
    InMux I__12253 (
            .O(N__53493),
            .I(N__53490));
    LocalMux I__12252 (
            .O(N__53490),
            .I(N__53487));
    Span4Mux_h I__12251 (
            .O(N__53487),
            .I(N__53484));
    Odrv4 I__12250 (
            .O(N__53484),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_16 ));
    InMux I__12249 (
            .O(N__53481),
            .I(N__53478));
    LocalMux I__12248 (
            .O(N__53478),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_16 ));
    CascadeMux I__12247 (
            .O(N__53475),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGHZ0Z5_cascade_ ));
    InMux I__12246 (
            .O(N__53472),
            .I(N__53469));
    LocalMux I__12245 (
            .O(N__53469),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16 ));
    InMux I__12244 (
            .O(N__53466),
            .I(N__53463));
    LocalMux I__12243 (
            .O(N__53463),
            .I(N__53460));
    Odrv12 I__12242 (
            .O(N__53460),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_15 ));
    CascadeMux I__12241 (
            .O(N__53457),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16_cascade_ ));
    InMux I__12240 (
            .O(N__53454),
            .I(N__53451));
    LocalMux I__12239 (
            .O(N__53451),
            .I(N__53448));
    Odrv4 I__12238 (
            .O(N__53448),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_16 ));
    InMux I__12237 (
            .O(N__53445),
            .I(N__53442));
    LocalMux I__12236 (
            .O(N__53442),
            .I(N__53439));
    Span12Mux_v I__12235 (
            .O(N__53439),
            .I(N__53436));
    Span12Mux_h I__12234 (
            .O(N__53436),
            .I(N__53433));
    Odrv12 I__12233 (
            .O(N__53433),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_31));
    CascadeMux I__12232 (
            .O(N__53430),
            .I(N__53427));
    InMux I__12231 (
            .O(N__53427),
            .I(N__53424));
    LocalMux I__12230 (
            .O(N__53424),
            .I(N__53421));
    Span4Mux_h I__12229 (
            .O(N__53421),
            .I(N__53416));
    InMux I__12228 (
            .O(N__53420),
            .I(N__53413));
    InMux I__12227 (
            .O(N__53419),
            .I(N__53410));
    Span4Mux_h I__12226 (
            .O(N__53416),
            .I(N__53407));
    LocalMux I__12225 (
            .O(N__53413),
            .I(N__53404));
    LocalMux I__12224 (
            .O(N__53410),
            .I(N__53401));
    Span4Mux_h I__12223 (
            .O(N__53407),
            .I(N__53398));
    Span4Mux_v I__12222 (
            .O(N__53404),
            .I(N__53393));
    Span4Mux_h I__12221 (
            .O(N__53401),
            .I(N__53393));
    Span4Mux_h I__12220 (
            .O(N__53398),
            .I(N__53390));
    Span4Mux_h I__12219 (
            .O(N__53393),
            .I(N__53387));
    Odrv4 I__12218 (
            .O(N__53390),
            .I(cemf_module_64ch_ctrl_inst1_data_config_14));
    Odrv4 I__12217 (
            .O(N__53387),
            .I(cemf_module_64ch_ctrl_inst1_data_config_14));
    CascadeMux I__12216 (
            .O(N__53382),
            .I(N__53379));
    InMux I__12215 (
            .O(N__53379),
            .I(N__53376));
    LocalMux I__12214 (
            .O(N__53376),
            .I(N__53372));
    InMux I__12213 (
            .O(N__53375),
            .I(N__53368));
    Span4Mux_v I__12212 (
            .O(N__53372),
            .I(N__53365));
    InMux I__12211 (
            .O(N__53371),
            .I(N__53362));
    LocalMux I__12210 (
            .O(N__53368),
            .I(N__53359));
    Span4Mux_h I__12209 (
            .O(N__53365),
            .I(N__53356));
    LocalMux I__12208 (
            .O(N__53362),
            .I(N__53351));
    Span4Mux_h I__12207 (
            .O(N__53359),
            .I(N__53351));
    Span4Mux_h I__12206 (
            .O(N__53356),
            .I(N__53348));
    Span4Mux_h I__12205 (
            .O(N__53351),
            .I(N__53345));
    Odrv4 I__12204 (
            .O(N__53348),
            .I(cemf_module_64ch_ctrl_inst1_data_config_15));
    Odrv4 I__12203 (
            .O(N__53345),
            .I(cemf_module_64ch_ctrl_inst1_data_config_15));
    InMux I__12202 (
            .O(N__53340),
            .I(N__53337));
    LocalMux I__12201 (
            .O(N__53337),
            .I(N__53334));
    Odrv4 I__12200 (
            .O(N__53334),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_25));
    InMux I__12199 (
            .O(N__53331),
            .I(N__53325));
    CascadeMux I__12198 (
            .O(N__53330),
            .I(N__53320));
    CascadeMux I__12197 (
            .O(N__53329),
            .I(N__53311));
    CascadeMux I__12196 (
            .O(N__53328),
            .I(N__53307));
    LocalMux I__12195 (
            .O(N__53325),
            .I(N__53303));
    CascadeMux I__12194 (
            .O(N__53324),
            .I(N__53300));
    CascadeMux I__12193 (
            .O(N__53323),
            .I(N__53297));
    InMux I__12192 (
            .O(N__53320),
            .I(N__53293));
    CascadeMux I__12191 (
            .O(N__53319),
            .I(N__53290));
    CascadeMux I__12190 (
            .O(N__53318),
            .I(N__53287));
    CascadeMux I__12189 (
            .O(N__53317),
            .I(N__53283));
    CascadeMux I__12188 (
            .O(N__53316),
            .I(N__53278));
    CascadeMux I__12187 (
            .O(N__53315),
            .I(N__53275));
    InMux I__12186 (
            .O(N__53314),
            .I(N__53272));
    InMux I__12185 (
            .O(N__53311),
            .I(N__53267));
    CascadeMux I__12184 (
            .O(N__53310),
            .I(N__53263));
    InMux I__12183 (
            .O(N__53307),
            .I(N__53259));
    CascadeMux I__12182 (
            .O(N__53306),
            .I(N__53253));
    Span4Mux_v I__12181 (
            .O(N__53303),
            .I(N__53250));
    InMux I__12180 (
            .O(N__53300),
            .I(N__53247));
    InMux I__12179 (
            .O(N__53297),
            .I(N__53244));
    InMux I__12178 (
            .O(N__53296),
            .I(N__53241));
    LocalMux I__12177 (
            .O(N__53293),
            .I(N__53238));
    InMux I__12176 (
            .O(N__53290),
            .I(N__53235));
    InMux I__12175 (
            .O(N__53287),
            .I(N__53232));
    InMux I__12174 (
            .O(N__53286),
            .I(N__53229));
    InMux I__12173 (
            .O(N__53283),
            .I(N__53226));
    InMux I__12172 (
            .O(N__53282),
            .I(N__53223));
    InMux I__12171 (
            .O(N__53281),
            .I(N__53220));
    InMux I__12170 (
            .O(N__53278),
            .I(N__53217));
    InMux I__12169 (
            .O(N__53275),
            .I(N__53214));
    LocalMux I__12168 (
            .O(N__53272),
            .I(N__53211));
    InMux I__12167 (
            .O(N__53271),
            .I(N__53208));
    InMux I__12166 (
            .O(N__53270),
            .I(N__53205));
    LocalMux I__12165 (
            .O(N__53267),
            .I(N__53202));
    InMux I__12164 (
            .O(N__53266),
            .I(N__53199));
    InMux I__12163 (
            .O(N__53263),
            .I(N__53196));
    CascadeMux I__12162 (
            .O(N__53262),
            .I(N__53191));
    LocalMux I__12161 (
            .O(N__53259),
            .I(N__53188));
    InMux I__12160 (
            .O(N__53258),
            .I(N__53185));
    InMux I__12159 (
            .O(N__53257),
            .I(N__53182));
    CascadeMux I__12158 (
            .O(N__53256),
            .I(N__53176));
    InMux I__12157 (
            .O(N__53253),
            .I(N__53172));
    Span4Mux_h I__12156 (
            .O(N__53250),
            .I(N__53167));
    LocalMux I__12155 (
            .O(N__53247),
            .I(N__53167));
    LocalMux I__12154 (
            .O(N__53244),
            .I(N__53162));
    LocalMux I__12153 (
            .O(N__53241),
            .I(N__53162));
    Span4Mux_v I__12152 (
            .O(N__53238),
            .I(N__53157));
    LocalMux I__12151 (
            .O(N__53235),
            .I(N__53157));
    LocalMux I__12150 (
            .O(N__53232),
            .I(N__53154));
    LocalMux I__12149 (
            .O(N__53229),
            .I(N__53147));
    LocalMux I__12148 (
            .O(N__53226),
            .I(N__53147));
    LocalMux I__12147 (
            .O(N__53223),
            .I(N__53147));
    LocalMux I__12146 (
            .O(N__53220),
            .I(N__53142));
    LocalMux I__12145 (
            .O(N__53217),
            .I(N__53142));
    LocalMux I__12144 (
            .O(N__53214),
            .I(N__53137));
    Span4Mux_h I__12143 (
            .O(N__53211),
            .I(N__53137));
    LocalMux I__12142 (
            .O(N__53208),
            .I(N__53130));
    LocalMux I__12141 (
            .O(N__53205),
            .I(N__53130));
    Span4Mux_h I__12140 (
            .O(N__53202),
            .I(N__53130));
    LocalMux I__12139 (
            .O(N__53199),
            .I(N__53127));
    LocalMux I__12138 (
            .O(N__53196),
            .I(N__53124));
    InMux I__12137 (
            .O(N__53195),
            .I(N__53119));
    InMux I__12136 (
            .O(N__53194),
            .I(N__53119));
    InMux I__12135 (
            .O(N__53191),
            .I(N__53116));
    Span4Mux_h I__12134 (
            .O(N__53188),
            .I(N__53111));
    LocalMux I__12133 (
            .O(N__53185),
            .I(N__53111));
    LocalMux I__12132 (
            .O(N__53182),
            .I(N__53108));
    InMux I__12131 (
            .O(N__53181),
            .I(N__53097));
    InMux I__12130 (
            .O(N__53180),
            .I(N__53097));
    InMux I__12129 (
            .O(N__53179),
            .I(N__53097));
    InMux I__12128 (
            .O(N__53176),
            .I(N__53097));
    InMux I__12127 (
            .O(N__53175),
            .I(N__53097));
    LocalMux I__12126 (
            .O(N__53172),
            .I(N__53090));
    Span4Mux_h I__12125 (
            .O(N__53167),
            .I(N__53090));
    Span4Mux_h I__12124 (
            .O(N__53162),
            .I(N__53090));
    Span4Mux_v I__12123 (
            .O(N__53157),
            .I(N__53087));
    Span4Mux_v I__12122 (
            .O(N__53154),
            .I(N__53082));
    Span4Mux_h I__12121 (
            .O(N__53147),
            .I(N__53082));
    Span4Mux_v I__12120 (
            .O(N__53142),
            .I(N__53075));
    Span4Mux_h I__12119 (
            .O(N__53137),
            .I(N__53075));
    Span4Mux_v I__12118 (
            .O(N__53130),
            .I(N__53075));
    Span4Mux_h I__12117 (
            .O(N__53127),
            .I(N__53068));
    Span4Mux_v I__12116 (
            .O(N__53124),
            .I(N__53068));
    LocalMux I__12115 (
            .O(N__53119),
            .I(N__53068));
    LocalMux I__12114 (
            .O(N__53116),
            .I(N__53059));
    Span4Mux_v I__12113 (
            .O(N__53111),
            .I(N__53059));
    Span4Mux_h I__12112 (
            .O(N__53108),
            .I(N__53059));
    LocalMux I__12111 (
            .O(N__53097),
            .I(N__53059));
    Span4Mux_v I__12110 (
            .O(N__53090),
            .I(N__53056));
    Sp12to4 I__12109 (
            .O(N__53087),
            .I(N__53053));
    Span4Mux_v I__12108 (
            .O(N__53082),
            .I(N__53048));
    Span4Mux_h I__12107 (
            .O(N__53075),
            .I(N__53048));
    Span4Mux_h I__12106 (
            .O(N__53068),
            .I(N__53043));
    Span4Mux_h I__12105 (
            .O(N__53059),
            .I(N__53043));
    Odrv4 I__12104 (
            .O(N__53056),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0 ));
    Odrv12 I__12103 (
            .O(N__53053),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0 ));
    Odrv4 I__12102 (
            .O(N__53048),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0 ));
    Odrv4 I__12101 (
            .O(N__53043),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0 ));
    CascadeMux I__12100 (
            .O(N__53034),
            .I(N__53031));
    InMux I__12099 (
            .O(N__53031),
            .I(N__53028));
    LocalMux I__12098 (
            .O(N__53028),
            .I(N__53025));
    Span4Mux_v I__12097 (
            .O(N__53025),
            .I(N__53022));
    Sp12to4 I__12096 (
            .O(N__53022),
            .I(N__53019));
    Odrv12 I__12095 (
            .O(N__53019),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_25));
    InMux I__12094 (
            .O(N__53016),
            .I(N__53005));
    InMux I__12093 (
            .O(N__53015),
            .I(N__53001));
    InMux I__12092 (
            .O(N__53014),
            .I(N__52995));
    CascadeMux I__12091 (
            .O(N__53013),
            .I(N__52991));
    InMux I__12090 (
            .O(N__53012),
            .I(N__52984));
    InMux I__12089 (
            .O(N__53011),
            .I(N__52979));
    InMux I__12088 (
            .O(N__53010),
            .I(N__52976));
    InMux I__12087 (
            .O(N__53009),
            .I(N__52973));
    InMux I__12086 (
            .O(N__53008),
            .I(N__52970));
    LocalMux I__12085 (
            .O(N__53005),
            .I(N__52967));
    InMux I__12084 (
            .O(N__53004),
            .I(N__52964));
    LocalMux I__12083 (
            .O(N__53001),
            .I(N__52961));
    InMux I__12082 (
            .O(N__53000),
            .I(N__52958));
    InMux I__12081 (
            .O(N__52999),
            .I(N__52955));
    InMux I__12080 (
            .O(N__52998),
            .I(N__52952));
    LocalMux I__12079 (
            .O(N__52995),
            .I(N__52949));
    InMux I__12078 (
            .O(N__52994),
            .I(N__52946));
    InMux I__12077 (
            .O(N__52991),
            .I(N__52943));
    InMux I__12076 (
            .O(N__52990),
            .I(N__52940));
    InMux I__12075 (
            .O(N__52989),
            .I(N__52937));
    InMux I__12074 (
            .O(N__52988),
            .I(N__52934));
    InMux I__12073 (
            .O(N__52987),
            .I(N__52931));
    LocalMux I__12072 (
            .O(N__52984),
            .I(N__52928));
    InMux I__12071 (
            .O(N__52983),
            .I(N__52919));
    InMux I__12070 (
            .O(N__52982),
            .I(N__52916));
    LocalMux I__12069 (
            .O(N__52979),
            .I(N__52911));
    LocalMux I__12068 (
            .O(N__52976),
            .I(N__52911));
    LocalMux I__12067 (
            .O(N__52973),
            .I(N__52908));
    LocalMux I__12066 (
            .O(N__52970),
            .I(N__52905));
    Span4Mux_h I__12065 (
            .O(N__52967),
            .I(N__52894));
    LocalMux I__12064 (
            .O(N__52964),
            .I(N__52894));
    Span4Mux_v I__12063 (
            .O(N__52961),
            .I(N__52894));
    LocalMux I__12062 (
            .O(N__52958),
            .I(N__52885));
    LocalMux I__12061 (
            .O(N__52955),
            .I(N__52885));
    LocalMux I__12060 (
            .O(N__52952),
            .I(N__52885));
    Span4Mux_v I__12059 (
            .O(N__52949),
            .I(N__52885));
    LocalMux I__12058 (
            .O(N__52946),
            .I(N__52882));
    LocalMux I__12057 (
            .O(N__52943),
            .I(N__52877));
    LocalMux I__12056 (
            .O(N__52940),
            .I(N__52877));
    LocalMux I__12055 (
            .O(N__52937),
            .I(N__52872));
    LocalMux I__12054 (
            .O(N__52934),
            .I(N__52872));
    LocalMux I__12053 (
            .O(N__52931),
            .I(N__52867));
    Span4Mux_v I__12052 (
            .O(N__52928),
            .I(N__52867));
    InMux I__12051 (
            .O(N__52927),
            .I(N__52854));
    InMux I__12050 (
            .O(N__52926),
            .I(N__52854));
    InMux I__12049 (
            .O(N__52925),
            .I(N__52854));
    InMux I__12048 (
            .O(N__52924),
            .I(N__52854));
    InMux I__12047 (
            .O(N__52923),
            .I(N__52854));
    InMux I__12046 (
            .O(N__52922),
            .I(N__52854));
    LocalMux I__12045 (
            .O(N__52919),
            .I(N__52847));
    LocalMux I__12044 (
            .O(N__52916),
            .I(N__52847));
    Span4Mux_h I__12043 (
            .O(N__52911),
            .I(N__52847));
    Span4Mux_h I__12042 (
            .O(N__52908),
            .I(N__52842));
    Span4Mux_v I__12041 (
            .O(N__52905),
            .I(N__52842));
    InMux I__12040 (
            .O(N__52904),
            .I(N__52833));
    InMux I__12039 (
            .O(N__52903),
            .I(N__52833));
    InMux I__12038 (
            .O(N__52902),
            .I(N__52833));
    InMux I__12037 (
            .O(N__52901),
            .I(N__52833));
    Span4Mux_h I__12036 (
            .O(N__52894),
            .I(N__52830));
    Span4Mux_h I__12035 (
            .O(N__52885),
            .I(N__52827));
    Span4Mux_v I__12034 (
            .O(N__52882),
            .I(N__52816));
    Span4Mux_v I__12033 (
            .O(N__52877),
            .I(N__52816));
    Span4Mux_v I__12032 (
            .O(N__52872),
            .I(N__52816));
    Span4Mux_h I__12031 (
            .O(N__52867),
            .I(N__52816));
    LocalMux I__12030 (
            .O(N__52854),
            .I(N__52816));
    Odrv4 I__12029 (
            .O(N__52847),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ));
    Odrv4 I__12028 (
            .O(N__52842),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ));
    LocalMux I__12027 (
            .O(N__52833),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ));
    Odrv4 I__12026 (
            .O(N__52830),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ));
    Odrv4 I__12025 (
            .O(N__52827),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ));
    Odrv4 I__12024 (
            .O(N__52816),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ));
    InMux I__12023 (
            .O(N__52803),
            .I(N__52800));
    LocalMux I__12022 (
            .O(N__52800),
            .I(N__52797));
    Span4Mux_v I__12021 (
            .O(N__52797),
            .I(N__52794));
    Span4Mux_h I__12020 (
            .O(N__52794),
            .I(N__52791));
    Span4Mux_v I__12019 (
            .O(N__52791),
            .I(N__52788));
    Sp12to4 I__12018 (
            .O(N__52788),
            .I(N__52785));
    Odrv12 I__12017 (
            .O(N__52785),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_25));
    InMux I__12016 (
            .O(N__52782),
            .I(N__52776));
    InMux I__12015 (
            .O(N__52781),
            .I(N__52773));
    InMux I__12014 (
            .O(N__52780),
            .I(N__52765));
    InMux I__12013 (
            .O(N__52779),
            .I(N__52762));
    LocalMux I__12012 (
            .O(N__52776),
            .I(N__52757));
    LocalMux I__12011 (
            .O(N__52773),
            .I(N__52752));
    InMux I__12010 (
            .O(N__52772),
            .I(N__52749));
    InMux I__12009 (
            .O(N__52771),
            .I(N__52746));
    InMux I__12008 (
            .O(N__52770),
            .I(N__52733));
    InMux I__12007 (
            .O(N__52769),
            .I(N__52730));
    InMux I__12006 (
            .O(N__52768),
            .I(N__52727));
    LocalMux I__12005 (
            .O(N__52765),
            .I(N__52722));
    LocalMux I__12004 (
            .O(N__52762),
            .I(N__52722));
    InMux I__12003 (
            .O(N__52761),
            .I(N__52719));
    InMux I__12002 (
            .O(N__52760),
            .I(N__52716));
    Span4Mux_v I__12001 (
            .O(N__52757),
            .I(N__52713));
    InMux I__12000 (
            .O(N__52756),
            .I(N__52710));
    InMux I__11999 (
            .O(N__52755),
            .I(N__52707));
    Span4Mux_h I__11998 (
            .O(N__52752),
            .I(N__52702));
    LocalMux I__11997 (
            .O(N__52749),
            .I(N__52702));
    LocalMux I__11996 (
            .O(N__52746),
            .I(N__52697));
    InMux I__11995 (
            .O(N__52745),
            .I(N__52694));
    InMux I__11994 (
            .O(N__52744),
            .I(N__52691));
    InMux I__11993 (
            .O(N__52743),
            .I(N__52688));
    InMux I__11992 (
            .O(N__52742),
            .I(N__52685));
    InMux I__11991 (
            .O(N__52741),
            .I(N__52682));
    InMux I__11990 (
            .O(N__52740),
            .I(N__52677));
    InMux I__11989 (
            .O(N__52739),
            .I(N__52677));
    InMux I__11988 (
            .O(N__52738),
            .I(N__52669));
    InMux I__11987 (
            .O(N__52737),
            .I(N__52666));
    InMux I__11986 (
            .O(N__52736),
            .I(N__52663));
    LocalMux I__11985 (
            .O(N__52733),
            .I(N__52660));
    LocalMux I__11984 (
            .O(N__52730),
            .I(N__52657));
    LocalMux I__11983 (
            .O(N__52727),
            .I(N__52648));
    Span4Mux_v I__11982 (
            .O(N__52722),
            .I(N__52648));
    LocalMux I__11981 (
            .O(N__52719),
            .I(N__52648));
    LocalMux I__11980 (
            .O(N__52716),
            .I(N__52648));
    Span4Mux_h I__11979 (
            .O(N__52713),
            .I(N__52643));
    LocalMux I__11978 (
            .O(N__52710),
            .I(N__52643));
    LocalMux I__11977 (
            .O(N__52707),
            .I(N__52640));
    Span4Mux_h I__11976 (
            .O(N__52702),
            .I(N__52637));
    InMux I__11975 (
            .O(N__52701),
            .I(N__52634));
    InMux I__11974 (
            .O(N__52700),
            .I(N__52631));
    Span4Mux_v I__11973 (
            .O(N__52697),
            .I(N__52626));
    LocalMux I__11972 (
            .O(N__52694),
            .I(N__52626));
    LocalMux I__11971 (
            .O(N__52691),
            .I(N__52621));
    LocalMux I__11970 (
            .O(N__52688),
            .I(N__52621));
    LocalMux I__11969 (
            .O(N__52685),
            .I(N__52614));
    LocalMux I__11968 (
            .O(N__52682),
            .I(N__52614));
    LocalMux I__11967 (
            .O(N__52677),
            .I(N__52614));
    InMux I__11966 (
            .O(N__52676),
            .I(N__52611));
    InMux I__11965 (
            .O(N__52675),
            .I(N__52608));
    InMux I__11964 (
            .O(N__52674),
            .I(N__52605));
    InMux I__11963 (
            .O(N__52673),
            .I(N__52602));
    InMux I__11962 (
            .O(N__52672),
            .I(N__52599));
    LocalMux I__11961 (
            .O(N__52669),
            .I(N__52592));
    LocalMux I__11960 (
            .O(N__52666),
            .I(N__52592));
    LocalMux I__11959 (
            .O(N__52663),
            .I(N__52592));
    Span4Mux_h I__11958 (
            .O(N__52660),
            .I(N__52585));
    Span4Mux_v I__11957 (
            .O(N__52657),
            .I(N__52585));
    Span4Mux_h I__11956 (
            .O(N__52648),
            .I(N__52585));
    Span4Mux_h I__11955 (
            .O(N__52643),
            .I(N__52578));
    Span4Mux_h I__11954 (
            .O(N__52640),
            .I(N__52578));
    Span4Mux_h I__11953 (
            .O(N__52637),
            .I(N__52578));
    LocalMux I__11952 (
            .O(N__52634),
            .I(N__52567));
    LocalMux I__11951 (
            .O(N__52631),
            .I(N__52567));
    Span4Mux_h I__11950 (
            .O(N__52626),
            .I(N__52567));
    Span4Mux_v I__11949 (
            .O(N__52621),
            .I(N__52567));
    Span4Mux_v I__11948 (
            .O(N__52614),
            .I(N__52567));
    LocalMux I__11947 (
            .O(N__52611),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    LocalMux I__11946 (
            .O(N__52608),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    LocalMux I__11945 (
            .O(N__52605),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    LocalMux I__11944 (
            .O(N__52602),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    LocalMux I__11943 (
            .O(N__52599),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    Odrv12 I__11942 (
            .O(N__52592),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    Odrv4 I__11941 (
            .O(N__52585),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    Odrv4 I__11940 (
            .O(N__52578),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    Odrv4 I__11939 (
            .O(N__52567),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ));
    CascadeMux I__11938 (
            .O(N__52548),
            .I(N__52545));
    InMux I__11937 (
            .O(N__52545),
            .I(N__52542));
    LocalMux I__11936 (
            .O(N__52542),
            .I(N__52539));
    Span4Mux_v I__11935 (
            .O(N__52539),
            .I(N__52536));
    Span4Mux_h I__11934 (
            .O(N__52536),
            .I(N__52533));
    Sp12to4 I__11933 (
            .O(N__52533),
            .I(N__52530));
    Odrv12 I__11932 (
            .O(N__52530),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_25));
    InMux I__11931 (
            .O(N__52527),
            .I(N__52517));
    InMux I__11930 (
            .O(N__52526),
            .I(N__52514));
    InMux I__11929 (
            .O(N__52525),
            .I(N__52509));
    InMux I__11928 (
            .O(N__52524),
            .I(N__52506));
    InMux I__11927 (
            .O(N__52523),
            .I(N__52503));
    InMux I__11926 (
            .O(N__52522),
            .I(N__52500));
    InMux I__11925 (
            .O(N__52521),
            .I(N__52497));
    InMux I__11924 (
            .O(N__52520),
            .I(N__52489));
    LocalMux I__11923 (
            .O(N__52517),
            .I(N__52481));
    LocalMux I__11922 (
            .O(N__52514),
            .I(N__52478));
    InMux I__11921 (
            .O(N__52513),
            .I(N__52475));
    InMux I__11920 (
            .O(N__52512),
            .I(N__52472));
    LocalMux I__11919 (
            .O(N__52509),
            .I(N__52468));
    LocalMux I__11918 (
            .O(N__52506),
            .I(N__52463));
    LocalMux I__11917 (
            .O(N__52503),
            .I(N__52463));
    LocalMux I__11916 (
            .O(N__52500),
            .I(N__52458));
    LocalMux I__11915 (
            .O(N__52497),
            .I(N__52458));
    InMux I__11914 (
            .O(N__52496),
            .I(N__52455));
    InMux I__11913 (
            .O(N__52495),
            .I(N__52450));
    InMux I__11912 (
            .O(N__52494),
            .I(N__52450));
    InMux I__11911 (
            .O(N__52493),
            .I(N__52447));
    InMux I__11910 (
            .O(N__52492),
            .I(N__52442));
    LocalMux I__11909 (
            .O(N__52489),
            .I(N__52434));
    InMux I__11908 (
            .O(N__52488),
            .I(N__52431));
    InMux I__11907 (
            .O(N__52487),
            .I(N__52428));
    InMux I__11906 (
            .O(N__52486),
            .I(N__52425));
    InMux I__11905 (
            .O(N__52485),
            .I(N__52422));
    InMux I__11904 (
            .O(N__52484),
            .I(N__52419));
    Span4Mux_h I__11903 (
            .O(N__52481),
            .I(N__52410));
    Span4Mux_h I__11902 (
            .O(N__52478),
            .I(N__52410));
    LocalMux I__11901 (
            .O(N__52475),
            .I(N__52410));
    LocalMux I__11900 (
            .O(N__52472),
            .I(N__52410));
    InMux I__11899 (
            .O(N__52471),
            .I(N__52407));
    Span4Mux_v I__11898 (
            .O(N__52468),
            .I(N__52404));
    Span4Mux_v I__11897 (
            .O(N__52463),
            .I(N__52399));
    Span4Mux_h I__11896 (
            .O(N__52458),
            .I(N__52399));
    LocalMux I__11895 (
            .O(N__52455),
            .I(N__52396));
    LocalMux I__11894 (
            .O(N__52450),
            .I(N__52391));
    LocalMux I__11893 (
            .O(N__52447),
            .I(N__52391));
    InMux I__11892 (
            .O(N__52446),
            .I(N__52388));
    InMux I__11891 (
            .O(N__52445),
            .I(N__52385));
    LocalMux I__11890 (
            .O(N__52442),
            .I(N__52382));
    InMux I__11889 (
            .O(N__52441),
            .I(N__52378));
    InMux I__11888 (
            .O(N__52440),
            .I(N__52375));
    InMux I__11887 (
            .O(N__52439),
            .I(N__52372));
    InMux I__11886 (
            .O(N__52438),
            .I(N__52367));
    InMux I__11885 (
            .O(N__52437),
            .I(N__52364));
    Span4Mux_h I__11884 (
            .O(N__52434),
            .I(N__52357));
    LocalMux I__11883 (
            .O(N__52431),
            .I(N__52357));
    LocalMux I__11882 (
            .O(N__52428),
            .I(N__52357));
    LocalMux I__11881 (
            .O(N__52425),
            .I(N__52354));
    LocalMux I__11880 (
            .O(N__52422),
            .I(N__52349));
    LocalMux I__11879 (
            .O(N__52419),
            .I(N__52349));
    Span4Mux_h I__11878 (
            .O(N__52410),
            .I(N__52344));
    LocalMux I__11877 (
            .O(N__52407),
            .I(N__52344));
    Span4Mux_h I__11876 (
            .O(N__52404),
            .I(N__52333));
    Span4Mux_h I__11875 (
            .O(N__52399),
            .I(N__52333));
    Span4Mux_v I__11874 (
            .O(N__52396),
            .I(N__52333));
    Span4Mux_v I__11873 (
            .O(N__52391),
            .I(N__52333));
    LocalMux I__11872 (
            .O(N__52388),
            .I(N__52333));
    LocalMux I__11871 (
            .O(N__52385),
            .I(N__52330));
    Span4Mux_h I__11870 (
            .O(N__52382),
            .I(N__52327));
    InMux I__11869 (
            .O(N__52381),
            .I(N__52324));
    LocalMux I__11868 (
            .O(N__52378),
            .I(N__52319));
    LocalMux I__11867 (
            .O(N__52375),
            .I(N__52319));
    LocalMux I__11866 (
            .O(N__52372),
            .I(N__52316));
    InMux I__11865 (
            .O(N__52371),
            .I(N__52311));
    InMux I__11864 (
            .O(N__52370),
            .I(N__52311));
    LocalMux I__11863 (
            .O(N__52367),
            .I(N__52308));
    LocalMux I__11862 (
            .O(N__52364),
            .I(N__52303));
    Span4Mux_v I__11861 (
            .O(N__52357),
            .I(N__52303));
    Span4Mux_h I__11860 (
            .O(N__52354),
            .I(N__52298));
    Span4Mux_h I__11859 (
            .O(N__52349),
            .I(N__52298));
    Span4Mux_v I__11858 (
            .O(N__52344),
            .I(N__52293));
    Span4Mux_h I__11857 (
            .O(N__52333),
            .I(N__52293));
    Span4Mux_h I__11856 (
            .O(N__52330),
            .I(N__52284));
    Span4Mux_h I__11855 (
            .O(N__52327),
            .I(N__52284));
    LocalMux I__11854 (
            .O(N__52324),
            .I(N__52284));
    Span4Mux_v I__11853 (
            .O(N__52319),
            .I(N__52284));
    Span4Mux_v I__11852 (
            .O(N__52316),
            .I(N__52279));
    LocalMux I__11851 (
            .O(N__52311),
            .I(N__52279));
    Span12Mux_v I__11850 (
            .O(N__52308),
            .I(N__52276));
    Span4Mux_h I__11849 (
            .O(N__52303),
            .I(N__52271));
    Span4Mux_v I__11848 (
            .O(N__52298),
            .I(N__52271));
    Span4Mux_v I__11847 (
            .O(N__52293),
            .I(N__52268));
    Span4Mux_v I__11846 (
            .O(N__52284),
            .I(N__52263));
    Span4Mux_h I__11845 (
            .O(N__52279),
            .I(N__52263));
    Odrv12 I__11844 (
            .O(N__52276),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1314 ));
    Odrv4 I__11843 (
            .O(N__52271),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1314 ));
    Odrv4 I__11842 (
            .O(N__52268),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1314 ));
    Odrv4 I__11841 (
            .O(N__52263),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1314 ));
    InMux I__11840 (
            .O(N__52254),
            .I(N__52251));
    LocalMux I__11839 (
            .O(N__52251),
            .I(N__52248));
    Span4Mux_h I__11838 (
            .O(N__52248),
            .I(N__52245));
    Span4Mux_v I__11837 (
            .O(N__52245),
            .I(N__52242));
    Odrv4 I__11836 (
            .O(N__52242),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_25));
    CascadeMux I__11835 (
            .O(N__52239),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_25_cascade_ ));
    InMux I__11834 (
            .O(N__52236),
            .I(N__52228));
    InMux I__11833 (
            .O(N__52235),
            .I(N__52224));
    InMux I__11832 (
            .O(N__52234),
            .I(N__52217));
    InMux I__11831 (
            .O(N__52233),
            .I(N__52210));
    InMux I__11830 (
            .O(N__52232),
            .I(N__52207));
    InMux I__11829 (
            .O(N__52231),
            .I(N__52200));
    LocalMux I__11828 (
            .O(N__52228),
            .I(N__52195));
    InMux I__11827 (
            .O(N__52227),
            .I(N__52192));
    LocalMux I__11826 (
            .O(N__52224),
            .I(N__52188));
    InMux I__11825 (
            .O(N__52223),
            .I(N__52183));
    InMux I__11824 (
            .O(N__52222),
            .I(N__52179));
    InMux I__11823 (
            .O(N__52221),
            .I(N__52176));
    InMux I__11822 (
            .O(N__52220),
            .I(N__52173));
    LocalMux I__11821 (
            .O(N__52217),
            .I(N__52170));
    InMux I__11820 (
            .O(N__52216),
            .I(N__52167));
    InMux I__11819 (
            .O(N__52215),
            .I(N__52164));
    InMux I__11818 (
            .O(N__52214),
            .I(N__52161));
    InMux I__11817 (
            .O(N__52213),
            .I(N__52158));
    LocalMux I__11816 (
            .O(N__52210),
            .I(N__52153));
    LocalMux I__11815 (
            .O(N__52207),
            .I(N__52153));
    InMux I__11814 (
            .O(N__52206),
            .I(N__52150));
    InMux I__11813 (
            .O(N__52205),
            .I(N__52147));
    InMux I__11812 (
            .O(N__52204),
            .I(N__52142));
    InMux I__11811 (
            .O(N__52203),
            .I(N__52139));
    LocalMux I__11810 (
            .O(N__52200),
            .I(N__52136));
    InMux I__11809 (
            .O(N__52199),
            .I(N__52133));
    InMux I__11808 (
            .O(N__52198),
            .I(N__52130));
    Span4Mux_h I__11807 (
            .O(N__52195),
            .I(N__52125));
    LocalMux I__11806 (
            .O(N__52192),
            .I(N__52125));
    InMux I__11805 (
            .O(N__52191),
            .I(N__52119));
    Span4Mux_v I__11804 (
            .O(N__52188),
            .I(N__52116));
    InMux I__11803 (
            .O(N__52187),
            .I(N__52113));
    InMux I__11802 (
            .O(N__52186),
            .I(N__52110));
    LocalMux I__11801 (
            .O(N__52183),
            .I(N__52107));
    InMux I__11800 (
            .O(N__52182),
            .I(N__52104));
    LocalMux I__11799 (
            .O(N__52179),
            .I(N__52099));
    LocalMux I__11798 (
            .O(N__52176),
            .I(N__52099));
    LocalMux I__11797 (
            .O(N__52173),
            .I(N__52090));
    Span4Mux_h I__11796 (
            .O(N__52170),
            .I(N__52090));
    LocalMux I__11795 (
            .O(N__52167),
            .I(N__52090));
    LocalMux I__11794 (
            .O(N__52164),
            .I(N__52090));
    LocalMux I__11793 (
            .O(N__52161),
            .I(N__52087));
    LocalMux I__11792 (
            .O(N__52158),
            .I(N__52080));
    Span4Mux_v I__11791 (
            .O(N__52153),
            .I(N__52080));
    LocalMux I__11790 (
            .O(N__52150),
            .I(N__52080));
    LocalMux I__11789 (
            .O(N__52147),
            .I(N__52077));
    InMux I__11788 (
            .O(N__52146),
            .I(N__52074));
    InMux I__11787 (
            .O(N__52145),
            .I(N__52071));
    LocalMux I__11786 (
            .O(N__52142),
            .I(N__52066));
    LocalMux I__11785 (
            .O(N__52139),
            .I(N__52066));
    Span4Mux_h I__11784 (
            .O(N__52136),
            .I(N__52061));
    LocalMux I__11783 (
            .O(N__52133),
            .I(N__52061));
    LocalMux I__11782 (
            .O(N__52130),
            .I(N__52058));
    Span4Mux_h I__11781 (
            .O(N__52125),
            .I(N__52055));
    InMux I__11780 (
            .O(N__52124),
            .I(N__52051));
    InMux I__11779 (
            .O(N__52123),
            .I(N__52048));
    InMux I__11778 (
            .O(N__52122),
            .I(N__52045));
    LocalMux I__11777 (
            .O(N__52119),
            .I(N__52038));
    Sp12to4 I__11776 (
            .O(N__52116),
            .I(N__52038));
    LocalMux I__11775 (
            .O(N__52113),
            .I(N__52038));
    LocalMux I__11774 (
            .O(N__52110),
            .I(N__52027));
    Span4Mux_v I__11773 (
            .O(N__52107),
            .I(N__52027));
    LocalMux I__11772 (
            .O(N__52104),
            .I(N__52027));
    Span4Mux_h I__11771 (
            .O(N__52099),
            .I(N__52027));
    Span4Mux_v I__11770 (
            .O(N__52090),
            .I(N__52027));
    Span4Mux_h I__11769 (
            .O(N__52087),
            .I(N__52020));
    Span4Mux_h I__11768 (
            .O(N__52080),
            .I(N__52020));
    Span4Mux_h I__11767 (
            .O(N__52077),
            .I(N__52020));
    LocalMux I__11766 (
            .O(N__52074),
            .I(N__52017));
    LocalMux I__11765 (
            .O(N__52071),
            .I(N__52006));
    Span4Mux_h I__11764 (
            .O(N__52066),
            .I(N__52006));
    Span4Mux_h I__11763 (
            .O(N__52061),
            .I(N__52006));
    Span4Mux_h I__11762 (
            .O(N__52058),
            .I(N__52006));
    Span4Mux_h I__11761 (
            .O(N__52055),
            .I(N__52006));
    InMux I__11760 (
            .O(N__52054),
            .I(N__52003));
    LocalMux I__11759 (
            .O(N__52051),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    LocalMux I__11758 (
            .O(N__52048),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    LocalMux I__11757 (
            .O(N__52045),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    Odrv12 I__11756 (
            .O(N__52038),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    Odrv4 I__11755 (
            .O(N__52027),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    Odrv4 I__11754 (
            .O(N__52020),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    Odrv4 I__11753 (
            .O(N__52017),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    Odrv4 I__11752 (
            .O(N__52006),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    LocalMux I__11751 (
            .O(N__52003),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ));
    InMux I__11750 (
            .O(N__51984),
            .I(N__51981));
    LocalMux I__11749 (
            .O(N__51981),
            .I(N__51978));
    Odrv12 I__11748 (
            .O(N__51978),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_25 ));
    InMux I__11747 (
            .O(N__51975),
            .I(N__51972));
    LocalMux I__11746 (
            .O(N__51972),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_25 ));
    CascadeMux I__11745 (
            .O(N__51969),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_25_cascade_ ));
    InMux I__11744 (
            .O(N__51966),
            .I(N__51963));
    LocalMux I__11743 (
            .O(N__51963),
            .I(N__51960));
    Span4Mux_h I__11742 (
            .O(N__51960),
            .I(N__51957));
    Span4Mux_h I__11741 (
            .O(N__51957),
            .I(N__51954));
    Odrv4 I__11740 (
            .O(N__51954),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_665 ));
    CascadeMux I__11739 (
            .O(N__51951),
            .I(N__51947));
    InMux I__11738 (
            .O(N__51950),
            .I(N__51943));
    InMux I__11737 (
            .O(N__51947),
            .I(N__51940));
    CascadeMux I__11736 (
            .O(N__51946),
            .I(N__51937));
    LocalMux I__11735 (
            .O(N__51943),
            .I(N__51931));
    LocalMux I__11734 (
            .O(N__51940),
            .I(N__51931));
    InMux I__11733 (
            .O(N__51937),
            .I(N__51928));
    InMux I__11732 (
            .O(N__51936),
            .I(N__51916));
    Span4Mux_v I__11731 (
            .O(N__51931),
            .I(N__51910));
    LocalMux I__11730 (
            .O(N__51928),
            .I(N__51910));
    InMux I__11729 (
            .O(N__51927),
            .I(N__51907));
    CascadeMux I__11728 (
            .O(N__51926),
            .I(N__51899));
    InMux I__11727 (
            .O(N__51925),
            .I(N__51896));
    InMux I__11726 (
            .O(N__51924),
            .I(N__51893));
    InMux I__11725 (
            .O(N__51923),
            .I(N__51887));
    InMux I__11724 (
            .O(N__51922),
            .I(N__51884));
    InMux I__11723 (
            .O(N__51921),
            .I(N__51881));
    InMux I__11722 (
            .O(N__51920),
            .I(N__51878));
    InMux I__11721 (
            .O(N__51919),
            .I(N__51875));
    LocalMux I__11720 (
            .O(N__51916),
            .I(N__51872));
    CascadeMux I__11719 (
            .O(N__51915),
            .I(N__51868));
    Span4Mux_h I__11718 (
            .O(N__51910),
            .I(N__51861));
    LocalMux I__11717 (
            .O(N__51907),
            .I(N__51861));
    InMux I__11716 (
            .O(N__51906),
            .I(N__51856));
    CascadeMux I__11715 (
            .O(N__51905),
            .I(N__51853));
    InMux I__11714 (
            .O(N__51904),
            .I(N__51850));
    InMux I__11713 (
            .O(N__51903),
            .I(N__51847));
    InMux I__11712 (
            .O(N__51902),
            .I(N__51843));
    InMux I__11711 (
            .O(N__51899),
            .I(N__51840));
    LocalMux I__11710 (
            .O(N__51896),
            .I(N__51837));
    LocalMux I__11709 (
            .O(N__51893),
            .I(N__51834));
    InMux I__11708 (
            .O(N__51892),
            .I(N__51831));
    InMux I__11707 (
            .O(N__51891),
            .I(N__51828));
    InMux I__11706 (
            .O(N__51890),
            .I(N__51825));
    LocalMux I__11705 (
            .O(N__51887),
            .I(N__51821));
    LocalMux I__11704 (
            .O(N__51884),
            .I(N__51814));
    LocalMux I__11703 (
            .O(N__51881),
            .I(N__51814));
    LocalMux I__11702 (
            .O(N__51878),
            .I(N__51814));
    LocalMux I__11701 (
            .O(N__51875),
            .I(N__51809));
    Span4Mux_h I__11700 (
            .O(N__51872),
            .I(N__51809));
    InMux I__11699 (
            .O(N__51871),
            .I(N__51804));
    InMux I__11698 (
            .O(N__51868),
            .I(N__51804));
    CascadeMux I__11697 (
            .O(N__51867),
            .I(N__51801));
    InMux I__11696 (
            .O(N__51866),
            .I(N__51798));
    Span4Mux_v I__11695 (
            .O(N__51861),
            .I(N__51795));
    InMux I__11694 (
            .O(N__51860),
            .I(N__51792));
    InMux I__11693 (
            .O(N__51859),
            .I(N__51787));
    LocalMux I__11692 (
            .O(N__51856),
            .I(N__51784));
    InMux I__11691 (
            .O(N__51853),
            .I(N__51781));
    LocalMux I__11690 (
            .O(N__51850),
            .I(N__51776));
    LocalMux I__11689 (
            .O(N__51847),
            .I(N__51776));
    InMux I__11688 (
            .O(N__51846),
            .I(N__51773));
    LocalMux I__11687 (
            .O(N__51843),
            .I(N__51770));
    LocalMux I__11686 (
            .O(N__51840),
            .I(N__51765));
    Span4Mux_h I__11685 (
            .O(N__51837),
            .I(N__51765));
    Span4Mux_v I__11684 (
            .O(N__51834),
            .I(N__51760));
    LocalMux I__11683 (
            .O(N__51831),
            .I(N__51760));
    LocalMux I__11682 (
            .O(N__51828),
            .I(N__51755));
    LocalMux I__11681 (
            .O(N__51825),
            .I(N__51755));
    InMux I__11680 (
            .O(N__51824),
            .I(N__51752));
    Span4Mux_h I__11679 (
            .O(N__51821),
            .I(N__51743));
    Span4Mux_v I__11678 (
            .O(N__51814),
            .I(N__51743));
    Span4Mux_h I__11677 (
            .O(N__51809),
            .I(N__51743));
    LocalMux I__11676 (
            .O(N__51804),
            .I(N__51743));
    InMux I__11675 (
            .O(N__51801),
            .I(N__51740));
    LocalMux I__11674 (
            .O(N__51798),
            .I(N__51733));
    Sp12to4 I__11673 (
            .O(N__51795),
            .I(N__51733));
    LocalMux I__11672 (
            .O(N__51792),
            .I(N__51733));
    InMux I__11671 (
            .O(N__51791),
            .I(N__51730));
    InMux I__11670 (
            .O(N__51790),
            .I(N__51727));
    LocalMux I__11669 (
            .O(N__51787),
            .I(N__51718));
    Span4Mux_v I__11668 (
            .O(N__51784),
            .I(N__51718));
    LocalMux I__11667 (
            .O(N__51781),
            .I(N__51718));
    Span4Mux_v I__11666 (
            .O(N__51776),
            .I(N__51718));
    LocalMux I__11665 (
            .O(N__51773),
            .I(N__51707));
    Span4Mux_v I__11664 (
            .O(N__51770),
            .I(N__51707));
    Span4Mux_v I__11663 (
            .O(N__51765),
            .I(N__51707));
    Span4Mux_h I__11662 (
            .O(N__51760),
            .I(N__51707));
    Span4Mux_v I__11661 (
            .O(N__51755),
            .I(N__51707));
    LocalMux I__11660 (
            .O(N__51752),
            .I(N__51702));
    Span4Mux_h I__11659 (
            .O(N__51743),
            .I(N__51702));
    LocalMux I__11658 (
            .O(N__51740),
            .I(N__51697));
    Span12Mux_h I__11657 (
            .O(N__51733),
            .I(N__51697));
    LocalMux I__11656 (
            .O(N__51730),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ));
    LocalMux I__11655 (
            .O(N__51727),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ));
    Odrv4 I__11654 (
            .O(N__51718),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ));
    Odrv4 I__11653 (
            .O(N__51707),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ));
    Odrv4 I__11652 (
            .O(N__51702),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ));
    Odrv12 I__11651 (
            .O(N__51697),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ));
    CascadeMux I__11650 (
            .O(N__51684),
            .I(N__51681));
    InMux I__11649 (
            .O(N__51681),
            .I(N__51678));
    LocalMux I__11648 (
            .O(N__51678),
            .I(N__51675));
    Odrv4 I__11647 (
            .O(N__51675),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_25));
    InMux I__11646 (
            .O(N__51672),
            .I(N__51669));
    LocalMux I__11645 (
            .O(N__51669),
            .I(N__51666));
    Odrv12 I__11644 (
            .O(N__51666),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_25 ));
    InMux I__11643 (
            .O(N__51663),
            .I(N__51660));
    LocalMux I__11642 (
            .O(N__51660),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_25 ));
    InMux I__11641 (
            .O(N__51657),
            .I(N__51653));
    CascadeMux I__11640 (
            .O(N__51656),
            .I(N__51649));
    LocalMux I__11639 (
            .O(N__51653),
            .I(N__51646));
    InMux I__11638 (
            .O(N__51652),
            .I(N__51643));
    InMux I__11637 (
            .O(N__51649),
            .I(N__51640));
    Span4Mux_h I__11636 (
            .O(N__51646),
            .I(N__51637));
    LocalMux I__11635 (
            .O(N__51643),
            .I(N__51634));
    LocalMux I__11634 (
            .O(N__51640),
            .I(N__51631));
    Odrv4 I__11633 (
            .O(N__51637),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_16));
    Odrv4 I__11632 (
            .O(N__51634),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_16));
    Odrv4 I__11631 (
            .O(N__51631),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_16));
    InMux I__11630 (
            .O(N__51624),
            .I(N__51621));
    LocalMux I__11629 (
            .O(N__51621),
            .I(N__51617));
    CascadeMux I__11628 (
            .O(N__51620),
            .I(N__51614));
    Span4Mux_v I__11627 (
            .O(N__51617),
            .I(N__51611));
    InMux I__11626 (
            .O(N__51614),
            .I(N__51607));
    Span4Mux_h I__11625 (
            .O(N__51611),
            .I(N__51604));
    InMux I__11624 (
            .O(N__51610),
            .I(N__51601));
    LocalMux I__11623 (
            .O(N__51607),
            .I(N__51598));
    Span4Mux_h I__11622 (
            .O(N__51604),
            .I(N__51591));
    LocalMux I__11621 (
            .O(N__51601),
            .I(N__51591));
    Span4Mux_h I__11620 (
            .O(N__51598),
            .I(N__51591));
    Odrv4 I__11619 (
            .O(N__51591),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_17));
    CascadeMux I__11618 (
            .O(N__51588),
            .I(N__51583));
    InMux I__11617 (
            .O(N__51587),
            .I(N__51580));
    InMux I__11616 (
            .O(N__51586),
            .I(N__51577));
    InMux I__11615 (
            .O(N__51583),
            .I(N__51574));
    LocalMux I__11614 (
            .O(N__51580),
            .I(N__51571));
    LocalMux I__11613 (
            .O(N__51577),
            .I(N__51568));
    LocalMux I__11612 (
            .O(N__51574),
            .I(N__51565));
    Span4Mux_h I__11611 (
            .O(N__51571),
            .I(N__51562));
    Odrv12 I__11610 (
            .O(N__51568),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_17));
    Odrv4 I__11609 (
            .O(N__51565),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_17));
    Odrv4 I__11608 (
            .O(N__51562),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_17));
    CascadeMux I__11607 (
            .O(N__51555),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_17_cascade_ ));
    InMux I__11606 (
            .O(N__51552),
            .I(N__51549));
    LocalMux I__11605 (
            .O(N__51549),
            .I(N__51546));
    Odrv4 I__11604 (
            .O(N__51546),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_17 ));
    InMux I__11603 (
            .O(N__51543),
            .I(N__51540));
    LocalMux I__11602 (
            .O(N__51540),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_19 ));
    CascadeMux I__11601 (
            .O(N__51537),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HHZ0Z5_cascade_ ));
    InMux I__11600 (
            .O(N__51534),
            .I(N__51531));
    LocalMux I__11599 (
            .O(N__51531),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19 ));
    CascadeMux I__11598 (
            .O(N__51528),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19_cascade_ ));
    InMux I__11597 (
            .O(N__51525),
            .I(N__51522));
    LocalMux I__11596 (
            .O(N__51522),
            .I(N__51519));
    Span4Mux_h I__11595 (
            .O(N__51519),
            .I(N__51516));
    Span4Mux_h I__11594 (
            .O(N__51516),
            .I(N__51513));
    Odrv4 I__11593 (
            .O(N__51513),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_19 ));
    InMux I__11592 (
            .O(N__51510),
            .I(N__51507));
    LocalMux I__11591 (
            .O(N__51507),
            .I(N__51502));
    CascadeMux I__11590 (
            .O(N__51506),
            .I(N__51499));
    CascadeMux I__11589 (
            .O(N__51505),
            .I(N__51496));
    Span4Mux_v I__11588 (
            .O(N__51502),
            .I(N__51493));
    InMux I__11587 (
            .O(N__51499),
            .I(N__51490));
    InMux I__11586 (
            .O(N__51496),
            .I(N__51487));
    Span4Mux_h I__11585 (
            .O(N__51493),
            .I(N__51482));
    LocalMux I__11584 (
            .O(N__51490),
            .I(N__51482));
    LocalMux I__11583 (
            .O(N__51487),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_19));
    Odrv4 I__11582 (
            .O(N__51482),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_19));
    InMux I__11581 (
            .O(N__51477),
            .I(N__51473));
    InMux I__11580 (
            .O(N__51476),
            .I(N__51470));
    LocalMux I__11579 (
            .O(N__51473),
            .I(N__51467));
    LocalMux I__11578 (
            .O(N__51470),
            .I(N__51464));
    Span4Mux_h I__11577 (
            .O(N__51467),
            .I(N__51460));
    Span4Mux_h I__11576 (
            .O(N__51464),
            .I(N__51457));
    InMux I__11575 (
            .O(N__51463),
            .I(N__51454));
    Odrv4 I__11574 (
            .O(N__51460),
            .I(cemf_module_64ch_ctrl_inst1_data_config_19));
    Odrv4 I__11573 (
            .O(N__51457),
            .I(cemf_module_64ch_ctrl_inst1_data_config_19));
    LocalMux I__11572 (
            .O(N__51454),
            .I(cemf_module_64ch_ctrl_inst1_data_config_19));
    CascadeMux I__11571 (
            .O(N__51447),
            .I(N__51444));
    InMux I__11570 (
            .O(N__51444),
            .I(N__51441));
    LocalMux I__11569 (
            .O(N__51441),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_19 ));
    InMux I__11568 (
            .O(N__51438),
            .I(N__51435));
    LocalMux I__11567 (
            .O(N__51435),
            .I(N__51431));
    CascadeMux I__11566 (
            .O(N__51434),
            .I(N__51427));
    Span4Mux_h I__11565 (
            .O(N__51431),
            .I(N__51424));
    CascadeMux I__11564 (
            .O(N__51430),
            .I(N__51421));
    InMux I__11563 (
            .O(N__51427),
            .I(N__51418));
    Span4Mux_h I__11562 (
            .O(N__51424),
            .I(N__51415));
    InMux I__11561 (
            .O(N__51421),
            .I(N__51412));
    LocalMux I__11560 (
            .O(N__51418),
            .I(N__51409));
    Odrv4 I__11559 (
            .O(N__51415),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_18));
    LocalMux I__11558 (
            .O(N__51412),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_18));
    Odrv4 I__11557 (
            .O(N__51409),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_18));
    InMux I__11556 (
            .O(N__51402),
            .I(N__51399));
    LocalMux I__11555 (
            .O(N__51399),
            .I(N__51396));
    Span4Mux_v I__11554 (
            .O(N__51396),
            .I(N__51392));
    InMux I__11553 (
            .O(N__51395),
            .I(N__51389));
    Span4Mux_h I__11552 (
            .O(N__51392),
            .I(N__51386));
    LocalMux I__11551 (
            .O(N__51389),
            .I(N__51383));
    Span4Mux_h I__11550 (
            .O(N__51386),
            .I(N__51377));
    Span4Mux_v I__11549 (
            .O(N__51383),
            .I(N__51377));
    InMux I__11548 (
            .O(N__51382),
            .I(N__51374));
    Odrv4 I__11547 (
            .O(N__51377),
            .I(cemf_module_64ch_ctrl_inst1_data_config_18));
    LocalMux I__11546 (
            .O(N__51374),
            .I(cemf_module_64ch_ctrl_inst1_data_config_18));
    InMux I__11545 (
            .O(N__51369),
            .I(N__51365));
    InMux I__11544 (
            .O(N__51368),
            .I(N__51361));
    LocalMux I__11543 (
            .O(N__51365),
            .I(N__51358));
    InMux I__11542 (
            .O(N__51364),
            .I(N__51355));
    LocalMux I__11541 (
            .O(N__51361),
            .I(N__51352));
    Span4Mux_v I__11540 (
            .O(N__51358),
            .I(N__51347));
    LocalMux I__11539 (
            .O(N__51355),
            .I(N__51347));
    Odrv4 I__11538 (
            .O(N__51352),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_18));
    Odrv4 I__11537 (
            .O(N__51347),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_18));
    CascadeMux I__11536 (
            .O(N__51342),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_18_cascade_ ));
    InMux I__11535 (
            .O(N__51339),
            .I(N__51336));
    LocalMux I__11534 (
            .O(N__51336),
            .I(N__51333));
    Span4Mux_h I__11533 (
            .O(N__51333),
            .I(N__51330));
    Odrv4 I__11532 (
            .O(N__51330),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_18 ));
    CascadeMux I__11531 (
            .O(N__51327),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGHZ0Z5_cascade_ ));
    InMux I__11530 (
            .O(N__51324),
            .I(N__51321));
    LocalMux I__11529 (
            .O(N__51321),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18 ));
    CascadeMux I__11528 (
            .O(N__51318),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18_cascade_ ));
    InMux I__11527 (
            .O(N__51315),
            .I(N__51312));
    LocalMux I__11526 (
            .O(N__51312),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_18 ));
    InMux I__11525 (
            .O(N__51309),
            .I(N__51306));
    LocalMux I__11524 (
            .O(N__51306),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_1 ));
    InMux I__11523 (
            .O(N__51303),
            .I(N__51300));
    LocalMux I__11522 (
            .O(N__51300),
            .I(N__51296));
    InMux I__11521 (
            .O(N__51299),
            .I(N__51293));
    Span12Mux_v I__11520 (
            .O(N__51296),
            .I(N__51290));
    LocalMux I__11519 (
            .O(N__51293),
            .I(\I2C_top_level_inst1.s_r_w ));
    Odrv12 I__11518 (
            .O(N__51290),
            .I(\I2C_top_level_inst1.s_r_w ));
    InMux I__11517 (
            .O(N__51285),
            .I(N__51282));
    LocalMux I__11516 (
            .O(N__51282),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_0 ));
    InMux I__11515 (
            .O(N__51279),
            .I(N__51276));
    LocalMux I__11514 (
            .O(N__51276),
            .I(N__51273));
    Span4Mux_v I__11513 (
            .O(N__51273),
            .I(N__51270));
    Span4Mux_h I__11512 (
            .O(N__51270),
            .I(N__51267));
    Odrv4 I__11511 (
            .O(N__51267),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_27));
    InMux I__11510 (
            .O(N__51264),
            .I(N__51261));
    LocalMux I__11509 (
            .O(N__51261),
            .I(N__51258));
    Span4Mux_h I__11508 (
            .O(N__51258),
            .I(N__51255));
    Odrv4 I__11507 (
            .O(N__51255),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_29));
    InMux I__11506 (
            .O(N__51252),
            .I(N__51248));
    InMux I__11505 (
            .O(N__51251),
            .I(N__51245));
    LocalMux I__11504 (
            .O(N__51248),
            .I(N__51242));
    LocalMux I__11503 (
            .O(N__51245),
            .I(N__51238));
    Span4Mux_v I__11502 (
            .O(N__51242),
            .I(N__51235));
    InMux I__11501 (
            .O(N__51241),
            .I(N__51232));
    Span4Mux_v I__11500 (
            .O(N__51238),
            .I(N__51229));
    Span4Mux_h I__11499 (
            .O(N__51235),
            .I(N__51224));
    LocalMux I__11498 (
            .O(N__51232),
            .I(N__51224));
    Span4Mux_h I__11497 (
            .O(N__51229),
            .I(N__51221));
    Span4Mux_v I__11496 (
            .O(N__51224),
            .I(N__51218));
    Odrv4 I__11495 (
            .O(N__51221),
            .I(cemf_module_64ch_ctrl_inst1_data_config_23));
    Odrv4 I__11494 (
            .O(N__51218),
            .I(cemf_module_64ch_ctrl_inst1_data_config_23));
    InMux I__11493 (
            .O(N__51213),
            .I(N__51210));
    LocalMux I__11492 (
            .O(N__51210),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_1 ));
    IoInMux I__11491 (
            .O(N__51207),
            .I(N__51203));
    InMux I__11490 (
            .O(N__51206),
            .I(N__51200));
    LocalMux I__11489 (
            .O(N__51203),
            .I(N__51197));
    LocalMux I__11488 (
            .O(N__51200),
            .I(N__51194));
    IoSpan4Mux I__11487 (
            .O(N__51197),
            .I(N__51191));
    Span4Mux_h I__11486 (
            .O(N__51194),
            .I(N__51187));
    Span4Mux_s2_v I__11485 (
            .O(N__51191),
            .I(N__51183));
    InMux I__11484 (
            .O(N__51190),
            .I(N__51180));
    Span4Mux_v I__11483 (
            .O(N__51187),
            .I(N__51177));
    InMux I__11482 (
            .O(N__51186),
            .I(N__51174));
    Sp12to4 I__11481 (
            .O(N__51183),
            .I(N__51171));
    LocalMux I__11480 (
            .O(N__51180),
            .I(N__51168));
    Span4Mux_h I__11479 (
            .O(N__51177),
            .I(N__51163));
    LocalMux I__11478 (
            .O(N__51174),
            .I(N__51163));
    Span12Mux_h I__11477 (
            .O(N__51171),
            .I(N__51160));
    Span4Mux_v I__11476 (
            .O(N__51168),
            .I(N__51157));
    Span4Mux_h I__11475 (
            .O(N__51163),
            .I(N__51154));
    Span12Mux_v I__11474 (
            .O(N__51160),
            .I(N__51151));
    Span4Mux_h I__11473 (
            .O(N__51157),
            .I(N__51148));
    Span4Mux_v I__11472 (
            .O(N__51154),
            .I(N__51145));
    Span12Mux_v I__11471 (
            .O(N__51151),
            .I(N__51142));
    Sp12to4 I__11470 (
            .O(N__51148),
            .I(N__51139));
    IoSpan4Mux I__11469 (
            .O(N__51145),
            .I(N__51136));
    Odrv12 I__11468 (
            .O(N__51142),
            .I(scl_c));
    Odrv12 I__11467 (
            .O(N__51139),
            .I(scl_c));
    Odrv4 I__11466 (
            .O(N__51136),
            .I(scl_c));
    InMux I__11465 (
            .O(N__51129),
            .I(N__51126));
    LocalMux I__11464 (
            .O(N__51126),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_0 ));
    InMux I__11463 (
            .O(N__51123),
            .I(N__51113));
    InMux I__11462 (
            .O(N__51122),
            .I(N__51113));
    InMux I__11461 (
            .O(N__51121),
            .I(N__51104));
    InMux I__11460 (
            .O(N__51120),
            .I(N__51104));
    InMux I__11459 (
            .O(N__51119),
            .I(N__51104));
    InMux I__11458 (
            .O(N__51118),
            .I(N__51104));
    LocalMux I__11457 (
            .O(N__51113),
            .I(N__51101));
    LocalMux I__11456 (
            .O(N__51104),
            .I(N__51098));
    Span4Mux_v I__11455 (
            .O(N__51101),
            .I(N__51095));
    Span4Mux_v I__11454 (
            .O(N__51098),
            .I(N__51092));
    Span4Mux_h I__11453 (
            .O(N__51095),
            .I(N__51089));
    Span4Mux_h I__11452 (
            .O(N__51092),
            .I(N__51086));
    Odrv4 I__11451 (
            .O(N__51089),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0 ));
    Odrv4 I__11450 (
            .O(N__51086),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0 ));
    InMux I__11449 (
            .O(N__51081),
            .I(N__51070));
    InMux I__11448 (
            .O(N__51080),
            .I(N__51070));
    InMux I__11447 (
            .O(N__51079),
            .I(N__51059));
    InMux I__11446 (
            .O(N__51078),
            .I(N__51059));
    InMux I__11445 (
            .O(N__51077),
            .I(N__51059));
    InMux I__11444 (
            .O(N__51076),
            .I(N__51059));
    InMux I__11443 (
            .O(N__51075),
            .I(N__51059));
    LocalMux I__11442 (
            .O(N__51070),
            .I(\I2C_top_level_inst1.s_command_1 ));
    LocalMux I__11441 (
            .O(N__51059),
            .I(\I2C_top_level_inst1.s_command_1 ));
    CascadeMux I__11440 (
            .O(N__51054),
            .I(N__51049));
    CascadeMux I__11439 (
            .O(N__51053),
            .I(N__51045));
    InMux I__11438 (
            .O(N__51052),
            .I(N__51037));
    InMux I__11437 (
            .O(N__51049),
            .I(N__51037));
    InMux I__11436 (
            .O(N__51048),
            .I(N__51037));
    InMux I__11435 (
            .O(N__51045),
            .I(N__51032));
    InMux I__11434 (
            .O(N__51044),
            .I(N__51032));
    LocalMux I__11433 (
            .O(N__51037),
            .I(N__51029));
    LocalMux I__11432 (
            .O(N__51032),
            .I(\I2C_top_level_inst1.s_command_2 ));
    Odrv4 I__11431 (
            .O(N__51029),
            .I(\I2C_top_level_inst1.s_command_2 ));
    CascadeMux I__11430 (
            .O(N__51024),
            .I(N__51019));
    CascadeMux I__11429 (
            .O(N__51023),
            .I(N__51016));
    InMux I__11428 (
            .O(N__51022),
            .I(N__51008));
    InMux I__11427 (
            .O(N__51019),
            .I(N__51008));
    InMux I__11426 (
            .O(N__51016),
            .I(N__50999));
    InMux I__11425 (
            .O(N__51015),
            .I(N__50999));
    InMux I__11424 (
            .O(N__51014),
            .I(N__50999));
    InMux I__11423 (
            .O(N__51013),
            .I(N__50999));
    LocalMux I__11422 (
            .O(N__51008),
            .I(\I2C_top_level_inst1.s_command_3 ));
    LocalMux I__11421 (
            .O(N__50999),
            .I(\I2C_top_level_inst1.s_command_3 ));
    InMux I__11420 (
            .O(N__50994),
            .I(N__50990));
    InMux I__11419 (
            .O(N__50993),
            .I(N__50987));
    LocalMux I__11418 (
            .O(N__50990),
            .I(N__50984));
    LocalMux I__11417 (
            .O(N__50987),
            .I(N__50980));
    Span4Mux_h I__11416 (
            .O(N__50984),
            .I(N__50976));
    InMux I__11415 (
            .O(N__50983),
            .I(N__50973));
    Span4Mux_h I__11414 (
            .O(N__50980),
            .I(N__50970));
    InMux I__11413 (
            .O(N__50979),
            .I(N__50967));
    Span4Mux_v I__11412 (
            .O(N__50976),
            .I(N__50960));
    LocalMux I__11411 (
            .O(N__50973),
            .I(N__50960));
    Span4Mux_v I__11410 (
            .O(N__50970),
            .I(N__50960));
    LocalMux I__11409 (
            .O(N__50967),
            .I(\I2C_top_level_inst1.s_load_wdata ));
    Odrv4 I__11408 (
            .O(N__50960),
            .I(\I2C_top_level_inst1.s_load_wdata ));
    InMux I__11407 (
            .O(N__50955),
            .I(N__50952));
    LocalMux I__11406 (
            .O(N__50952),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_0 ));
    InMux I__11405 (
            .O(N__50949),
            .I(N__50946));
    LocalMux I__11404 (
            .O(N__50946),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_1 ));
    InMux I__11403 (
            .O(N__50943),
            .I(N__50940));
    LocalMux I__11402 (
            .O(N__50940),
            .I(N__50937));
    Span4Mux_v I__11401 (
            .O(N__50937),
            .I(N__50934));
    Span4Mux_v I__11400 (
            .O(N__50934),
            .I(N__50927));
    InMux I__11399 (
            .O(N__50933),
            .I(N__50924));
    InMux I__11398 (
            .O(N__50932),
            .I(N__50914));
    InMux I__11397 (
            .O(N__50931),
            .I(N__50914));
    InMux I__11396 (
            .O(N__50930),
            .I(N__50914));
    Span4Mux_h I__11395 (
            .O(N__50927),
            .I(N__50909));
    LocalMux I__11394 (
            .O(N__50924),
            .I(N__50909));
    InMux I__11393 (
            .O(N__50923),
            .I(N__50902));
    InMux I__11392 (
            .O(N__50922),
            .I(N__50902));
    InMux I__11391 (
            .O(N__50921),
            .I(N__50902));
    LocalMux I__11390 (
            .O(N__50914),
            .I(N__50899));
    Span4Mux_h I__11389 (
            .O(N__50909),
            .I(N__50896));
    LocalMux I__11388 (
            .O(N__50902),
            .I(N__50893));
    Odrv4 I__11387 (
            .O(N__50899),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2 ));
    Odrv4 I__11386 (
            .O(N__50896),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2 ));
    Odrv4 I__11385 (
            .O(N__50893),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2 ));
    InMux I__11384 (
            .O(N__50886),
            .I(N__50878));
    CascadeMux I__11383 (
            .O(N__50885),
            .I(N__50875));
    InMux I__11382 (
            .O(N__50884),
            .I(N__50866));
    InMux I__11381 (
            .O(N__50883),
            .I(N__50866));
    InMux I__11380 (
            .O(N__50882),
            .I(N__50861));
    InMux I__11379 (
            .O(N__50881),
            .I(N__50858));
    LocalMux I__11378 (
            .O(N__50878),
            .I(N__50855));
    InMux I__11377 (
            .O(N__50875),
            .I(N__50844));
    InMux I__11376 (
            .O(N__50874),
            .I(N__50844));
    InMux I__11375 (
            .O(N__50873),
            .I(N__50844));
    InMux I__11374 (
            .O(N__50872),
            .I(N__50844));
    InMux I__11373 (
            .O(N__50871),
            .I(N__50844));
    LocalMux I__11372 (
            .O(N__50866),
            .I(N__50841));
    InMux I__11371 (
            .O(N__50865),
            .I(N__50836));
    InMux I__11370 (
            .O(N__50864),
            .I(N__50836));
    LocalMux I__11369 (
            .O(N__50861),
            .I(N__50833));
    LocalMux I__11368 (
            .O(N__50858),
            .I(N__50830));
    Span4Mux_h I__11367 (
            .O(N__50855),
            .I(N__50821));
    LocalMux I__11366 (
            .O(N__50844),
            .I(N__50821));
    Span4Mux_v I__11365 (
            .O(N__50841),
            .I(N__50821));
    LocalMux I__11364 (
            .O(N__50836),
            .I(N__50821));
    Span4Mux_v I__11363 (
            .O(N__50833),
            .I(N__50817));
    Span4Mux_h I__11362 (
            .O(N__50830),
            .I(N__50814));
    Span4Mux_h I__11361 (
            .O(N__50821),
            .I(N__50811));
    InMux I__11360 (
            .O(N__50820),
            .I(N__50808));
    Sp12to4 I__11359 (
            .O(N__50817),
            .I(N__50805));
    Span4Mux_v I__11358 (
            .O(N__50814),
            .I(N__50802));
    Span4Mux_v I__11357 (
            .O(N__50811),
            .I(N__50797));
    LocalMux I__11356 (
            .O(N__50808),
            .I(N__50797));
    Odrv12 I__11355 (
            .O(N__50805),
            .I(\I2C_top_level_inst1.s_start ));
    Odrv4 I__11354 (
            .O(N__50802),
            .I(\I2C_top_level_inst1.s_start ));
    Odrv4 I__11353 (
            .O(N__50797),
            .I(\I2C_top_level_inst1.s_start ));
    InMux I__11352 (
            .O(N__50790),
            .I(N__50787));
    LocalMux I__11351 (
            .O(N__50787),
            .I(N__50784));
    Span4Mux_h I__11350 (
            .O(N__50784),
            .I(N__50781));
    Span4Mux_h I__11349 (
            .O(N__50781),
            .I(N__50778));
    Odrv4 I__11348 (
            .O(N__50778),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_0 ));
    CascadeMux I__11347 (
            .O(N__50775),
            .I(N__50772));
    InMux I__11346 (
            .O(N__50772),
            .I(N__50769));
    LocalMux I__11345 (
            .O(N__50769),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_86_0 ));
    InMux I__11344 (
            .O(N__50766),
            .I(N__50763));
    LocalMux I__11343 (
            .O(N__50763),
            .I(N__50760));
    Odrv4 I__11342 (
            .O(N__50760),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_95_0 ));
    InMux I__11341 (
            .O(N__50757),
            .I(N__50754));
    LocalMux I__11340 (
            .O(N__50754),
            .I(N__50751));
    Span4Mux_h I__11339 (
            .O(N__50751),
            .I(N__50748));
    Span4Mux_h I__11338 (
            .O(N__50748),
            .I(N__50743));
    InMux I__11337 (
            .O(N__50747),
            .I(N__50738));
    InMux I__11336 (
            .O(N__50746),
            .I(N__50738));
    Span4Mux_h I__11335 (
            .O(N__50743),
            .I(N__50735));
    LocalMux I__11334 (
            .O(N__50738),
            .I(N__50732));
    Odrv4 I__11333 (
            .O(N__50735),
            .I(\I2C_top_level_inst1.s_stop ));
    Odrv4 I__11332 (
            .O(N__50732),
            .I(\I2C_top_level_inst1.s_stop ));
    InMux I__11331 (
            .O(N__50727),
            .I(N__50724));
    LocalMux I__11330 (
            .O(N__50724),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_0 ));
    InMux I__11329 (
            .O(N__50721),
            .I(N__50718));
    LocalMux I__11328 (
            .O(N__50718),
            .I(N__50711));
    InMux I__11327 (
            .O(N__50717),
            .I(N__50706));
    InMux I__11326 (
            .O(N__50716),
            .I(N__50706));
    InMux I__11325 (
            .O(N__50715),
            .I(N__50701));
    InMux I__11324 (
            .O(N__50714),
            .I(N__50701));
    Span4Mux_v I__11323 (
            .O(N__50711),
            .I(N__50698));
    LocalMux I__11322 (
            .O(N__50706),
            .I(N__50693));
    LocalMux I__11321 (
            .O(N__50701),
            .I(N__50693));
    Span4Mux_h I__11320 (
            .O(N__50698),
            .I(N__50690));
    Span12Mux_v I__11319 (
            .O(N__50693),
            .I(N__50687));
    Odrv4 I__11318 (
            .O(N__50690),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2 ));
    Odrv12 I__11317 (
            .O(N__50687),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2 ));
    InMux I__11316 (
            .O(N__50682),
            .I(N__50678));
    InMux I__11315 (
            .O(N__50681),
            .I(N__50675));
    LocalMux I__11314 (
            .O(N__50678),
            .I(N__50670));
    LocalMux I__11313 (
            .O(N__50675),
            .I(N__50670));
    Odrv4 I__11312 (
            .O(N__50670),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_844_2 ));
    InMux I__11311 (
            .O(N__50667),
            .I(N__50663));
    InMux I__11310 (
            .O(N__50666),
            .I(N__50660));
    LocalMux I__11309 (
            .O(N__50663),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2 ));
    LocalMux I__11308 (
            .O(N__50660),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2 ));
    InMux I__11307 (
            .O(N__50655),
            .I(N__50652));
    LocalMux I__11306 (
            .O(N__50652),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_1 ));
    InMux I__11305 (
            .O(N__50649),
            .I(N__50646));
    LocalMux I__11304 (
            .O(N__50646),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_1 ));
    InMux I__11303 (
            .O(N__50643),
            .I(N__50637));
    InMux I__11302 (
            .O(N__50642),
            .I(N__50637));
    LocalMux I__11301 (
            .O(N__50637),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1754_1 ));
    CascadeMux I__11300 (
            .O(N__50634),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0_cascade_ ));
    InMux I__11299 (
            .O(N__50631),
            .I(N__50628));
    LocalMux I__11298 (
            .O(N__50628),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_25 ));
    CascadeMux I__11297 (
            .O(N__50625),
            .I(N__50622));
    InMux I__11296 (
            .O(N__50622),
            .I(N__50618));
    InMux I__11295 (
            .O(N__50621),
            .I(N__50615));
    LocalMux I__11294 (
            .O(N__50618),
            .I(N__50612));
    LocalMux I__11293 (
            .O(N__50615),
            .I(N__50608));
    Span4Mux_h I__11292 (
            .O(N__50612),
            .I(N__50605));
    InMux I__11291 (
            .O(N__50611),
            .I(N__50602));
    Span4Mux_v I__11290 (
            .O(N__50608),
            .I(N__50597));
    Span4Mux_h I__11289 (
            .O(N__50605),
            .I(N__50597));
    LocalMux I__11288 (
            .O(N__50602),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2 ));
    Odrv4 I__11287 (
            .O(N__50597),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2 ));
    InMux I__11286 (
            .O(N__50592),
            .I(N__50589));
    LocalMux I__11285 (
            .O(N__50589),
            .I(N__50586));
    Span4Mux_h I__11284 (
            .O(N__50586),
            .I(N__50582));
    InMux I__11283 (
            .O(N__50585),
            .I(N__50578));
    Span4Mux_v I__11282 (
            .O(N__50582),
            .I(N__50575));
    InMux I__11281 (
            .O(N__50581),
            .I(N__50572));
    LocalMux I__11280 (
            .O(N__50578),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i ));
    Odrv4 I__11279 (
            .O(N__50575),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i ));
    LocalMux I__11278 (
            .O(N__50572),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i ));
    CascadeMux I__11277 (
            .O(N__50565),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_24_cascade_ ));
    CascadeMux I__11276 (
            .O(N__50562),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_11_cascade_ ));
    InMux I__11275 (
            .O(N__50559),
            .I(N__50555));
    InMux I__11274 (
            .O(N__50558),
            .I(N__50552));
    LocalMux I__11273 (
            .O(N__50555),
            .I(N__50546));
    LocalMux I__11272 (
            .O(N__50552),
            .I(N__50546));
    InMux I__11271 (
            .O(N__50551),
            .I(N__50540));
    Span4Mux_v I__11270 (
            .O(N__50546),
            .I(N__50533));
    InMux I__11269 (
            .O(N__50545),
            .I(N__50530));
    InMux I__11268 (
            .O(N__50544),
            .I(N__50525));
    InMux I__11267 (
            .O(N__50543),
            .I(N__50525));
    LocalMux I__11266 (
            .O(N__50540),
            .I(N__50522));
    InMux I__11265 (
            .O(N__50539),
            .I(N__50517));
    InMux I__11264 (
            .O(N__50538),
            .I(N__50517));
    InMux I__11263 (
            .O(N__50537),
            .I(N__50512));
    InMux I__11262 (
            .O(N__50536),
            .I(N__50512));
    Span4Mux_h I__11261 (
            .O(N__50533),
            .I(N__50509));
    LocalMux I__11260 (
            .O(N__50530),
            .I(N__50506));
    LocalMux I__11259 (
            .O(N__50525),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ));
    Odrv4 I__11258 (
            .O(N__50522),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ));
    LocalMux I__11257 (
            .O(N__50517),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ));
    LocalMux I__11256 (
            .O(N__50512),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ));
    Odrv4 I__11255 (
            .O(N__50509),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ));
    Odrv12 I__11254 (
            .O(N__50506),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ));
    CascadeMux I__11253 (
            .O(N__50493),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_11_cascade_ ));
    CascadeMux I__11252 (
            .O(N__50490),
            .I(N__50487));
    InMux I__11251 (
            .O(N__50487),
            .I(N__50484));
    LocalMux I__11250 (
            .O(N__50484),
            .I(N__50481));
    Span4Mux_v I__11249 (
            .O(N__50481),
            .I(N__50478));
    Span4Mux_h I__11248 (
            .O(N__50478),
            .I(N__50475));
    Span4Mux_h I__11247 (
            .O(N__50475),
            .I(N__50472));
    Odrv4 I__11246 (
            .O(N__50472),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_2_11 ));
    CascadeMux I__11245 (
            .O(N__50469),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_1_2_0_cascade_ ));
    CascadeMux I__11244 (
            .O(N__50466),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i_cascade_ ));
    CascadeMux I__11243 (
            .O(N__50463),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_372_cascade_ ));
    InMux I__11242 (
            .O(N__50460),
            .I(N__50457));
    LocalMux I__11241 (
            .O(N__50457),
            .I(N__50453));
    InMux I__11240 (
            .O(N__50456),
            .I(N__50450));
    Span4Mux_h I__11239 (
            .O(N__50453),
            .I(N__50446));
    LocalMux I__11238 (
            .O(N__50450),
            .I(N__50443));
    InMux I__11237 (
            .O(N__50449),
            .I(N__50440));
    Span4Mux_h I__11236 (
            .O(N__50446),
            .I(N__50437));
    Span12Mux_h I__11235 (
            .O(N__50443),
            .I(N__50434));
    LocalMux I__11234 (
            .O(N__50440),
            .I(N_409));
    Odrv4 I__11233 (
            .O(N__50437),
            .I(N_409));
    Odrv12 I__11232 (
            .O(N__50434),
            .I(N_409));
    InMux I__11231 (
            .O(N__50427),
            .I(N__50424));
    LocalMux I__11230 (
            .O(N__50424),
            .I(N__50421));
    Odrv4 I__11229 (
            .O(N__50421),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_a3_1_0_14 ));
    CascadeMux I__11228 (
            .O(N__50418),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_412_0_cascade_ ));
    InMux I__11227 (
            .O(N__50415),
            .I(N__50412));
    LocalMux I__11226 (
            .O(N__50412),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_1_14 ));
    CascadeMux I__11225 (
            .O(N__50409),
            .I(N__50398));
    InMux I__11224 (
            .O(N__50408),
            .I(N__50381));
    InMux I__11223 (
            .O(N__50407),
            .I(N__50381));
    InMux I__11222 (
            .O(N__50406),
            .I(N__50368));
    InMux I__11221 (
            .O(N__50405),
            .I(N__50368));
    InMux I__11220 (
            .O(N__50404),
            .I(N__50368));
    InMux I__11219 (
            .O(N__50403),
            .I(N__50368));
    InMux I__11218 (
            .O(N__50402),
            .I(N__50368));
    InMux I__11217 (
            .O(N__50401),
            .I(N__50359));
    InMux I__11216 (
            .O(N__50398),
            .I(N__50359));
    InMux I__11215 (
            .O(N__50397),
            .I(N__50359));
    InMux I__11214 (
            .O(N__50396),
            .I(N__50359));
    CascadeMux I__11213 (
            .O(N__50395),
            .I(N__50356));
    InMux I__11212 (
            .O(N__50394),
            .I(N__50334));
    InMux I__11211 (
            .O(N__50393),
            .I(N__50334));
    InMux I__11210 (
            .O(N__50392),
            .I(N__50334));
    InMux I__11209 (
            .O(N__50391),
            .I(N__50334));
    InMux I__11208 (
            .O(N__50390),
            .I(N__50334));
    InMux I__11207 (
            .O(N__50389),
            .I(N__50334));
    InMux I__11206 (
            .O(N__50388),
            .I(N__50329));
    InMux I__11205 (
            .O(N__50387),
            .I(N__50329));
    CascadeMux I__11204 (
            .O(N__50386),
            .I(N__50326));
    LocalMux I__11203 (
            .O(N__50381),
            .I(N__50323));
    InMux I__11202 (
            .O(N__50380),
            .I(N__50318));
    InMux I__11201 (
            .O(N__50379),
            .I(N__50318));
    LocalMux I__11200 (
            .O(N__50368),
            .I(N__50313));
    LocalMux I__11199 (
            .O(N__50359),
            .I(N__50313));
    InMux I__11198 (
            .O(N__50356),
            .I(N__50308));
    InMux I__11197 (
            .O(N__50355),
            .I(N__50308));
    InMux I__11196 (
            .O(N__50354),
            .I(N__50301));
    InMux I__11195 (
            .O(N__50353),
            .I(N__50301));
    InMux I__11194 (
            .O(N__50352),
            .I(N__50301));
    InMux I__11193 (
            .O(N__50351),
            .I(N__50290));
    InMux I__11192 (
            .O(N__50350),
            .I(N__50290));
    InMux I__11191 (
            .O(N__50349),
            .I(N__50290));
    InMux I__11190 (
            .O(N__50348),
            .I(N__50290));
    InMux I__11189 (
            .O(N__50347),
            .I(N__50290));
    LocalMux I__11188 (
            .O(N__50334),
            .I(N__50285));
    LocalMux I__11187 (
            .O(N__50329),
            .I(N__50285));
    InMux I__11186 (
            .O(N__50326),
            .I(N__50282));
    Span4Mux_v I__11185 (
            .O(N__50323),
            .I(N__50277));
    LocalMux I__11184 (
            .O(N__50318),
            .I(N__50277));
    Span4Mux_h I__11183 (
            .O(N__50313),
            .I(N__50274));
    LocalMux I__11182 (
            .O(N__50308),
            .I(N__50265));
    LocalMux I__11181 (
            .O(N__50301),
            .I(N__50265));
    LocalMux I__11180 (
            .O(N__50290),
            .I(N__50265));
    Span4Mux_v I__11179 (
            .O(N__50285),
            .I(N__50265));
    LocalMux I__11178 (
            .O(N__50282),
            .I(N__50262));
    Span4Mux_h I__11177 (
            .O(N__50277),
            .I(N__50257));
    Span4Mux_v I__11176 (
            .O(N__50274),
            .I(N__50257));
    Span4Mux_h I__11175 (
            .O(N__50265),
            .I(N__50254));
    Span4Mux_h I__11174 (
            .O(N__50262),
            .I(N__50251));
    Span4Mux_v I__11173 (
            .O(N__50257),
            .I(N__50248));
    Span4Mux_v I__11172 (
            .O(N__50254),
            .I(N__50245));
    Span4Mux_h I__11171 (
            .O(N__50251),
            .I(N__50239));
    Span4Mux_h I__11170 (
            .O(N__50248),
            .I(N__50239));
    Span4Mux_h I__11169 (
            .O(N__50245),
            .I(N__50236));
    InMux I__11168 (
            .O(N__50244),
            .I(N__50233));
    Odrv4 I__11167 (
            .O(N__50239),
            .I(N_410));
    Odrv4 I__11166 (
            .O(N__50236),
            .I(N_410));
    LocalMux I__11165 (
            .O(N__50233),
            .I(N_410));
    InMux I__11164 (
            .O(N__50226),
            .I(N__50223));
    LocalMux I__11163 (
            .O(N__50223),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_1_0_14 ));
    CascadeMux I__11162 (
            .O(N__50220),
            .I(N__50215));
    InMux I__11161 (
            .O(N__50219),
            .I(N__50208));
    InMux I__11160 (
            .O(N__50218),
            .I(N__50208));
    InMux I__11159 (
            .O(N__50215),
            .I(N__50208));
    LocalMux I__11158 (
            .O(N__50208),
            .I(N__50205));
    Span4Mux_v I__11157 (
            .O(N__50205),
            .I(N__50202));
    Span4Mux_h I__11156 (
            .O(N__50202),
            .I(N__50199));
    Odrv4 I__11155 (
            .O(N__50199),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_322 ));
    CascadeMux I__11154 (
            .O(N__50196),
            .I(N__50193));
    InMux I__11153 (
            .O(N__50193),
            .I(N__50188));
    InMux I__11152 (
            .O(N__50192),
            .I(N__50185));
    InMux I__11151 (
            .O(N__50191),
            .I(N__50182));
    LocalMux I__11150 (
            .O(N__50188),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0 ));
    LocalMux I__11149 (
            .O(N__50185),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0 ));
    LocalMux I__11148 (
            .O(N__50182),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0 ));
    InMux I__11147 (
            .O(N__50175),
            .I(N__50172));
    LocalMux I__11146 (
            .O(N__50172),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0 ));
    CascadeMux I__11145 (
            .O(N__50169),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0_cascade_ ));
    InMux I__11144 (
            .O(N__50166),
            .I(N__50163));
    LocalMux I__11143 (
            .O(N__50163),
            .I(N__50160));
    Span4Mux_v I__11142 (
            .O(N__50160),
            .I(N__50157));
    Odrv4 I__11141 (
            .O(N__50157),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_267 ));
    InMux I__11140 (
            .O(N__50154),
            .I(N__50151));
    LocalMux I__11139 (
            .O(N__50151),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_394 ));
    CascadeMux I__11138 (
            .O(N__50148),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_267_cascade_ ));
    InMux I__11137 (
            .O(N__50145),
            .I(N__50142));
    LocalMux I__11136 (
            .O(N__50142),
            .I(N__50134));
    InMux I__11135 (
            .O(N__50141),
            .I(N__50131));
    InMux I__11134 (
            .O(N__50140),
            .I(N__50126));
    InMux I__11133 (
            .O(N__50139),
            .I(N__50126));
    InMux I__11132 (
            .O(N__50138),
            .I(N__50121));
    InMux I__11131 (
            .O(N__50137),
            .I(N__50121));
    Span4Mux_h I__11130 (
            .O(N__50134),
            .I(N__50114));
    LocalMux I__11129 (
            .O(N__50131),
            .I(N__50114));
    LocalMux I__11128 (
            .O(N__50126),
            .I(N__50114));
    LocalMux I__11127 (
            .O(N__50121),
            .I(N__50109));
    Span4Mux_v I__11126 (
            .O(N__50114),
            .I(N__50106));
    InMux I__11125 (
            .O(N__50113),
            .I(N__50103));
    InMux I__11124 (
            .O(N__50112),
            .I(N__50100));
    Odrv4 I__11123 (
            .O(N__50109),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0 ));
    Odrv4 I__11122 (
            .O(N__50106),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0 ));
    LocalMux I__11121 (
            .O(N__50103),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0 ));
    LocalMux I__11120 (
            .O(N__50100),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0 ));
    CEMux I__11119 (
            .O(N__50091),
            .I(N__50088));
    LocalMux I__11118 (
            .O(N__50088),
            .I(N__50084));
    CEMux I__11117 (
            .O(N__50087),
            .I(N__50081));
    Span4Mux_h I__11116 (
            .O(N__50084),
            .I(N__50077));
    LocalMux I__11115 (
            .O(N__50081),
            .I(N__50073));
    CEMux I__11114 (
            .O(N__50080),
            .I(N__50070));
    Span4Mux_v I__11113 (
            .O(N__50077),
            .I(N__50067));
    CEMux I__11112 (
            .O(N__50076),
            .I(N__50064));
    Span4Mux_h I__11111 (
            .O(N__50073),
            .I(N__50061));
    LocalMux I__11110 (
            .O(N__50070),
            .I(N__50058));
    Span4Mux_v I__11109 (
            .O(N__50067),
            .I(N__50053));
    LocalMux I__11108 (
            .O(N__50064),
            .I(N__50053));
    Span4Mux_h I__11107 (
            .O(N__50061),
            .I(N__50046));
    Span4Mux_h I__11106 (
            .O(N__50058),
            .I(N__50043));
    Span4Mux_h I__11105 (
            .O(N__50053),
            .I(N__50040));
    CEMux I__11104 (
            .O(N__50052),
            .I(N__50037));
    InMux I__11103 (
            .O(N__50051),
            .I(N__50030));
    InMux I__11102 (
            .O(N__50050),
            .I(N__50030));
    InMux I__11101 (
            .O(N__50049),
            .I(N__50030));
    Odrv4 I__11100 (
            .O(N__50046),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ));
    Odrv4 I__11099 (
            .O(N__50043),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ));
    Odrv4 I__11098 (
            .O(N__50040),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ));
    LocalMux I__11097 (
            .O(N__50037),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ));
    LocalMux I__11096 (
            .O(N__50030),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ));
    CascadeMux I__11095 (
            .O(N__50019),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_1_1_i_m2_1_9_cascade_ ));
    InMux I__11094 (
            .O(N__50016),
            .I(N__50012));
    InMux I__11093 (
            .O(N__50015),
            .I(N__50009));
    LocalMux I__11092 (
            .O(N__50012),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_101 ));
    LocalMux I__11091 (
            .O(N__50009),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_101 ));
    InMux I__11090 (
            .O(N__50004),
            .I(N__50001));
    LocalMux I__11089 (
            .O(N__50001),
            .I(N__49998));
    Span4Mux_v I__11088 (
            .O(N__49998),
            .I(N__49994));
    InMux I__11087 (
            .O(N__49997),
            .I(N__49991));
    Odrv4 I__11086 (
            .O(N__49994),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0 ));
    LocalMux I__11085 (
            .O(N__49991),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0 ));
    CascadeMux I__11084 (
            .O(N__49986),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3_cascade_ ));
    InMux I__11083 (
            .O(N__49983),
            .I(N__49980));
    LocalMux I__11082 (
            .O(N__49980),
            .I(N__49977));
    Span4Mux_v I__11081 (
            .O(N__49977),
            .I(N__49974));
    Span4Mux_h I__11080 (
            .O(N__49974),
            .I(N__49971));
    Span4Mux_h I__11079 (
            .O(N__49971),
            .I(N__49968));
    Odrv4 I__11078 (
            .O(N__49968),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_3 ));
    InMux I__11077 (
            .O(N__49965),
            .I(N__49962));
    LocalMux I__11076 (
            .O(N__49962),
            .I(N__49958));
    InMux I__11075 (
            .O(N__49961),
            .I(N__49955));
    Span4Mux_h I__11074 (
            .O(N__49958),
            .I(N__49952));
    LocalMux I__11073 (
            .O(N__49955),
            .I(N__49949));
    Span4Mux_v I__11072 (
            .O(N__49952),
            .I(N__49943));
    Span4Mux_h I__11071 (
            .O(N__49949),
            .I(N__49943));
    InMux I__11070 (
            .O(N__49948),
            .I(N__49940));
    Odrv4 I__11069 (
            .O(N__49943),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_2));
    LocalMux I__11068 (
            .O(N__49940),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_2));
    CascadeMux I__11067 (
            .O(N__49935),
            .I(N__49932));
    InMux I__11066 (
            .O(N__49932),
            .I(N__49929));
    LocalMux I__11065 (
            .O(N__49929),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_2 ));
    InMux I__11064 (
            .O(N__49926),
            .I(N__49923));
    LocalMux I__11063 (
            .O(N__49923),
            .I(N__49920));
    Odrv4 I__11062 (
            .O(N__49920),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_2 ));
    CascadeMux I__11061 (
            .O(N__49917),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2QZ0Z5_cascade_ ));
    InMux I__11060 (
            .O(N__49914),
            .I(N__49911));
    LocalMux I__11059 (
            .O(N__49911),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2 ));
    CascadeMux I__11058 (
            .O(N__49908),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2_cascade_ ));
    InMux I__11057 (
            .O(N__49905),
            .I(N__49902));
    LocalMux I__11056 (
            .O(N__49902),
            .I(N__49899));
    Sp12to4 I__11055 (
            .O(N__49899),
            .I(N__49896));
    Odrv12 I__11054 (
            .O(N__49896),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_2 ));
    CascadeMux I__11053 (
            .O(N__49893),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_6_0_0_cascade_ ));
    InMux I__11052 (
            .O(N__49890),
            .I(N__49887));
    LocalMux I__11051 (
            .O(N__49887),
            .I(N__49884));
    Span12Mux_v I__11050 (
            .O(N__49884),
            .I(N__49881));
    Odrv12 I__11049 (
            .O(N__49881),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_607 ));
    CascadeMux I__11048 (
            .O(N__49878),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_15_cascade_ ));
    InMux I__11047 (
            .O(N__49875),
            .I(N__49872));
    LocalMux I__11046 (
            .O(N__49872),
            .I(N__49869));
    Span4Mux_h I__11045 (
            .O(N__49869),
            .I(N__49866));
    Span4Mux_h I__11044 (
            .O(N__49866),
            .I(N__49863));
    Odrv4 I__11043 (
            .O(N__49863),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_1_15 ));
    CascadeMux I__11042 (
            .O(N__49860),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10_cascade_ ));
    InMux I__11041 (
            .O(N__49857),
            .I(N__49854));
    LocalMux I__11040 (
            .O(N__49854),
            .I(N__49851));
    Span4Mux_v I__11039 (
            .O(N__49851),
            .I(N__49848));
    Span4Mux_h I__11038 (
            .O(N__49848),
            .I(N__49845));
    Odrv4 I__11037 (
            .O(N__49845),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_10 ));
    InMux I__11036 (
            .O(N__49842),
            .I(N__49839));
    LocalMux I__11035 (
            .O(N__49839),
            .I(N__49836));
    Span4Mux_h I__11034 (
            .O(N__49836),
            .I(N__49833));
    Span4Mux_v I__11033 (
            .O(N__49833),
            .I(N__49829));
    InMux I__11032 (
            .O(N__49832),
            .I(N__49826));
    Sp12to4 I__11031 (
            .O(N__49829),
            .I(N__49823));
    LocalMux I__11030 (
            .O(N__49826),
            .I(N__49820));
    Span12Mux_h I__11029 (
            .O(N__49823),
            .I(N__49816));
    Span4Mux_v I__11028 (
            .O(N__49820),
            .I(N__49813));
    InMux I__11027 (
            .O(N__49819),
            .I(N__49810));
    Odrv12 I__11026 (
            .O(N__49816),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_9));
    Odrv4 I__11025 (
            .O(N__49813),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_9));
    LocalMux I__11024 (
            .O(N__49810),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_9));
    CascadeMux I__11023 (
            .O(N__49803),
            .I(N__49800));
    InMux I__11022 (
            .O(N__49800),
            .I(N__49797));
    LocalMux I__11021 (
            .O(N__49797),
            .I(N__49794));
    Odrv4 I__11020 (
            .O(N__49794),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_9 ));
    InMux I__11019 (
            .O(N__49791),
            .I(N__49788));
    LocalMux I__11018 (
            .O(N__49788),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_9 ));
    CascadeMux I__11017 (
            .O(N__49785),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044QZ0Z5_cascade_ ));
    InMux I__11016 (
            .O(N__49782),
            .I(N__49779));
    LocalMux I__11015 (
            .O(N__49779),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9 ));
    InMux I__11014 (
            .O(N__49776),
            .I(N__49773));
    LocalMux I__11013 (
            .O(N__49773),
            .I(N__49770));
    Span4Mux_v I__11012 (
            .O(N__49770),
            .I(N__49767));
    Span4Mux_v I__11011 (
            .O(N__49767),
            .I(N__49764));
    Odrv4 I__11010 (
            .O(N__49764),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_8 ));
    CascadeMux I__11009 (
            .O(N__49761),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9_cascade_ ));
    InMux I__11008 (
            .O(N__49758),
            .I(N__49755));
    LocalMux I__11007 (
            .O(N__49755),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_9 ));
    InMux I__11006 (
            .O(N__49752),
            .I(N__49748));
    InMux I__11005 (
            .O(N__49751),
            .I(N__49744));
    LocalMux I__11004 (
            .O(N__49748),
            .I(N__49741));
    CascadeMux I__11003 (
            .O(N__49747),
            .I(N__49738));
    LocalMux I__11002 (
            .O(N__49744),
            .I(N__49735));
    Span12Mux_v I__11001 (
            .O(N__49741),
            .I(N__49732));
    InMux I__11000 (
            .O(N__49738),
            .I(N__49729));
    Span4Mux_v I__10999 (
            .O(N__49735),
            .I(N__49726));
    Odrv12 I__10998 (
            .O(N__49732),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_2));
    LocalMux I__10997 (
            .O(N__49729),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_2));
    Odrv4 I__10996 (
            .O(N__49726),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_2));
    InMux I__10995 (
            .O(N__49719),
            .I(N__49715));
    CascadeMux I__10994 (
            .O(N__49718),
            .I(N__49712));
    LocalMux I__10993 (
            .O(N__49715),
            .I(N__49709));
    InMux I__10992 (
            .O(N__49712),
            .I(N__49706));
    Span4Mux_v I__10991 (
            .O(N__49709),
            .I(N__49703));
    LocalMux I__10990 (
            .O(N__49706),
            .I(N__49700));
    Sp12to4 I__10989 (
            .O(N__49703),
            .I(N__49697));
    Span4Mux_h I__10988 (
            .O(N__49700),
            .I(N__49694));
    Span12Mux_h I__10987 (
            .O(N__49697),
            .I(N__49690));
    Span4Mux_v I__10986 (
            .O(N__49694),
            .I(N__49687));
    InMux I__10985 (
            .O(N__49693),
            .I(N__49684));
    Odrv12 I__10984 (
            .O(N__49690),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_3));
    Odrv4 I__10983 (
            .O(N__49687),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_3));
    LocalMux I__10982 (
            .O(N__49684),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_3));
    InMux I__10981 (
            .O(N__49677),
            .I(N__49673));
    InMux I__10980 (
            .O(N__49676),
            .I(N__49670));
    LocalMux I__10979 (
            .O(N__49673),
            .I(N__49666));
    LocalMux I__10978 (
            .O(N__49670),
            .I(N__49663));
    InMux I__10977 (
            .O(N__49669),
            .I(N__49660));
    Span4Mux_v I__10976 (
            .O(N__49666),
            .I(N__49657));
    Span4Mux_v I__10975 (
            .O(N__49663),
            .I(N__49654));
    LocalMux I__10974 (
            .O(N__49660),
            .I(N__49651));
    Span4Mux_h I__10973 (
            .O(N__49657),
            .I(N__49648));
    Odrv4 I__10972 (
            .O(N__49654),
            .I(cemf_module_64ch_ctrl_inst1_data_config_3));
    Odrv4 I__10971 (
            .O(N__49651),
            .I(cemf_module_64ch_ctrl_inst1_data_config_3));
    Odrv4 I__10970 (
            .O(N__49648),
            .I(cemf_module_64ch_ctrl_inst1_data_config_3));
    InMux I__10969 (
            .O(N__49641),
            .I(N__49638));
    LocalMux I__10968 (
            .O(N__49638),
            .I(N__49633));
    InMux I__10967 (
            .O(N__49637),
            .I(N__49630));
    CascadeMux I__10966 (
            .O(N__49636),
            .I(N__49627));
    Span4Mux_v I__10965 (
            .O(N__49633),
            .I(N__49624));
    LocalMux I__10964 (
            .O(N__49630),
            .I(N__49621));
    InMux I__10963 (
            .O(N__49627),
            .I(N__49618));
    Span4Mux_h I__10962 (
            .O(N__49624),
            .I(N__49615));
    Span4Mux_v I__10961 (
            .O(N__49621),
            .I(N__49612));
    LocalMux I__10960 (
            .O(N__49618),
            .I(N__49609));
    Span4Mux_h I__10959 (
            .O(N__49615),
            .I(N__49602));
    Span4Mux_v I__10958 (
            .O(N__49612),
            .I(N__49602));
    Span4Mux_v I__10957 (
            .O(N__49609),
            .I(N__49602));
    Odrv4 I__10956 (
            .O(N__49602),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_3));
    CascadeMux I__10955 (
            .O(N__49599),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_3_cascade_ ));
    InMux I__10954 (
            .O(N__49596),
            .I(N__49593));
    LocalMux I__10953 (
            .O(N__49593),
            .I(N__49590));
    Span4Mux_h I__10952 (
            .O(N__49590),
            .I(N__49587));
    Span4Mux_h I__10951 (
            .O(N__49587),
            .I(N__49584));
    Odrv4 I__10950 (
            .O(N__49584),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_3 ));
    CascadeMux I__10949 (
            .O(N__49581),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253QZ0Z5_cascade_ ));
    InMux I__10948 (
            .O(N__49578),
            .I(N__49575));
    LocalMux I__10947 (
            .O(N__49575),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3 ));
    CascadeMux I__10946 (
            .O(N__49572),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLHZ0Z5_cascade_ ));
    InMux I__10945 (
            .O(N__49569),
            .I(N__49566));
    LocalMux I__10944 (
            .O(N__49566),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23 ));
    CascadeMux I__10943 (
            .O(N__49563),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23_cascade_ ));
    InMux I__10942 (
            .O(N__49560),
            .I(N__49557));
    LocalMux I__10941 (
            .O(N__49557),
            .I(N__49554));
    Span4Mux_v I__10940 (
            .O(N__49554),
            .I(N__49551));
    Span4Mux_v I__10939 (
            .O(N__49551),
            .I(N__49548));
    Sp12to4 I__10938 (
            .O(N__49548),
            .I(N__49545));
    Span12Mux_h I__10937 (
            .O(N__49545),
            .I(N__49542));
    Odrv12 I__10936 (
            .O(N__49542),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.dout_conf ));
    CascadeMux I__10935 (
            .O(N__49539),
            .I(N__49536));
    InMux I__10934 (
            .O(N__49536),
            .I(N__49533));
    LocalMux I__10933 (
            .O(N__49533),
            .I(N__49530));
    Odrv12 I__10932 (
            .O(N__49530),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALHZ0Z5 ));
    InMux I__10931 (
            .O(N__49527),
            .I(N__49524));
    LocalMux I__10930 (
            .O(N__49524),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22 ));
    InMux I__10929 (
            .O(N__49521),
            .I(N__49518));
    LocalMux I__10928 (
            .O(N__49518),
            .I(N__49515));
    Span4Mux_v I__10927 (
            .O(N__49515),
            .I(N__49512));
    Sp12to4 I__10926 (
            .O(N__49512),
            .I(N__49509));
    Odrv12 I__10925 (
            .O(N__49509),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_21 ));
    CascadeMux I__10924 (
            .O(N__49506),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22_cascade_ ));
    InMux I__10923 (
            .O(N__49503),
            .I(N__49500));
    LocalMux I__10922 (
            .O(N__49500),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_22 ));
    InMux I__10921 (
            .O(N__49497),
            .I(N__49494));
    LocalMux I__10920 (
            .O(N__49494),
            .I(N__49490));
    CascadeMux I__10919 (
            .O(N__49493),
            .I(N__49487));
    Span4Mux_h I__10918 (
            .O(N__49490),
            .I(N__49484));
    InMux I__10917 (
            .O(N__49487),
            .I(N__49481));
    Span4Mux_v I__10916 (
            .O(N__49484),
            .I(N__49477));
    LocalMux I__10915 (
            .O(N__49481),
            .I(N__49474));
    InMux I__10914 (
            .O(N__49480),
            .I(N__49471));
    Odrv4 I__10913 (
            .O(N__49477),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_23));
    Odrv12 I__10912 (
            .O(N__49474),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_23));
    LocalMux I__10911 (
            .O(N__49471),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_23));
    InMux I__10910 (
            .O(N__49464),
            .I(N__49461));
    LocalMux I__10909 (
            .O(N__49461),
            .I(N__49458));
    Span4Mux_h I__10908 (
            .O(N__49458),
            .I(N__49455));
    Span4Mux_v I__10907 (
            .O(N__49455),
            .I(N__49450));
    InMux I__10906 (
            .O(N__49454),
            .I(N__49447));
    InMux I__10905 (
            .O(N__49453),
            .I(N__49444));
    Odrv4 I__10904 (
            .O(N__49450),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_23));
    LocalMux I__10903 (
            .O(N__49447),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_23));
    LocalMux I__10902 (
            .O(N__49444),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_23));
    InMux I__10901 (
            .O(N__49437),
            .I(N__49434));
    LocalMux I__10900 (
            .O(N__49434),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_23 ));
    CascadeMux I__10899 (
            .O(N__49431),
            .I(N__49428));
    InMux I__10898 (
            .O(N__49428),
            .I(N__49424));
    InMux I__10897 (
            .O(N__49427),
            .I(N__49420));
    LocalMux I__10896 (
            .O(N__49424),
            .I(N__49417));
    InMux I__10895 (
            .O(N__49423),
            .I(N__49414));
    LocalMux I__10894 (
            .O(N__49420),
            .I(N__49411));
    Span4Mux_h I__10893 (
            .O(N__49417),
            .I(N__49408));
    LocalMux I__10892 (
            .O(N__49414),
            .I(N__49405));
    Span4Mux_v I__10891 (
            .O(N__49411),
            .I(N__49402));
    Span4Mux_v I__10890 (
            .O(N__49408),
            .I(N__49399));
    Span4Mux_v I__10889 (
            .O(N__49405),
            .I(N__49394));
    Span4Mux_h I__10888 (
            .O(N__49402),
            .I(N__49394));
    Span4Mux_h I__10887 (
            .O(N__49399),
            .I(N__49391));
    Odrv4 I__10886 (
            .O(N__49394),
            .I(cemf_module_64ch_ctrl_inst1_data_config_9));
    Odrv4 I__10885 (
            .O(N__49391),
            .I(cemf_module_64ch_ctrl_inst1_data_config_9));
    InMux I__10884 (
            .O(N__49386),
            .I(N__49383));
    LocalMux I__10883 (
            .O(N__49383),
            .I(N__49379));
    CascadeMux I__10882 (
            .O(N__49382),
            .I(N__49375));
    Span4Mux_v I__10881 (
            .O(N__49379),
            .I(N__49372));
    InMux I__10880 (
            .O(N__49378),
            .I(N__49369));
    InMux I__10879 (
            .O(N__49375),
            .I(N__49366));
    Span4Mux_h I__10878 (
            .O(N__49372),
            .I(N__49363));
    LocalMux I__10877 (
            .O(N__49369),
            .I(N__49360));
    LocalMux I__10876 (
            .O(N__49366),
            .I(N__49357));
    Span4Mux_v I__10875 (
            .O(N__49363),
            .I(N__49354));
    Span4Mux_h I__10874 (
            .O(N__49360),
            .I(N__49349));
    Span4Mux_h I__10873 (
            .O(N__49357),
            .I(N__49349));
    Odrv4 I__10872 (
            .O(N__49354),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_9));
    Odrv4 I__10871 (
            .O(N__49349),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_9));
    CascadeMux I__10870 (
            .O(N__49344),
            .I(N__49341));
    InMux I__10869 (
            .O(N__49341),
            .I(N__49336));
    InMux I__10868 (
            .O(N__49340),
            .I(N__49333));
    CascadeMux I__10867 (
            .O(N__49339),
            .I(N__49330));
    LocalMux I__10866 (
            .O(N__49336),
            .I(N__49327));
    LocalMux I__10865 (
            .O(N__49333),
            .I(N__49324));
    InMux I__10864 (
            .O(N__49330),
            .I(N__49321));
    Span4Mux_h I__10863 (
            .O(N__49327),
            .I(N__49318));
    Span12Mux_v I__10862 (
            .O(N__49324),
            .I(N__49313));
    LocalMux I__10861 (
            .O(N__49321),
            .I(N__49313));
    Odrv4 I__10860 (
            .O(N__49318),
            .I(cemf_module_64ch_ctrl_inst1_data_config_10));
    Odrv12 I__10859 (
            .O(N__49313),
            .I(cemf_module_64ch_ctrl_inst1_data_config_10));
    InMux I__10858 (
            .O(N__49308),
            .I(N__49304));
    InMux I__10857 (
            .O(N__49307),
            .I(N__49301));
    LocalMux I__10856 (
            .O(N__49304),
            .I(N__49298));
    LocalMux I__10855 (
            .O(N__49301),
            .I(N__49295));
    Span4Mux_v I__10854 (
            .O(N__49298),
            .I(N__49292));
    Span4Mux_h I__10853 (
            .O(N__49295),
            .I(N__49289));
    Span4Mux_h I__10852 (
            .O(N__49292),
            .I(N__49286));
    Span4Mux_h I__10851 (
            .O(N__49289),
            .I(N__49282));
    Sp12to4 I__10850 (
            .O(N__49286),
            .I(N__49279));
    InMux I__10849 (
            .O(N__49285),
            .I(N__49276));
    Odrv4 I__10848 (
            .O(N__49282),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_10));
    Odrv12 I__10847 (
            .O(N__49279),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_10));
    LocalMux I__10846 (
            .O(N__49276),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_10));
    InMux I__10845 (
            .O(N__49269),
            .I(N__49265));
    InMux I__10844 (
            .O(N__49268),
            .I(N__49262));
    LocalMux I__10843 (
            .O(N__49265),
            .I(N__49259));
    LocalMux I__10842 (
            .O(N__49262),
            .I(N__49256));
    Span4Mux_v I__10841 (
            .O(N__49259),
            .I(N__49252));
    Span4Mux_v I__10840 (
            .O(N__49256),
            .I(N__49249));
    CascadeMux I__10839 (
            .O(N__49255),
            .I(N__49246));
    Span4Mux_h I__10838 (
            .O(N__49252),
            .I(N__49241));
    Span4Mux_h I__10837 (
            .O(N__49249),
            .I(N__49241));
    InMux I__10836 (
            .O(N__49246),
            .I(N__49238));
    Odrv4 I__10835 (
            .O(N__49241),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_10));
    LocalMux I__10834 (
            .O(N__49238),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_10));
    CascadeMux I__10833 (
            .O(N__49233),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_10_cascade_ ));
    InMux I__10832 (
            .O(N__49230),
            .I(N__49227));
    LocalMux I__10831 (
            .O(N__49227),
            .I(N__49224));
    Span4Mux_v I__10830 (
            .O(N__49224),
            .I(N__49221));
    Odrv4 I__10829 (
            .O(N__49221),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_10 ));
    CascadeMux I__10828 (
            .O(N__49218),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFHZ0Z5_cascade_ ));
    InMux I__10827 (
            .O(N__49215),
            .I(N__49212));
    LocalMux I__10826 (
            .O(N__49212),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10 ));
    CascadeMux I__10825 (
            .O(N__49209),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9DZ0Z7_cascade_ ));
    InMux I__10824 (
            .O(N__49206),
            .I(N__49203));
    LocalMux I__10823 (
            .O(N__49203),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19 ));
    CascadeMux I__10822 (
            .O(N__49200),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19_cascade_ ));
    InMux I__10821 (
            .O(N__49197),
            .I(N__49194));
    LocalMux I__10820 (
            .O(N__49194),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_18 ));
    InMux I__10819 (
            .O(N__49191),
            .I(N__49188));
    LocalMux I__10818 (
            .O(N__49188),
            .I(N__49185));
    Span4Mux_h I__10817 (
            .O(N__49185),
            .I(N__49182));
    Span4Mux_h I__10816 (
            .O(N__49182),
            .I(N__49179));
    Span4Mux_v I__10815 (
            .O(N__49179),
            .I(N__49176));
    Odrv4 I__10814 (
            .O(N__49176),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_19 ));
    InMux I__10813 (
            .O(N__49173),
            .I(N__49170));
    LocalMux I__10812 (
            .O(N__49170),
            .I(N__49167));
    Span4Mux_h I__10811 (
            .O(N__49167),
            .I(N__49164));
    Span4Mux_h I__10810 (
            .O(N__49164),
            .I(N__49160));
    CascadeMux I__10809 (
            .O(N__49163),
            .I(N__49157));
    Span4Mux_h I__10808 (
            .O(N__49160),
            .I(N__49153));
    InMux I__10807 (
            .O(N__49157),
            .I(N__49148));
    InMux I__10806 (
            .O(N__49156),
            .I(N__49148));
    Odrv4 I__10805 (
            .O(N__49153),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_18));
    LocalMux I__10804 (
            .O(N__49148),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_18));
    InMux I__10803 (
            .O(N__49143),
            .I(N__49140));
    LocalMux I__10802 (
            .O(N__49140),
            .I(N__49137));
    Span4Mux_v I__10801 (
            .O(N__49137),
            .I(N__49134));
    Span4Mux_v I__10800 (
            .O(N__49134),
            .I(N__49131));
    Odrv4 I__10799 (
            .O(N__49131),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_27));
    InMux I__10798 (
            .O(N__49128),
            .I(N__49125));
    LocalMux I__10797 (
            .O(N__49125),
            .I(N__49122));
    Span4Mux_h I__10796 (
            .O(N__49122),
            .I(N__49119));
    Span4Mux_h I__10795 (
            .O(N__49119),
            .I(N__49116));
    Span4Mux_h I__10794 (
            .O(N__49116),
            .I(N__49113));
    Odrv4 I__10793 (
            .O(N__49113),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_28));
    InMux I__10792 (
            .O(N__49110),
            .I(N__49107));
    LocalMux I__10791 (
            .O(N__49107),
            .I(N__49104));
    Span4Mux_h I__10790 (
            .O(N__49104),
            .I(N__49101));
    Span4Mux_v I__10789 (
            .O(N__49101),
            .I(N__49098));
    Odrv4 I__10788 (
            .O(N__49098),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_29));
    CEMux I__10787 (
            .O(N__49095),
            .I(N__49090));
    CEMux I__10786 (
            .O(N__49094),
            .I(N__49087));
    CEMux I__10785 (
            .O(N__49093),
            .I(N__49084));
    LocalMux I__10784 (
            .O(N__49090),
            .I(N__49080));
    LocalMux I__10783 (
            .O(N__49087),
            .I(N__49075));
    LocalMux I__10782 (
            .O(N__49084),
            .I(N__49075));
    CEMux I__10781 (
            .O(N__49083),
            .I(N__49072));
    Span4Mux_v I__10780 (
            .O(N__49080),
            .I(N__49064));
    Span4Mux_v I__10779 (
            .O(N__49075),
            .I(N__49064));
    LocalMux I__10778 (
            .O(N__49072),
            .I(N__49064));
    CEMux I__10777 (
            .O(N__49071),
            .I(N__49060));
    Span4Mux_h I__10776 (
            .O(N__49064),
            .I(N__49056));
    CEMux I__10775 (
            .O(N__49063),
            .I(N__49053));
    LocalMux I__10774 (
            .O(N__49060),
            .I(N__49050));
    CEMux I__10773 (
            .O(N__49059),
            .I(N__49047));
    Span4Mux_v I__10772 (
            .O(N__49056),
            .I(N__49044));
    LocalMux I__10771 (
            .O(N__49053),
            .I(N__49041));
    Span4Mux_v I__10770 (
            .O(N__49050),
            .I(N__49038));
    LocalMux I__10769 (
            .O(N__49047),
            .I(N__49035));
    Span4Mux_h I__10768 (
            .O(N__49044),
            .I(N__49028));
    Span4Mux_h I__10767 (
            .O(N__49041),
            .I(N__49028));
    Span4Mux_h I__10766 (
            .O(N__49038),
            .I(N__49023));
    Span4Mux_h I__10765 (
            .O(N__49035),
            .I(N__49023));
    CEMux I__10764 (
            .O(N__49034),
            .I(N__49020));
    CEMux I__10763 (
            .O(N__49033),
            .I(N__49017));
    Odrv4 I__10762 (
            .O(N__49028),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0 ));
    Odrv4 I__10761 (
            .O(N__49023),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0 ));
    LocalMux I__10760 (
            .O(N__49020),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0 ));
    LocalMux I__10759 (
            .O(N__49017),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0 ));
    CascadeMux I__10758 (
            .O(N__49008),
            .I(N__49005));
    InMux I__10757 (
            .O(N__49005),
            .I(N__49000));
    InMux I__10756 (
            .O(N__49004),
            .I(N__48997));
    InMux I__10755 (
            .O(N__49003),
            .I(N__48994));
    LocalMux I__10754 (
            .O(N__49000),
            .I(N__48991));
    LocalMux I__10753 (
            .O(N__48997),
            .I(N__48988));
    LocalMux I__10752 (
            .O(N__48994),
            .I(N__48985));
    Span4Mux_h I__10751 (
            .O(N__48991),
            .I(N__48982));
    Odrv12 I__10750 (
            .O(N__48988),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_23));
    Odrv4 I__10749 (
            .O(N__48985),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_23));
    Odrv4 I__10748 (
            .O(N__48982),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_23));
    InMux I__10747 (
            .O(N__48975),
            .I(N__48971));
    InMux I__10746 (
            .O(N__48974),
            .I(N__48968));
    LocalMux I__10745 (
            .O(N__48971),
            .I(N__48965));
    LocalMux I__10744 (
            .O(N__48968),
            .I(N__48961));
    Span4Mux_h I__10743 (
            .O(N__48965),
            .I(N__48958));
    InMux I__10742 (
            .O(N__48964),
            .I(N__48955));
    Span4Mux_h I__10741 (
            .O(N__48961),
            .I(N__48950));
    Span4Mux_h I__10740 (
            .O(N__48958),
            .I(N__48950));
    LocalMux I__10739 (
            .O(N__48955),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_23));
    Odrv4 I__10738 (
            .O(N__48950),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_23));
    CascadeMux I__10737 (
            .O(N__48945),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_23_cascade_ ));
    InMux I__10736 (
            .O(N__48942),
            .I(N__48939));
    LocalMux I__10735 (
            .O(N__48939),
            .I(N__48936));
    Span4Mux_h I__10734 (
            .O(N__48936),
            .I(N__48931));
    InMux I__10733 (
            .O(N__48935),
            .I(N__48926));
    InMux I__10732 (
            .O(N__48934),
            .I(N__48926));
    Odrv4 I__10731 (
            .O(N__48931),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_0));
    LocalMux I__10730 (
            .O(N__48926),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_0));
    InMux I__10729 (
            .O(N__48921),
            .I(N__48918));
    LocalMux I__10728 (
            .O(N__48918),
            .I(N__48915));
    Span4Mux_h I__10727 (
            .O(N__48915),
            .I(N__48911));
    CascadeMux I__10726 (
            .O(N__48914),
            .I(N__48907));
    Span4Mux_h I__10725 (
            .O(N__48911),
            .I(N__48904));
    InMux I__10724 (
            .O(N__48910),
            .I(N__48901));
    InMux I__10723 (
            .O(N__48907),
            .I(N__48898));
    Odrv4 I__10722 (
            .O(N__48904),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_0));
    LocalMux I__10721 (
            .O(N__48901),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_0));
    LocalMux I__10720 (
            .O(N__48898),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_0));
    InMux I__10719 (
            .O(N__48891),
            .I(N__48888));
    LocalMux I__10718 (
            .O(N__48888),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_0 ));
    CascadeMux I__10717 (
            .O(N__48885),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_0_cascade_ ));
    CascadeMux I__10716 (
            .O(N__48882),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQLZ0Z7_cascade_ ));
    InMux I__10715 (
            .O(N__48879),
            .I(N__48875));
    InMux I__10714 (
            .O(N__48878),
            .I(N__48872));
    LocalMux I__10713 (
            .O(N__48875),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0 ));
    LocalMux I__10712 (
            .O(N__48872),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0 ));
    CascadeMux I__10711 (
            .O(N__48867),
            .I(N__48863));
    InMux I__10710 (
            .O(N__48866),
            .I(N__48859));
    InMux I__10709 (
            .O(N__48863),
            .I(N__48856));
    InMux I__10708 (
            .O(N__48862),
            .I(N__48853));
    LocalMux I__10707 (
            .O(N__48859),
            .I(N__48848));
    LocalMux I__10706 (
            .O(N__48856),
            .I(N__48848));
    LocalMux I__10705 (
            .O(N__48853),
            .I(N__48845));
    Span4Mux_v I__10704 (
            .O(N__48848),
            .I(N__48842));
    Odrv12 I__10703 (
            .O(N__48845),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_18));
    Odrv4 I__10702 (
            .O(N__48842),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_18));
    CascadeMux I__10701 (
            .O(N__48837),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_18_cascade_ ));
    InMux I__10700 (
            .O(N__48834),
            .I(N__48831));
    LocalMux I__10699 (
            .O(N__48831),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_18 ));
    CascadeMux I__10698 (
            .O(N__48828),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579DZ0Z7_cascade_ ));
    InMux I__10697 (
            .O(N__48825),
            .I(N__48822));
    LocalMux I__10696 (
            .O(N__48822),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18 ));
    InMux I__10695 (
            .O(N__48819),
            .I(N__48816));
    LocalMux I__10694 (
            .O(N__48816),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_17 ));
    CascadeMux I__10693 (
            .O(N__48813),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18_cascade_ ));
    CascadeMux I__10692 (
            .O(N__48810),
            .I(N__48807));
    InMux I__10691 (
            .O(N__48807),
            .I(N__48804));
    LocalMux I__10690 (
            .O(N__48804),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_19 ));
    InMux I__10689 (
            .O(N__48801),
            .I(N__48798));
    LocalMux I__10688 (
            .O(N__48798),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_19 ));
    CascadeMux I__10687 (
            .O(N__48795),
            .I(N__48792));
    InMux I__10686 (
            .O(N__48792),
            .I(N__48789));
    LocalMux I__10685 (
            .O(N__48789),
            .I(N__48786));
    Span4Mux_v I__10684 (
            .O(N__48786),
            .I(N__48783));
    Span4Mux_h I__10683 (
            .O(N__48783),
            .I(N__48780));
    Span4Mux_h I__10682 (
            .O(N__48780),
            .I(N__48777));
    Odrv4 I__10681 (
            .O(N__48777),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_28));
    CascadeMux I__10680 (
            .O(N__48774),
            .I(N__48771));
    InMux I__10679 (
            .O(N__48771),
            .I(N__48768));
    LocalMux I__10678 (
            .O(N__48768),
            .I(N__48765));
    Span4Mux_h I__10677 (
            .O(N__48765),
            .I(N__48762));
    Odrv4 I__10676 (
            .O(N__48762),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_29));
    InMux I__10675 (
            .O(N__48759),
            .I(N__48756));
    LocalMux I__10674 (
            .O(N__48756),
            .I(N__48753));
    Span4Mux_v I__10673 (
            .O(N__48753),
            .I(N__48750));
    Sp12to4 I__10672 (
            .O(N__48750),
            .I(N__48746));
    InMux I__10671 (
            .O(N__48749),
            .I(N__48742));
    Span12Mux_h I__10670 (
            .O(N__48746),
            .I(N__48739));
    InMux I__10669 (
            .O(N__48745),
            .I(N__48736));
    LocalMux I__10668 (
            .O(N__48742),
            .I(N__48733));
    Odrv12 I__10667 (
            .O(N__48739),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_7));
    LocalMux I__10666 (
            .O(N__48736),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_7));
    Odrv4 I__10665 (
            .O(N__48733),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_7));
    CEMux I__10664 (
            .O(N__48726),
            .I(N__48711));
    CEMux I__10663 (
            .O(N__48725),
            .I(N__48711));
    CEMux I__10662 (
            .O(N__48724),
            .I(N__48711));
    CEMux I__10661 (
            .O(N__48723),
            .I(N__48711));
    CEMux I__10660 (
            .O(N__48722),
            .I(N__48711));
    GlobalMux I__10659 (
            .O(N__48711),
            .I(N__48708));
    gio2CtrlBuf I__10658 (
            .O(N__48708),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g ));
    InMux I__10657 (
            .O(N__48705),
            .I(N__48702));
    LocalMux I__10656 (
            .O(N__48702),
            .I(N__48698));
    CascadeMux I__10655 (
            .O(N__48701),
            .I(N__48695));
    Span4Mux_v I__10654 (
            .O(N__48698),
            .I(N__48691));
    InMux I__10653 (
            .O(N__48695),
            .I(N__48686));
    InMux I__10652 (
            .O(N__48694),
            .I(N__48686));
    Odrv4 I__10651 (
            .O(N__48691),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_19));
    LocalMux I__10650 (
            .O(N__48686),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_19));
    InMux I__10649 (
            .O(N__48681),
            .I(N__48678));
    LocalMux I__10648 (
            .O(N__48678),
            .I(N__48674));
    CascadeMux I__10647 (
            .O(N__48677),
            .I(N__48671));
    Span12Mux_s10_v I__10646 (
            .O(N__48674),
            .I(N__48667));
    InMux I__10645 (
            .O(N__48671),
            .I(N__48664));
    InMux I__10644 (
            .O(N__48670),
            .I(N__48661));
    Odrv12 I__10643 (
            .O(N__48667),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_19));
    LocalMux I__10642 (
            .O(N__48664),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_19));
    LocalMux I__10641 (
            .O(N__48661),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_19));
    InMux I__10640 (
            .O(N__48654),
            .I(N__48642));
    InMux I__10639 (
            .O(N__48653),
            .I(N__48642));
    InMux I__10638 (
            .O(N__48652),
            .I(N__48642));
    InMux I__10637 (
            .O(N__48651),
            .I(N__48642));
    LocalMux I__10636 (
            .O(N__48642),
            .I(N__48635));
    InMux I__10635 (
            .O(N__48641),
            .I(N__48626));
    InMux I__10634 (
            .O(N__48640),
            .I(N__48626));
    InMux I__10633 (
            .O(N__48639),
            .I(N__48626));
    InMux I__10632 (
            .O(N__48638),
            .I(N__48626));
    Odrv4 I__10631 (
            .O(N__48635),
            .I(\serializer_mod_inst.next_state32_i ));
    LocalMux I__10630 (
            .O(N__48626),
            .I(\serializer_mod_inst.next_state32_i ));
    InMux I__10629 (
            .O(N__48621),
            .I(\serializer_mod_inst.counter_sr_cry_6 ));
    InMux I__10628 (
            .O(N__48618),
            .I(N__48613));
    InMux I__10627 (
            .O(N__48617),
            .I(N__48610));
    InMux I__10626 (
            .O(N__48616),
            .I(N__48607));
    LocalMux I__10625 (
            .O(N__48613),
            .I(\serializer_mod_inst.counter_srZ0Z_7 ));
    LocalMux I__10624 (
            .O(N__48610),
            .I(\serializer_mod_inst.counter_srZ0Z_7 ));
    LocalMux I__10623 (
            .O(N__48607),
            .I(\serializer_mod_inst.counter_srZ0Z_7 ));
    CEMux I__10622 (
            .O(N__48600),
            .I(N__48597));
    LocalMux I__10621 (
            .O(N__48597),
            .I(N__48594));
    Span4Mux_v I__10620 (
            .O(N__48594),
            .I(N__48591));
    Span4Mux_h I__10619 (
            .O(N__48591),
            .I(N__48588));
    Odrv4 I__10618 (
            .O(N__48588),
            .I(\serializer_mod_inst.counter_sre_0_i ));
    CascadeMux I__10617 (
            .O(N__48585),
            .I(N__48582));
    InMux I__10616 (
            .O(N__48582),
            .I(N__48578));
    InMux I__10615 (
            .O(N__48581),
            .I(N__48575));
    LocalMux I__10614 (
            .O(N__48578),
            .I(N__48572));
    LocalMux I__10613 (
            .O(N__48575),
            .I(N__48569));
    Span4Mux_v I__10612 (
            .O(N__48572),
            .I(N__48566));
    Span4Mux_v I__10611 (
            .O(N__48569),
            .I(N__48562));
    Span4Mux_v I__10610 (
            .O(N__48566),
            .I(N__48559));
    CascadeMux I__10609 (
            .O(N__48565),
            .I(N__48556));
    Span4Mux_h I__10608 (
            .O(N__48562),
            .I(N__48551));
    Span4Mux_h I__10607 (
            .O(N__48559),
            .I(N__48551));
    InMux I__10606 (
            .O(N__48556),
            .I(N__48548));
    Span4Mux_h I__10605 (
            .O(N__48551),
            .I(N__48545));
    LocalMux I__10604 (
            .O(N__48548),
            .I(N__48542));
    Odrv4 I__10603 (
            .O(N__48545),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_15));
    Odrv4 I__10602 (
            .O(N__48542),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_15));
    CascadeMux I__10601 (
            .O(N__48537),
            .I(N__48534));
    InMux I__10600 (
            .O(N__48534),
            .I(N__48531));
    LocalMux I__10599 (
            .O(N__48531),
            .I(N__48528));
    Span4Mux_v I__10598 (
            .O(N__48528),
            .I(N__48525));
    Span4Mux_h I__10597 (
            .O(N__48525),
            .I(N__48522));
    Odrv4 I__10596 (
            .O(N__48522),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_24));
    InMux I__10595 (
            .O(N__48519),
            .I(N__48516));
    LocalMux I__10594 (
            .O(N__48516),
            .I(N__48513));
    Span4Mux_v I__10593 (
            .O(N__48513),
            .I(N__48510));
    Span4Mux_h I__10592 (
            .O(N__48510),
            .I(N__48507));
    Odrv4 I__10591 (
            .O(N__48507),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_2Z0Z_26 ));
    CascadeMux I__10590 (
            .O(N__48504),
            .I(N__48501));
    InMux I__10589 (
            .O(N__48501),
            .I(N__48498));
    LocalMux I__10588 (
            .O(N__48498),
            .I(N__48495));
    Span4Mux_h I__10587 (
            .O(N__48495),
            .I(N__48492));
    Odrv4 I__10586 (
            .O(N__48492),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_27));
    InMux I__10585 (
            .O(N__48489),
            .I(N__48486));
    LocalMux I__10584 (
            .O(N__48486),
            .I(\serializer_mod_inst.un22_next_state_5 ));
    InMux I__10583 (
            .O(N__48483),
            .I(N__48479));
    InMux I__10582 (
            .O(N__48482),
            .I(N__48475));
    LocalMux I__10581 (
            .O(N__48479),
            .I(N__48472));
    InMux I__10580 (
            .O(N__48478),
            .I(N__48469));
    LocalMux I__10579 (
            .O(N__48475),
            .I(\serializer_mod_inst.counter_srZ0Z_0 ));
    Odrv4 I__10578 (
            .O(N__48472),
            .I(\serializer_mod_inst.counter_srZ0Z_0 ));
    LocalMux I__10577 (
            .O(N__48469),
            .I(\serializer_mod_inst.counter_srZ0Z_0 ));
    InMux I__10576 (
            .O(N__48462),
            .I(bfn_21_27_0_));
    CascadeMux I__10575 (
            .O(N__48459),
            .I(N__48454));
    InMux I__10574 (
            .O(N__48458),
            .I(N__48451));
    InMux I__10573 (
            .O(N__48457),
            .I(N__48448));
    InMux I__10572 (
            .O(N__48454),
            .I(N__48445));
    LocalMux I__10571 (
            .O(N__48451),
            .I(\serializer_mod_inst.counter_srZ0Z_1 ));
    LocalMux I__10570 (
            .O(N__48448),
            .I(\serializer_mod_inst.counter_srZ0Z_1 ));
    LocalMux I__10569 (
            .O(N__48445),
            .I(\serializer_mod_inst.counter_srZ0Z_1 ));
    InMux I__10568 (
            .O(N__48438),
            .I(\serializer_mod_inst.counter_sr_cry_0 ));
    InMux I__10567 (
            .O(N__48435),
            .I(N__48431));
    InMux I__10566 (
            .O(N__48434),
            .I(N__48427));
    LocalMux I__10565 (
            .O(N__48431),
            .I(N__48424));
    InMux I__10564 (
            .O(N__48430),
            .I(N__48421));
    LocalMux I__10563 (
            .O(N__48427),
            .I(\serializer_mod_inst.counter_srZ0Z_2 ));
    Odrv4 I__10562 (
            .O(N__48424),
            .I(\serializer_mod_inst.counter_srZ0Z_2 ));
    LocalMux I__10561 (
            .O(N__48421),
            .I(\serializer_mod_inst.counter_srZ0Z_2 ));
    InMux I__10560 (
            .O(N__48414),
            .I(\serializer_mod_inst.counter_sr_cry_1 ));
    InMux I__10559 (
            .O(N__48411),
            .I(N__48406));
    InMux I__10558 (
            .O(N__48410),
            .I(N__48401));
    InMux I__10557 (
            .O(N__48409),
            .I(N__48401));
    LocalMux I__10556 (
            .O(N__48406),
            .I(\serializer_mod_inst.counter_srZ0Z_3 ));
    LocalMux I__10555 (
            .O(N__48401),
            .I(\serializer_mod_inst.counter_srZ0Z_3 ));
    InMux I__10554 (
            .O(N__48396),
            .I(\serializer_mod_inst.counter_sr_cry_2 ));
    InMux I__10553 (
            .O(N__48393),
            .I(N__48388));
    InMux I__10552 (
            .O(N__48392),
            .I(N__48383));
    InMux I__10551 (
            .O(N__48391),
            .I(N__48383));
    LocalMux I__10550 (
            .O(N__48388),
            .I(\serializer_mod_inst.counter_srZ0Z_4 ));
    LocalMux I__10549 (
            .O(N__48383),
            .I(\serializer_mod_inst.counter_srZ0Z_4 ));
    InMux I__10548 (
            .O(N__48378),
            .I(\serializer_mod_inst.counter_sr_cry_3 ));
    InMux I__10547 (
            .O(N__48375),
            .I(N__48370));
    InMux I__10546 (
            .O(N__48374),
            .I(N__48365));
    InMux I__10545 (
            .O(N__48373),
            .I(N__48365));
    LocalMux I__10544 (
            .O(N__48370),
            .I(\serializer_mod_inst.counter_srZ0Z_5 ));
    LocalMux I__10543 (
            .O(N__48365),
            .I(\serializer_mod_inst.counter_srZ0Z_5 ));
    InMux I__10542 (
            .O(N__48360),
            .I(\serializer_mod_inst.counter_sr_cry_4 ));
    InMux I__10541 (
            .O(N__48357),
            .I(N__48352));
    CascadeMux I__10540 (
            .O(N__48356),
            .I(N__48349));
    InMux I__10539 (
            .O(N__48355),
            .I(N__48346));
    LocalMux I__10538 (
            .O(N__48352),
            .I(N__48343));
    InMux I__10537 (
            .O(N__48349),
            .I(N__48340));
    LocalMux I__10536 (
            .O(N__48346),
            .I(\serializer_mod_inst.counter_srZ0Z_6 ));
    Odrv4 I__10535 (
            .O(N__48343),
            .I(\serializer_mod_inst.counter_srZ0Z_6 ));
    LocalMux I__10534 (
            .O(N__48340),
            .I(\serializer_mod_inst.counter_srZ0Z_6 ));
    InMux I__10533 (
            .O(N__48333),
            .I(\serializer_mod_inst.counter_sr_cry_5 ));
    CascadeMux I__10532 (
            .O(N__48330),
            .I(N__48326));
    InMux I__10531 (
            .O(N__48329),
            .I(N__48322));
    InMux I__10530 (
            .O(N__48326),
            .I(N__48317));
    InMux I__10529 (
            .O(N__48325),
            .I(N__48317));
    LocalMux I__10528 (
            .O(N__48322),
            .I(N__48314));
    LocalMux I__10527 (
            .O(N__48317),
            .I(N__48311));
    Span12Mux_v I__10526 (
            .O(N__48314),
            .I(N__48307));
    Span4Mux_h I__10525 (
            .O(N__48311),
            .I(N__48304));
    InMux I__10524 (
            .O(N__48310),
            .I(N__48301));
    Odrv12 I__10523 (
            .O(N__48307),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0 ));
    Odrv4 I__10522 (
            .O(N__48304),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0 ));
    LocalMux I__10521 (
            .O(N__48301),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0 ));
    InMux I__10520 (
            .O(N__48294),
            .I(N__48287));
    InMux I__10519 (
            .O(N__48293),
            .I(N__48284));
    InMux I__10518 (
            .O(N__48292),
            .I(N__48281));
    InMux I__10517 (
            .O(N__48291),
            .I(N__48278));
    InMux I__10516 (
            .O(N__48290),
            .I(N__48275));
    LocalMux I__10515 (
            .O(N__48287),
            .I(N__48272));
    LocalMux I__10514 (
            .O(N__48284),
            .I(N__48263));
    LocalMux I__10513 (
            .O(N__48281),
            .I(N__48263));
    LocalMux I__10512 (
            .O(N__48278),
            .I(N__48263));
    LocalMux I__10511 (
            .O(N__48275),
            .I(N__48263));
    Span4Mux_v I__10510 (
            .O(N__48272),
            .I(N__48259));
    Span4Mux_v I__10509 (
            .O(N__48263),
            .I(N__48253));
    InMux I__10508 (
            .O(N__48262),
            .I(N__48250));
    Span4Mux_h I__10507 (
            .O(N__48259),
            .I(N__48247));
    InMux I__10506 (
            .O(N__48258),
            .I(N__48244));
    InMux I__10505 (
            .O(N__48257),
            .I(N__48241));
    InMux I__10504 (
            .O(N__48256),
            .I(N__48238));
    Span4Mux_h I__10503 (
            .O(N__48253),
            .I(N__48235));
    LocalMux I__10502 (
            .O(N__48250),
            .I(\I2C_top_level_inst1.s_data_ireg_0 ));
    Odrv4 I__10501 (
            .O(N__48247),
            .I(\I2C_top_level_inst1.s_data_ireg_0 ));
    LocalMux I__10500 (
            .O(N__48244),
            .I(\I2C_top_level_inst1.s_data_ireg_0 ));
    LocalMux I__10499 (
            .O(N__48241),
            .I(\I2C_top_level_inst1.s_data_ireg_0 ));
    LocalMux I__10498 (
            .O(N__48238),
            .I(\I2C_top_level_inst1.s_data_ireg_0 ));
    Odrv4 I__10497 (
            .O(N__48235),
            .I(\I2C_top_level_inst1.s_data_ireg_0 ));
    CascadeMux I__10496 (
            .O(N__48222),
            .I(N__48216));
    CascadeMux I__10495 (
            .O(N__48221),
            .I(N__48213));
    CascadeMux I__10494 (
            .O(N__48220),
            .I(N__48210));
    CascadeMux I__10493 (
            .O(N__48219),
            .I(N__48206));
    InMux I__10492 (
            .O(N__48216),
            .I(N__48196));
    InMux I__10491 (
            .O(N__48213),
            .I(N__48196));
    InMux I__10490 (
            .O(N__48210),
            .I(N__48196));
    InMux I__10489 (
            .O(N__48209),
            .I(N__48196));
    InMux I__10488 (
            .O(N__48206),
            .I(N__48190));
    InMux I__10487 (
            .O(N__48205),
            .I(N__48190));
    LocalMux I__10486 (
            .O(N__48196),
            .I(N__48187));
    InMux I__10485 (
            .O(N__48195),
            .I(N__48184));
    LocalMux I__10484 (
            .O(N__48190),
            .I(N__48174));
    Span4Mux_h I__10483 (
            .O(N__48187),
            .I(N__48174));
    LocalMux I__10482 (
            .O(N__48184),
            .I(N__48174));
    InMux I__10481 (
            .O(N__48183),
            .I(N__48167));
    InMux I__10480 (
            .O(N__48182),
            .I(N__48167));
    InMux I__10479 (
            .O(N__48181),
            .I(N__48167));
    Odrv4 I__10478 (
            .O(N__48174),
            .I(\I2C_top_level_inst1.s_command_0 ));
    LocalMux I__10477 (
            .O(N__48167),
            .I(\I2C_top_level_inst1.s_command_0 ));
    InMux I__10476 (
            .O(N__48162),
            .I(N__48159));
    LocalMux I__10475 (
            .O(N__48159),
            .I(N__48153));
    InMux I__10474 (
            .O(N__48158),
            .I(N__48150));
    InMux I__10473 (
            .O(N__48157),
            .I(N__48147));
    InMux I__10472 (
            .O(N__48156),
            .I(N__48144));
    Span4Mux_v I__10471 (
            .O(N__48153),
            .I(N__48141));
    LocalMux I__10470 (
            .O(N__48150),
            .I(N__48133));
    LocalMux I__10469 (
            .O(N__48147),
            .I(N__48133));
    LocalMux I__10468 (
            .O(N__48144),
            .I(N__48133));
    Span4Mux_h I__10467 (
            .O(N__48141),
            .I(N__48129));
    InMux I__10466 (
            .O(N__48140),
            .I(N__48126));
    Span4Mux_v I__10465 (
            .O(N__48133),
            .I(N__48123));
    InMux I__10464 (
            .O(N__48132),
            .I(N__48120));
    Odrv4 I__10463 (
            .O(N__48129),
            .I(\I2C_top_level_inst1.s_data_ireg_1 ));
    LocalMux I__10462 (
            .O(N__48126),
            .I(\I2C_top_level_inst1.s_data_ireg_1 ));
    Odrv4 I__10461 (
            .O(N__48123),
            .I(\I2C_top_level_inst1.s_data_ireg_1 ));
    LocalMux I__10460 (
            .O(N__48120),
            .I(\I2C_top_level_inst1.s_data_ireg_1 ));
    InMux I__10459 (
            .O(N__48111),
            .I(N__48108));
    LocalMux I__10458 (
            .O(N__48108),
            .I(N__48102));
    InMux I__10457 (
            .O(N__48107),
            .I(N__48099));
    InMux I__10456 (
            .O(N__48106),
            .I(N__48096));
    InMux I__10455 (
            .O(N__48105),
            .I(N__48093));
    Span4Mux_v I__10454 (
            .O(N__48102),
            .I(N__48090));
    LocalMux I__10453 (
            .O(N__48099),
            .I(N__48085));
    LocalMux I__10452 (
            .O(N__48096),
            .I(N__48085));
    LocalMux I__10451 (
            .O(N__48093),
            .I(N__48082));
    Span4Mux_h I__10450 (
            .O(N__48090),
            .I(N__48077));
    Span4Mux_v I__10449 (
            .O(N__48085),
            .I(N__48074));
    Span4Mux_v I__10448 (
            .O(N__48082),
            .I(N__48071));
    InMux I__10447 (
            .O(N__48081),
            .I(N__48066));
    InMux I__10446 (
            .O(N__48080),
            .I(N__48066));
    Odrv4 I__10445 (
            .O(N__48077),
            .I(\I2C_top_level_inst1.s_data_ireg_2 ));
    Odrv4 I__10444 (
            .O(N__48074),
            .I(\I2C_top_level_inst1.s_data_ireg_2 ));
    Odrv4 I__10443 (
            .O(N__48071),
            .I(\I2C_top_level_inst1.s_data_ireg_2 ));
    LocalMux I__10442 (
            .O(N__48066),
            .I(\I2C_top_level_inst1.s_data_ireg_2 ));
    InMux I__10441 (
            .O(N__48057),
            .I(N__48053));
    InMux I__10440 (
            .O(N__48056),
            .I(N__48050));
    LocalMux I__10439 (
            .O(N__48053),
            .I(N__48045));
    LocalMux I__10438 (
            .O(N__48050),
            .I(N__48042));
    InMux I__10437 (
            .O(N__48049),
            .I(N__48039));
    InMux I__10436 (
            .O(N__48048),
            .I(N__48036));
    Span4Mux_v I__10435 (
            .O(N__48045),
            .I(N__48033));
    Span4Mux_v I__10434 (
            .O(N__48042),
            .I(N__48029));
    LocalMux I__10433 (
            .O(N__48039),
            .I(N__48024));
    LocalMux I__10432 (
            .O(N__48036),
            .I(N__48024));
    Span4Mux_v I__10431 (
            .O(N__48033),
            .I(N__48021));
    InMux I__10430 (
            .O(N__48032),
            .I(N__48017));
    Span4Mux_h I__10429 (
            .O(N__48029),
            .I(N__48014));
    Span4Mux_v I__10428 (
            .O(N__48024),
            .I(N__48009));
    Span4Mux_h I__10427 (
            .O(N__48021),
            .I(N__48009));
    InMux I__10426 (
            .O(N__48020),
            .I(N__48006));
    LocalMux I__10425 (
            .O(N__48017),
            .I(\I2C_top_level_inst1.s_data_ireg_3 ));
    Odrv4 I__10424 (
            .O(N__48014),
            .I(\I2C_top_level_inst1.s_data_ireg_3 ));
    Odrv4 I__10423 (
            .O(N__48009),
            .I(\I2C_top_level_inst1.s_data_ireg_3 ));
    LocalMux I__10422 (
            .O(N__48006),
            .I(\I2C_top_level_inst1.s_data_ireg_3 ));
    ClkMux I__10421 (
            .O(N__47997),
            .I(N__47937));
    ClkMux I__10420 (
            .O(N__47996),
            .I(N__47937));
    ClkMux I__10419 (
            .O(N__47995),
            .I(N__47937));
    ClkMux I__10418 (
            .O(N__47994),
            .I(N__47937));
    ClkMux I__10417 (
            .O(N__47993),
            .I(N__47937));
    ClkMux I__10416 (
            .O(N__47992),
            .I(N__47937));
    ClkMux I__10415 (
            .O(N__47991),
            .I(N__47937));
    ClkMux I__10414 (
            .O(N__47990),
            .I(N__47937));
    ClkMux I__10413 (
            .O(N__47989),
            .I(N__47937));
    ClkMux I__10412 (
            .O(N__47988),
            .I(N__47937));
    ClkMux I__10411 (
            .O(N__47987),
            .I(N__47937));
    ClkMux I__10410 (
            .O(N__47986),
            .I(N__47937));
    ClkMux I__10409 (
            .O(N__47985),
            .I(N__47937));
    ClkMux I__10408 (
            .O(N__47984),
            .I(N__47937));
    ClkMux I__10407 (
            .O(N__47983),
            .I(N__47937));
    ClkMux I__10406 (
            .O(N__47982),
            .I(N__47937));
    ClkMux I__10405 (
            .O(N__47981),
            .I(N__47937));
    ClkMux I__10404 (
            .O(N__47980),
            .I(N__47937));
    ClkMux I__10403 (
            .O(N__47979),
            .I(N__47937));
    ClkMux I__10402 (
            .O(N__47978),
            .I(N__47937));
    GlobalMux I__10401 (
            .O(N__47937),
            .I(N__47934));
    gio2CtrlBuf I__10400 (
            .O(N__47934),
            .I(scl_c_g));
    CEMux I__10399 (
            .O(N__47931),
            .I(N__47928));
    LocalMux I__10398 (
            .O(N__47928),
            .I(N__47925));
    Span4Mux_h I__10397 (
            .O(N__47925),
            .I(N__47922));
    Span4Mux_h I__10396 (
            .O(N__47922),
            .I(N__47918));
    CEMux I__10395 (
            .O(N__47921),
            .I(N__47915));
    Sp12to4 I__10394 (
            .O(N__47918),
            .I(N__47907));
    LocalMux I__10393 (
            .O(N__47915),
            .I(N__47907));
    InMux I__10392 (
            .O(N__47914),
            .I(N__47904));
    InMux I__10391 (
            .O(N__47913),
            .I(N__47899));
    InMux I__10390 (
            .O(N__47912),
            .I(N__47899));
    Odrv12 I__10389 (
            .O(N__47907),
            .I(\I2C_top_level_inst1.s_load_command ));
    LocalMux I__10388 (
            .O(N__47904),
            .I(\I2C_top_level_inst1.s_load_command ));
    LocalMux I__10387 (
            .O(N__47899),
            .I(\I2C_top_level_inst1.s_load_command ));
    InMux I__10386 (
            .O(N__47892),
            .I(N__47889));
    LocalMux I__10385 (
            .O(N__47889),
            .I(\serializer_mod_inst.un1_counter_srlto6_3 ));
    CascadeMux I__10384 (
            .O(N__47886),
            .I(\serializer_mod_inst.un1_counter_srlto6_4_cascade_ ));
    InMux I__10383 (
            .O(N__47883),
            .I(N__47860));
    InMux I__10382 (
            .O(N__47882),
            .I(N__47833));
    InMux I__10381 (
            .O(N__47881),
            .I(N__47833));
    InMux I__10380 (
            .O(N__47880),
            .I(N__47833));
    InMux I__10379 (
            .O(N__47879),
            .I(N__47833));
    InMux I__10378 (
            .O(N__47878),
            .I(N__47828));
    InMux I__10377 (
            .O(N__47877),
            .I(N__47828));
    InMux I__10376 (
            .O(N__47876),
            .I(N__47823));
    InMux I__10375 (
            .O(N__47875),
            .I(N__47823));
    InMux I__10374 (
            .O(N__47874),
            .I(N__47820));
    InMux I__10373 (
            .O(N__47873),
            .I(N__47815));
    InMux I__10372 (
            .O(N__47872),
            .I(N__47815));
    InMux I__10371 (
            .O(N__47871),
            .I(N__47803));
    InMux I__10370 (
            .O(N__47870),
            .I(N__47803));
    InMux I__10369 (
            .O(N__47869),
            .I(N__47803));
    InMux I__10368 (
            .O(N__47868),
            .I(N__47798));
    InMux I__10367 (
            .O(N__47867),
            .I(N__47798));
    InMux I__10366 (
            .O(N__47866),
            .I(N__47795));
    InMux I__10365 (
            .O(N__47865),
            .I(N__47788));
    InMux I__10364 (
            .O(N__47864),
            .I(N__47788));
    InMux I__10363 (
            .O(N__47863),
            .I(N__47788));
    LocalMux I__10362 (
            .O(N__47860),
            .I(N__47785));
    InMux I__10361 (
            .O(N__47859),
            .I(N__47778));
    InMux I__10360 (
            .O(N__47858),
            .I(N__47778));
    InMux I__10359 (
            .O(N__47857),
            .I(N__47778));
    InMux I__10358 (
            .O(N__47856),
            .I(N__47771));
    InMux I__10357 (
            .O(N__47855),
            .I(N__47771));
    InMux I__10356 (
            .O(N__47854),
            .I(N__47771));
    InMux I__10355 (
            .O(N__47853),
            .I(N__47764));
    InMux I__10354 (
            .O(N__47852),
            .I(N__47764));
    InMux I__10353 (
            .O(N__47851),
            .I(N__47764));
    InMux I__10352 (
            .O(N__47850),
            .I(N__47759));
    InMux I__10351 (
            .O(N__47849),
            .I(N__47759));
    InMux I__10350 (
            .O(N__47848),
            .I(N__47756));
    InMux I__10349 (
            .O(N__47847),
            .I(N__47743));
    InMux I__10348 (
            .O(N__47846),
            .I(N__47743));
    InMux I__10347 (
            .O(N__47845),
            .I(N__47743));
    InMux I__10346 (
            .O(N__47844),
            .I(N__47743));
    InMux I__10345 (
            .O(N__47843),
            .I(N__47743));
    InMux I__10344 (
            .O(N__47842),
            .I(N__47743));
    LocalMux I__10343 (
            .O(N__47833),
            .I(N__47732));
    LocalMux I__10342 (
            .O(N__47828),
            .I(N__47732));
    LocalMux I__10341 (
            .O(N__47823),
            .I(N__47732));
    LocalMux I__10340 (
            .O(N__47820),
            .I(N__47732));
    LocalMux I__10339 (
            .O(N__47815),
            .I(N__47721));
    InMux I__10338 (
            .O(N__47814),
            .I(N__47716));
    InMux I__10337 (
            .O(N__47813),
            .I(N__47716));
    InMux I__10336 (
            .O(N__47812),
            .I(N__47711));
    InMux I__10335 (
            .O(N__47811),
            .I(N__47711));
    InMux I__10334 (
            .O(N__47810),
            .I(N__47708));
    LocalMux I__10333 (
            .O(N__47803),
            .I(N__47703));
    LocalMux I__10332 (
            .O(N__47798),
            .I(N__47696));
    LocalMux I__10331 (
            .O(N__47795),
            .I(N__47696));
    LocalMux I__10330 (
            .O(N__47788),
            .I(N__47696));
    Span4Mux_h I__10329 (
            .O(N__47785),
            .I(N__47681));
    LocalMux I__10328 (
            .O(N__47778),
            .I(N__47681));
    LocalMux I__10327 (
            .O(N__47771),
            .I(N__47681));
    LocalMux I__10326 (
            .O(N__47764),
            .I(N__47681));
    LocalMux I__10325 (
            .O(N__47759),
            .I(N__47681));
    LocalMux I__10324 (
            .O(N__47756),
            .I(N__47681));
    LocalMux I__10323 (
            .O(N__47743),
            .I(N__47681));
    InMux I__10322 (
            .O(N__47742),
            .I(N__47676));
    InMux I__10321 (
            .O(N__47741),
            .I(N__47676));
    Span4Mux_v I__10320 (
            .O(N__47732),
            .I(N__47673));
    InMux I__10319 (
            .O(N__47731),
            .I(N__47664));
    InMux I__10318 (
            .O(N__47730),
            .I(N__47664));
    InMux I__10317 (
            .O(N__47729),
            .I(N__47664));
    InMux I__10316 (
            .O(N__47728),
            .I(N__47664));
    InMux I__10315 (
            .O(N__47727),
            .I(N__47655));
    InMux I__10314 (
            .O(N__47726),
            .I(N__47655));
    InMux I__10313 (
            .O(N__47725),
            .I(N__47655));
    InMux I__10312 (
            .O(N__47724),
            .I(N__47655));
    Span4Mux_h I__10311 (
            .O(N__47721),
            .I(N__47639));
    LocalMux I__10310 (
            .O(N__47716),
            .I(N__47639));
    LocalMux I__10309 (
            .O(N__47711),
            .I(N__47634));
    LocalMux I__10308 (
            .O(N__47708),
            .I(N__47634));
    InMux I__10307 (
            .O(N__47707),
            .I(N__47629));
    InMux I__10306 (
            .O(N__47706),
            .I(N__47629));
    Span4Mux_h I__10305 (
            .O(N__47703),
            .I(N__47620));
    Span4Mux_v I__10304 (
            .O(N__47696),
            .I(N__47620));
    Span4Mux_v I__10303 (
            .O(N__47681),
            .I(N__47620));
    LocalMux I__10302 (
            .O(N__47676),
            .I(N__47620));
    Span4Mux_h I__10301 (
            .O(N__47673),
            .I(N__47613));
    LocalMux I__10300 (
            .O(N__47664),
            .I(N__47613));
    LocalMux I__10299 (
            .O(N__47655),
            .I(N__47613));
    InMux I__10298 (
            .O(N__47654),
            .I(N__47602));
    InMux I__10297 (
            .O(N__47653),
            .I(N__47602));
    InMux I__10296 (
            .O(N__47652),
            .I(N__47602));
    InMux I__10295 (
            .O(N__47651),
            .I(N__47602));
    InMux I__10294 (
            .O(N__47650),
            .I(N__47602));
    InMux I__10293 (
            .O(N__47649),
            .I(N__47591));
    InMux I__10292 (
            .O(N__47648),
            .I(N__47591));
    InMux I__10291 (
            .O(N__47647),
            .I(N__47591));
    InMux I__10290 (
            .O(N__47646),
            .I(N__47591));
    InMux I__10289 (
            .O(N__47645),
            .I(N__47591));
    InMux I__10288 (
            .O(N__47644),
            .I(N__47588));
    Odrv4 I__10287 (
            .O(N__47639),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    Odrv12 I__10286 (
            .O(N__47634),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    LocalMux I__10285 (
            .O(N__47629),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    Odrv4 I__10284 (
            .O(N__47620),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    Odrv4 I__10283 (
            .O(N__47613),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    LocalMux I__10282 (
            .O(N__47602),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    LocalMux I__10281 (
            .O(N__47591),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    LocalMux I__10280 (
            .O(N__47588),
            .I(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ));
    CascadeMux I__10279 (
            .O(N__47571),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_10_cascade_ ));
    CascadeMux I__10278 (
            .O(N__47568),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_18_cascade_ ));
    InMux I__10277 (
            .O(N__47565),
            .I(N__47557));
    InMux I__10276 (
            .O(N__47564),
            .I(N__47557));
    InMux I__10275 (
            .O(N__47563),
            .I(N__47552));
    InMux I__10274 (
            .O(N__47562),
            .I(N__47552));
    LocalMux I__10273 (
            .O(N__47557),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18 ));
    LocalMux I__10272 (
            .O(N__47552),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18 ));
    InMux I__10271 (
            .O(N__47547),
            .I(N__47538));
    InMux I__10270 (
            .O(N__47546),
            .I(N__47538));
    InMux I__10269 (
            .O(N__47545),
            .I(N__47538));
    LocalMux I__10268 (
            .O(N__47538),
            .I(N__47535));
    Span4Mux_h I__10267 (
            .O(N__47535),
            .I(N__47532));
    Span4Mux_v I__10266 (
            .O(N__47532),
            .I(N__47529));
    Odrv4 I__10265 (
            .O(N__47529),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1605_0 ));
    InMux I__10264 (
            .O(N__47526),
            .I(N__47523));
    LocalMux I__10263 (
            .O(N__47523),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0 ));
    CascadeMux I__10262 (
            .O(N__47520),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0_cascade_ ));
    InMux I__10261 (
            .O(N__47517),
            .I(N__47514));
    LocalMux I__10260 (
            .O(N__47514),
            .I(N__47511));
    Span4Mux_v I__10259 (
            .O(N__47511),
            .I(N__47507));
    InMux I__10258 (
            .O(N__47510),
            .I(N__47504));
    Span4Mux_v I__10257 (
            .O(N__47507),
            .I(N__47501));
    LocalMux I__10256 (
            .O(N__47504),
            .I(N__47498));
    Odrv4 I__10255 (
            .O(N__47501),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0 ));
    Odrv4 I__10254 (
            .O(N__47498),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0 ));
    InMux I__10253 (
            .O(N__47493),
            .I(N__47490));
    LocalMux I__10252 (
            .O(N__47490),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_0_1_14 ));
    CascadeMux I__10251 (
            .O(N__47487),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_279_cascade_ ));
    CascadeMux I__10250 (
            .O(N__47484),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_0_1_7_cascade_ ));
    CascadeMux I__10249 (
            .O(N__47481),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_268_cascade_ ));
    InMux I__10248 (
            .O(N__47478),
            .I(N__47475));
    LocalMux I__10247 (
            .O(N__47475),
            .I(N__47472));
    Odrv4 I__10246 (
            .O(N__47472),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_7_3_i_a2_0 ));
    InMux I__10245 (
            .O(N__47469),
            .I(N__47463));
    InMux I__10244 (
            .O(N__47468),
            .I(N__47463));
    LocalMux I__10243 (
            .O(N__47463),
            .I(N__47460));
    Span4Mux_h I__10242 (
            .O(N__47460),
            .I(N__47457));
    Span4Mux_h I__10241 (
            .O(N__47457),
            .I(N__47453));
    InMux I__10240 (
            .O(N__47456),
            .I(N__47450));
    Odrv4 I__10239 (
            .O(N__47453),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0 ));
    LocalMux I__10238 (
            .O(N__47450),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0 ));
    InMux I__10237 (
            .O(N__47445),
            .I(N__47442));
    LocalMux I__10236 (
            .O(N__47442),
            .I(N__47439));
    Odrv12 I__10235 (
            .O(N__47439),
            .I(\I2C_top_level_inst1.s_addr1_o_0 ));
    CascadeMux I__10234 (
            .O(N__47436),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0_cascade_ ));
    InMux I__10233 (
            .O(N__47433),
            .I(N__47430));
    LocalMux I__10232 (
            .O(N__47430),
            .I(N__47427));
    Span4Mux_h I__10231 (
            .O(N__47427),
            .I(N__47423));
    InMux I__10230 (
            .O(N__47426),
            .I(N__47420));
    Odrv4 I__10229 (
            .O(N__47423),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1 ));
    LocalMux I__10228 (
            .O(N__47420),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1 ));
    InMux I__10227 (
            .O(N__47415),
            .I(N__47404));
    InMux I__10226 (
            .O(N__47414),
            .I(N__47404));
    InMux I__10225 (
            .O(N__47413),
            .I(N__47400));
    InMux I__10224 (
            .O(N__47412),
            .I(N__47391));
    InMux I__10223 (
            .O(N__47411),
            .I(N__47391));
    InMux I__10222 (
            .O(N__47410),
            .I(N__47391));
    InMux I__10221 (
            .O(N__47409),
            .I(N__47391));
    LocalMux I__10220 (
            .O(N__47404),
            .I(N__47388));
    CascadeMux I__10219 (
            .O(N__47403),
            .I(N__47385));
    LocalMux I__10218 (
            .O(N__47400),
            .I(N__47375));
    LocalMux I__10217 (
            .O(N__47391),
            .I(N__47372));
    Span4Mux_h I__10216 (
            .O(N__47388),
            .I(N__47369));
    InMux I__10215 (
            .O(N__47385),
            .I(N__47366));
    InMux I__10214 (
            .O(N__47384),
            .I(N__47357));
    InMux I__10213 (
            .O(N__47383),
            .I(N__47357));
    InMux I__10212 (
            .O(N__47382),
            .I(N__47357));
    InMux I__10211 (
            .O(N__47381),
            .I(N__47357));
    InMux I__10210 (
            .O(N__47380),
            .I(N__47350));
    InMux I__10209 (
            .O(N__47379),
            .I(N__47350));
    InMux I__10208 (
            .O(N__47378),
            .I(N__47350));
    Span4Mux_h I__10207 (
            .O(N__47375),
            .I(N__47347));
    Span4Mux_h I__10206 (
            .O(N__47372),
            .I(N__47344));
    Sp12to4 I__10205 (
            .O(N__47369),
            .I(N__47341));
    LocalMux I__10204 (
            .O(N__47366),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ));
    LocalMux I__10203 (
            .O(N__47357),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ));
    LocalMux I__10202 (
            .O(N__47350),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ));
    Odrv4 I__10201 (
            .O(N__47347),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ));
    Odrv4 I__10200 (
            .O(N__47344),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ));
    Odrv12 I__10199 (
            .O(N__47341),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ));
    CascadeMux I__10198 (
            .O(N__47328),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_8_cascade_ ));
    InMux I__10197 (
            .O(N__47325),
            .I(N__47322));
    LocalMux I__10196 (
            .O(N__47322),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_CO ));
    InMux I__10195 (
            .O(N__47319),
            .I(N__47316));
    LocalMux I__10194 (
            .O(N__47316),
            .I(N__47313));
    Span4Mux_v I__10193 (
            .O(N__47313),
            .I(N__47310));
    Odrv4 I__10192 (
            .O(N__47310),
            .I(\I2C_top_level_inst1.s_addr0_o_1 ));
    CascadeMux I__10191 (
            .O(N__47307),
            .I(N__47304));
    InMux I__10190 (
            .O(N__47304),
            .I(N__47301));
    LocalMux I__10189 (
            .O(N__47301),
            .I(N__47298));
    Span4Mux_v I__10188 (
            .O(N__47298),
            .I(N__47295));
    Span4Mux_h I__10187 (
            .O(N__47295),
            .I(N__47292));
    Span4Mux_v I__10186 (
            .O(N__47292),
            .I(N__47289));
    Odrv4 I__10185 (
            .O(N__47289),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1651 ));
    InMux I__10184 (
            .O(N__47286),
            .I(N__47283));
    LocalMux I__10183 (
            .O(N__47283),
            .I(N__47280));
    Span4Mux_h I__10182 (
            .O(N__47280),
            .I(N__47277));
    Span4Mux_h I__10181 (
            .O(N__47277),
            .I(N__47274));
    Odrv4 I__10180 (
            .O(N__47274),
            .I(\I2C_top_level_inst1.s_addr0_o_2 ));
    CascadeMux I__10179 (
            .O(N__47271),
            .I(N__47268));
    InMux I__10178 (
            .O(N__47268),
            .I(N__47265));
    LocalMux I__10177 (
            .O(N__47265),
            .I(N__47262));
    Span4Mux_h I__10176 (
            .O(N__47262),
            .I(N__47259));
    Sp12to4 I__10175 (
            .O(N__47259),
            .I(N__47256));
    Span12Mux_v I__10174 (
            .O(N__47256),
            .I(N__47253));
    Odrv12 I__10173 (
            .O(N__47253),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1652 ));
    CascadeMux I__10172 (
            .O(N__47250),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_0_4_cascade_ ));
    InMux I__10171 (
            .O(N__47247),
            .I(N__47240));
    InMux I__10170 (
            .O(N__47246),
            .I(N__47237));
    InMux I__10169 (
            .O(N__47245),
            .I(N__47232));
    InMux I__10168 (
            .O(N__47244),
            .I(N__47232));
    InMux I__10167 (
            .O(N__47243),
            .I(N__47229));
    LocalMux I__10166 (
            .O(N__47240),
            .I(N__47222));
    LocalMux I__10165 (
            .O(N__47237),
            .I(N__47222));
    LocalMux I__10164 (
            .O(N__47232),
            .I(N__47222));
    LocalMux I__10163 (
            .O(N__47229),
            .I(N__47219));
    Span4Mux_h I__10162 (
            .O(N__47222),
            .I(N__47216));
    Span4Mux_v I__10161 (
            .O(N__47219),
            .I(N__47213));
    Odrv4 I__10160 (
            .O(N__47216),
            .I(s_paddr_I2C_5));
    Odrv4 I__10159 (
            .O(N__47213),
            .I(s_paddr_I2C_5));
    InMux I__10158 (
            .O(N__47208),
            .I(N__47201));
    InMux I__10157 (
            .O(N__47207),
            .I(N__47201));
    InMux I__10156 (
            .O(N__47206),
            .I(N__47198));
    LocalMux I__10155 (
            .O(N__47201),
            .I(N__47193));
    LocalMux I__10154 (
            .O(N__47198),
            .I(N__47190));
    InMux I__10153 (
            .O(N__47197),
            .I(N__47187));
    InMux I__10152 (
            .O(N__47196),
            .I(N__47184));
    Span4Mux_v I__10151 (
            .O(N__47193),
            .I(N__47179));
    Span4Mux_v I__10150 (
            .O(N__47190),
            .I(N__47179));
    LocalMux I__10149 (
            .O(N__47187),
            .I(s_paddr_I2C_4));
    LocalMux I__10148 (
            .O(N__47184),
            .I(s_paddr_I2C_4));
    Odrv4 I__10147 (
            .O(N__47179),
            .I(s_paddr_I2C_4));
    InMux I__10146 (
            .O(N__47172),
            .I(N__47165));
    InMux I__10145 (
            .O(N__47171),
            .I(N__47161));
    InMux I__10144 (
            .O(N__47170),
            .I(N__47158));
    InMux I__10143 (
            .O(N__47169),
            .I(N__47153));
    InMux I__10142 (
            .O(N__47168),
            .I(N__47153));
    LocalMux I__10141 (
            .O(N__47165),
            .I(N__47150));
    InMux I__10140 (
            .O(N__47164),
            .I(N__47147));
    LocalMux I__10139 (
            .O(N__47161),
            .I(N__47140));
    LocalMux I__10138 (
            .O(N__47158),
            .I(N__47140));
    LocalMux I__10137 (
            .O(N__47153),
            .I(N__47140));
    Span4Mux_v I__10136 (
            .O(N__47150),
            .I(N__47137));
    LocalMux I__10135 (
            .O(N__47147),
            .I(N__47134));
    Span4Mux_v I__10134 (
            .O(N__47140),
            .I(N__47129));
    Span4Mux_h I__10133 (
            .O(N__47137),
            .I(N__47129));
    Odrv4 I__10132 (
            .O(N__47134),
            .I(s_paddr_I2C_6));
    Odrv4 I__10131 (
            .O(N__47129),
            .I(s_paddr_I2C_6));
    CascadeMux I__10130 (
            .O(N__47124),
            .I(N__47119));
    CascadeMux I__10129 (
            .O(N__47123),
            .I(N__47115));
    CascadeMux I__10128 (
            .O(N__47122),
            .I(N__47112));
    InMux I__10127 (
            .O(N__47119),
            .I(N__47107));
    InMux I__10126 (
            .O(N__47118),
            .I(N__47104));
    InMux I__10125 (
            .O(N__47115),
            .I(N__47099));
    InMux I__10124 (
            .O(N__47112),
            .I(N__47099));
    InMux I__10123 (
            .O(N__47111),
            .I(N__47094));
    InMux I__10122 (
            .O(N__47110),
            .I(N__47094));
    LocalMux I__10121 (
            .O(N__47107),
            .I(N__47090));
    LocalMux I__10120 (
            .O(N__47104),
            .I(N__47085));
    LocalMux I__10119 (
            .O(N__47099),
            .I(N__47085));
    LocalMux I__10118 (
            .O(N__47094),
            .I(N__47082));
    InMux I__10117 (
            .O(N__47093),
            .I(N__47079));
    Span4Mux_h I__10116 (
            .O(N__47090),
            .I(N__47076));
    Span4Mux_h I__10115 (
            .O(N__47085),
            .I(N__47073));
    Span4Mux_h I__10114 (
            .O(N__47082),
            .I(N__47068));
    LocalMux I__10113 (
            .O(N__47079),
            .I(N__47068));
    Odrv4 I__10112 (
            .O(N__47076),
            .I(s_paddr_I2C_7));
    Odrv4 I__10111 (
            .O(N__47073),
            .I(s_paddr_I2C_7));
    Odrv4 I__10110 (
            .O(N__47068),
            .I(s_paddr_I2C_7));
    InMux I__10109 (
            .O(N__47061),
            .I(N__47058));
    LocalMux I__10108 (
            .O(N__47058),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_2 ));
    InMux I__10107 (
            .O(N__47055),
            .I(N__47052));
    LocalMux I__10106 (
            .O(N__47052),
            .I(N__47049));
    Span4Mux_v I__10105 (
            .O(N__47049),
            .I(N__47046));
    Odrv4 I__10104 (
            .O(N__47046),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_5 ));
    InMux I__10103 (
            .O(N__47043),
            .I(N__47038));
    InMux I__10102 (
            .O(N__47042),
            .I(N__47034));
    InMux I__10101 (
            .O(N__47041),
            .I(N__47031));
    LocalMux I__10100 (
            .O(N__47038),
            .I(N__47028));
    InMux I__10099 (
            .O(N__47037),
            .I(N__47025));
    LocalMux I__10098 (
            .O(N__47034),
            .I(N__47018));
    LocalMux I__10097 (
            .O(N__47031),
            .I(N__47018));
    Span4Mux_v I__10096 (
            .O(N__47028),
            .I(N__47018));
    LocalMux I__10095 (
            .O(N__47025),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10 ));
    Odrv4 I__10094 (
            .O(N__47018),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10 ));
    InMux I__10093 (
            .O(N__47013),
            .I(N__47009));
    InMux I__10092 (
            .O(N__47012),
            .I(N__47004));
    LocalMux I__10091 (
            .O(N__47009),
            .I(N__47001));
    InMux I__10090 (
            .O(N__47008),
            .I(N__46998));
    InMux I__10089 (
            .O(N__47007),
            .I(N__46995));
    LocalMux I__10088 (
            .O(N__47004),
            .I(N__46992));
    Span4Mux_h I__10087 (
            .O(N__47001),
            .I(N__46989));
    LocalMux I__10086 (
            .O(N__46998),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9 ));
    LocalMux I__10085 (
            .O(N__46995),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9 ));
    Odrv4 I__10084 (
            .O(N__46992),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9 ));
    Odrv4 I__10083 (
            .O(N__46989),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9 ));
    InMux I__10082 (
            .O(N__46980),
            .I(N__46977));
    LocalMux I__10081 (
            .O(N__46977),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_3 ));
    InMux I__10080 (
            .O(N__46974),
            .I(N__46971));
    LocalMux I__10079 (
            .O(N__46971),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_2_2 ));
    CascadeMux I__10078 (
            .O(N__46968),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0_cascade_ ));
    CascadeMux I__10077 (
            .O(N__46965),
            .I(N__46962));
    InMux I__10076 (
            .O(N__46962),
            .I(N__46959));
    LocalMux I__10075 (
            .O(N__46959),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0 ));
    InMux I__10074 (
            .O(N__46956),
            .I(N__46953));
    LocalMux I__10073 (
            .O(N__46953),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_1_0 ));
    CascadeMux I__10072 (
            .O(N__46950),
            .I(N__46947));
    InMux I__10071 (
            .O(N__46947),
            .I(N__46943));
    InMux I__10070 (
            .O(N__46946),
            .I(N__46939));
    LocalMux I__10069 (
            .O(N__46943),
            .I(N__46935));
    InMux I__10068 (
            .O(N__46942),
            .I(N__46932));
    LocalMux I__10067 (
            .O(N__46939),
            .I(N__46929));
    InMux I__10066 (
            .O(N__46938),
            .I(N__46926));
    Span4Mux_h I__10065 (
            .O(N__46935),
            .I(N__46923));
    LocalMux I__10064 (
            .O(N__46932),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11 ));
    Odrv4 I__10063 (
            .O(N__46929),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11 ));
    LocalMux I__10062 (
            .O(N__46926),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11 ));
    Odrv4 I__10061 (
            .O(N__46923),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11 ));
    CascadeMux I__10060 (
            .O(N__46914),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0_cascade_ ));
    InMux I__10059 (
            .O(N__46911),
            .I(N__46904));
    CascadeMux I__10058 (
            .O(N__46910),
            .I(N__46901));
    CascadeMux I__10057 (
            .O(N__46909),
            .I(N__46897));
    CascadeMux I__10056 (
            .O(N__46908),
            .I(N__46893));
    InMux I__10055 (
            .O(N__46907),
            .I(N__46888));
    LocalMux I__10054 (
            .O(N__46904),
            .I(N__46885));
    InMux I__10053 (
            .O(N__46901),
            .I(N__46876));
    InMux I__10052 (
            .O(N__46900),
            .I(N__46876));
    InMux I__10051 (
            .O(N__46897),
            .I(N__46876));
    InMux I__10050 (
            .O(N__46896),
            .I(N__46876));
    InMux I__10049 (
            .O(N__46893),
            .I(N__46869));
    InMux I__10048 (
            .O(N__46892),
            .I(N__46869));
    InMux I__10047 (
            .O(N__46891),
            .I(N__46869));
    LocalMux I__10046 (
            .O(N__46888),
            .I(N__46866));
    Span4Mux_v I__10045 (
            .O(N__46885),
            .I(N__46863));
    LocalMux I__10044 (
            .O(N__46876),
            .I(N__46860));
    LocalMux I__10043 (
            .O(N__46869),
            .I(N__46857));
    Span4Mux_v I__10042 (
            .O(N__46866),
            .I(N__46854));
    Span4Mux_h I__10041 (
            .O(N__46863),
            .I(N__46849));
    Span4Mux_v I__10040 (
            .O(N__46860),
            .I(N__46849));
    Span4Mux_h I__10039 (
            .O(N__46857),
            .I(N__46846));
    Sp12to4 I__10038 (
            .O(N__46854),
            .I(N__46843));
    Sp12to4 I__10037 (
            .O(N__46849),
            .I(N__46840));
    Span4Mux_v I__10036 (
            .O(N__46846),
            .I(N__46837));
    Span12Mux_h I__10035 (
            .O(N__46843),
            .I(N__46832));
    Span12Mux_h I__10034 (
            .O(N__46840),
            .I(N__46832));
    Span4Mux_v I__10033 (
            .O(N__46837),
            .I(N__46829));
    Odrv12 I__10032 (
            .O(N__46832),
            .I(s_paddr_I2C_2));
    Odrv4 I__10031 (
            .O(N__46829),
            .I(s_paddr_I2C_2));
    InMux I__10030 (
            .O(N__46824),
            .I(N__46821));
    LocalMux I__10029 (
            .O(N__46821),
            .I(N__46818));
    Span4Mux_v I__10028 (
            .O(N__46818),
            .I(N__46814));
    InMux I__10027 (
            .O(N__46817),
            .I(N__46808));
    Span4Mux_h I__10026 (
            .O(N__46814),
            .I(N__46804));
    InMux I__10025 (
            .O(N__46813),
            .I(N__46799));
    InMux I__10024 (
            .O(N__46812),
            .I(N__46799));
    InMux I__10023 (
            .O(N__46811),
            .I(N__46796));
    LocalMux I__10022 (
            .O(N__46808),
            .I(N__46793));
    InMux I__10021 (
            .O(N__46807),
            .I(N__46790));
    Sp12to4 I__10020 (
            .O(N__46804),
            .I(N__46787));
    LocalMux I__10019 (
            .O(N__46799),
            .I(N__46782));
    LocalMux I__10018 (
            .O(N__46796),
            .I(N__46782));
    Span4Mux_v I__10017 (
            .O(N__46793),
            .I(N__46779));
    LocalMux I__10016 (
            .O(N__46790),
            .I(N__46772));
    Span12Mux_v I__10015 (
            .O(N__46787),
            .I(N__46772));
    Span12Mux_h I__10014 (
            .O(N__46782),
            .I(N__46772));
    Span4Mux_v I__10013 (
            .O(N__46779),
            .I(N__46769));
    Odrv12 I__10012 (
            .O(N__46772),
            .I(s_paddr_I2C_1));
    Odrv4 I__10011 (
            .O(N__46769),
            .I(s_paddr_I2C_1));
    InMux I__10010 (
            .O(N__46764),
            .I(N__46757));
    CascadeMux I__10009 (
            .O(N__46763),
            .I(N__46753));
    InMux I__10008 (
            .O(N__46762),
            .I(N__46746));
    InMux I__10007 (
            .O(N__46761),
            .I(N__46746));
    InMux I__10006 (
            .O(N__46760),
            .I(N__46746));
    LocalMux I__10005 (
            .O(N__46757),
            .I(N__46743));
    InMux I__10004 (
            .O(N__46756),
            .I(N__46740));
    InMux I__10003 (
            .O(N__46753),
            .I(N__46737));
    LocalMux I__10002 (
            .O(N__46746),
            .I(N__46732));
    Span4Mux_v I__10001 (
            .O(N__46743),
            .I(N__46732));
    LocalMux I__10000 (
            .O(N__46740),
            .I(s_paddr_I2C_0));
    LocalMux I__9999 (
            .O(N__46737),
            .I(s_paddr_I2C_0));
    Odrv4 I__9998 (
            .O(N__46732),
            .I(s_paddr_I2C_0));
    InMux I__9997 (
            .O(N__46725),
            .I(N__46722));
    LocalMux I__9996 (
            .O(N__46722),
            .I(N__46719));
    Span4Mux_v I__9995 (
            .O(N__46719),
            .I(N__46716));
    Span4Mux_h I__9994 (
            .O(N__46716),
            .I(N__46713));
    Odrv4 I__9993 (
            .O(N__46713),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_10 ));
    InMux I__9992 (
            .O(N__46710),
            .I(N__46707));
    LocalMux I__9991 (
            .O(N__46707),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_10 ));
    CascadeMux I__9990 (
            .O(N__46704),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7DZ0Z7_cascade_ ));
    InMux I__9989 (
            .O(N__46701),
            .I(N__46698));
    LocalMux I__9988 (
            .O(N__46698),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10 ));
    InMux I__9987 (
            .O(N__46695),
            .I(N__46692));
    LocalMux I__9986 (
            .O(N__46692),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_9 ));
    CascadeMux I__9985 (
            .O(N__46689),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10_cascade_ ));
    InMux I__9984 (
            .O(N__46686),
            .I(N__46683));
    LocalMux I__9983 (
            .O(N__46683),
            .I(N__46680));
    Span4Mux_h I__9982 (
            .O(N__46680),
            .I(N__46677));
    Span4Mux_v I__9981 (
            .O(N__46677),
            .I(N__46674));
    Odrv4 I__9980 (
            .O(N__46674),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_10 ));
    InMux I__9979 (
            .O(N__46671),
            .I(N__46668));
    LocalMux I__9978 (
            .O(N__46668),
            .I(N__46664));
    CascadeMux I__9977 (
            .O(N__46667),
            .I(N__46661));
    Span4Mux_v I__9976 (
            .O(N__46664),
            .I(N__46657));
    InMux I__9975 (
            .O(N__46661),
            .I(N__46654));
    InMux I__9974 (
            .O(N__46660),
            .I(N__46651));
    Span4Mux_h I__9973 (
            .O(N__46657),
            .I(N__46644));
    LocalMux I__9972 (
            .O(N__46654),
            .I(N__46644));
    LocalMux I__9971 (
            .O(N__46651),
            .I(N__46644));
    Odrv4 I__9970 (
            .O(N__46644),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_9));
    InMux I__9969 (
            .O(N__46641),
            .I(N__46638));
    LocalMux I__9968 (
            .O(N__46638),
            .I(N__46635));
    Span4Mux_h I__9967 (
            .O(N__46635),
            .I(N__46631));
    CascadeMux I__9966 (
            .O(N__46634),
            .I(N__46628));
    Span4Mux_h I__9965 (
            .O(N__46631),
            .I(N__46624));
    InMux I__9964 (
            .O(N__46628),
            .I(N__46619));
    InMux I__9963 (
            .O(N__46627),
            .I(N__46619));
    Odrv4 I__9962 (
            .O(N__46624),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_9));
    LocalMux I__9961 (
            .O(N__46619),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_9));
    InMux I__9960 (
            .O(N__46614),
            .I(N__46611));
    LocalMux I__9959 (
            .O(N__46611),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_9 ));
    CascadeMux I__9958 (
            .O(N__46608),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i_cascade_ ));
    InMux I__9957 (
            .O(N__46605),
            .I(N__46602));
    LocalMux I__9956 (
            .O(N__46602),
            .I(N__46599));
    Sp12to4 I__9955 (
            .O(N__46599),
            .I(N__46594));
    InMux I__9954 (
            .O(N__46598),
            .I(N__46589));
    InMux I__9953 (
            .O(N__46597),
            .I(N__46589));
    Span12Mux_v I__9952 (
            .O(N__46594),
            .I(N__46586));
    LocalMux I__9951 (
            .O(N__46589),
            .I(N__46583));
    Odrv12 I__9950 (
            .O(N__46586),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_15));
    Odrv4 I__9949 (
            .O(N__46583),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_15));
    InMux I__9948 (
            .O(N__46578),
            .I(N__46575));
    LocalMux I__9947 (
            .O(N__46575),
            .I(N__46572));
    Span4Mux_v I__9946 (
            .O(N__46572),
            .I(N__46569));
    Span4Mux_v I__9945 (
            .O(N__46569),
            .I(N__46566));
    Odrv4 I__9944 (
            .O(N__46566),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_24));
    InMux I__9943 (
            .O(N__46563),
            .I(N__46560));
    LocalMux I__9942 (
            .O(N__46560),
            .I(N__46557));
    Span4Mux_v I__9941 (
            .O(N__46557),
            .I(N__46553));
    CascadeMux I__9940 (
            .O(N__46556),
            .I(N__46549));
    Span4Mux_v I__9939 (
            .O(N__46553),
            .I(N__46546));
    InMux I__9938 (
            .O(N__46552),
            .I(N__46541));
    InMux I__9937 (
            .O(N__46549),
            .I(N__46541));
    Span4Mux_h I__9936 (
            .O(N__46546),
            .I(N__46538));
    LocalMux I__9935 (
            .O(N__46541),
            .I(N__46535));
    Odrv4 I__9934 (
            .O(N__46538),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_17));
    Odrv12 I__9933 (
            .O(N__46535),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_17));
    InMux I__9932 (
            .O(N__46530),
            .I(N__46527));
    LocalMux I__9931 (
            .O(N__46527),
            .I(N__46520));
    InMux I__9930 (
            .O(N__46526),
            .I(N__46517));
    InMux I__9929 (
            .O(N__46525),
            .I(N__46514));
    InMux I__9928 (
            .O(N__46524),
            .I(N__46511));
    InMux I__9927 (
            .O(N__46523),
            .I(N__46508));
    Span4Mux_v I__9926 (
            .O(N__46520),
            .I(N__46502));
    LocalMux I__9925 (
            .O(N__46517),
            .I(N__46502));
    LocalMux I__9924 (
            .O(N__46514),
            .I(N__46497));
    LocalMux I__9923 (
            .O(N__46511),
            .I(N__46494));
    LocalMux I__9922 (
            .O(N__46508),
            .I(N__46491));
    CascadeMux I__9921 (
            .O(N__46507),
            .I(N__46488));
    Span4Mux_h I__9920 (
            .O(N__46502),
            .I(N__46485));
    InMux I__9919 (
            .O(N__46501),
            .I(N__46482));
    InMux I__9918 (
            .O(N__46500),
            .I(N__46479));
    Span4Mux_v I__9917 (
            .O(N__46497),
            .I(N__46476));
    Span4Mux_v I__9916 (
            .O(N__46494),
            .I(N__46471));
    Span4Mux_h I__9915 (
            .O(N__46491),
            .I(N__46471));
    InMux I__9914 (
            .O(N__46488),
            .I(N__46468));
    Span4Mux_h I__9913 (
            .O(N__46485),
            .I(N__46465));
    LocalMux I__9912 (
            .O(N__46482),
            .I(N__46462));
    LocalMux I__9911 (
            .O(N__46479),
            .I(N__46458));
    Span4Mux_v I__9910 (
            .O(N__46476),
            .I(N__46453));
    Span4Mux_h I__9909 (
            .O(N__46471),
            .I(N__46453));
    LocalMux I__9908 (
            .O(N__46468),
            .I(N__46450));
    Span4Mux_h I__9907 (
            .O(N__46465),
            .I(N__46447));
    Span4Mux_v I__9906 (
            .O(N__46462),
            .I(N__46444));
    InMux I__9905 (
            .O(N__46461),
            .I(N__46441));
    Span12Mux_v I__9904 (
            .O(N__46458),
            .I(N__46438));
    Span4Mux_h I__9903 (
            .O(N__46453),
            .I(N__46435));
    Span4Mux_h I__9902 (
            .O(N__46450),
            .I(N__46428));
    Span4Mux_h I__9901 (
            .O(N__46447),
            .I(N__46428));
    Span4Mux_h I__9900 (
            .O(N__46444),
            .I(N__46428));
    LocalMux I__9899 (
            .O(N__46441),
            .I(I2C_top_level_inst1_s_data_oreg_9));
    Odrv12 I__9898 (
            .O(N__46438),
            .I(I2C_top_level_inst1_s_data_oreg_9));
    Odrv4 I__9897 (
            .O(N__46435),
            .I(I2C_top_level_inst1_s_data_oreg_9));
    Odrv4 I__9896 (
            .O(N__46428),
            .I(I2C_top_level_inst1_s_data_oreg_9));
    CascadeMux I__9895 (
            .O(N__46419),
            .I(N__46416));
    InMux I__9894 (
            .O(N__46416),
            .I(N__46413));
    LocalMux I__9893 (
            .O(N__46413),
            .I(N__46410));
    Span4Mux_v I__9892 (
            .O(N__46410),
            .I(N__46407));
    Odrv4 I__9891 (
            .O(N__46407),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_9 ));
    CascadeMux I__9890 (
            .O(N__46404),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSLZ0Z7_cascade_ ));
    InMux I__9889 (
            .O(N__46401),
            .I(N__46398));
    LocalMux I__9888 (
            .O(N__46398),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9 ));
    CascadeMux I__9887 (
            .O(N__46395),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9_cascade_ ));
    InMux I__9886 (
            .O(N__46392),
            .I(N__46389));
    LocalMux I__9885 (
            .O(N__46389),
            .I(N__46386));
    Span4Mux_h I__9884 (
            .O(N__46386),
            .I(N__46383));
    Odrv4 I__9883 (
            .O(N__46383),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_8 ));
    InMux I__9882 (
            .O(N__46380),
            .I(N__46377));
    LocalMux I__9881 (
            .O(N__46377),
            .I(N__46373));
    InMux I__9880 (
            .O(N__46376),
            .I(N__46370));
    Span4Mux_v I__9879 (
            .O(N__46373),
            .I(N__46366));
    LocalMux I__9878 (
            .O(N__46370),
            .I(N__46363));
    InMux I__9877 (
            .O(N__46369),
            .I(N__46360));
    Span4Mux_h I__9876 (
            .O(N__46366),
            .I(N__46355));
    Span4Mux_v I__9875 (
            .O(N__46363),
            .I(N__46355));
    LocalMux I__9874 (
            .O(N__46360),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_11));
    Odrv4 I__9873 (
            .O(N__46355),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_11));
    InMux I__9872 (
            .O(N__46350),
            .I(N__46347));
    LocalMux I__9871 (
            .O(N__46347),
            .I(N__46343));
    InMux I__9870 (
            .O(N__46346),
            .I(N__46340));
    Span4Mux_v I__9869 (
            .O(N__46343),
            .I(N__46336));
    LocalMux I__9868 (
            .O(N__46340),
            .I(N__46333));
    InMux I__9867 (
            .O(N__46339),
            .I(N__46330));
    Span4Mux_h I__9866 (
            .O(N__46336),
            .I(N__46327));
    Span4Mux_v I__9865 (
            .O(N__46333),
            .I(N__46322));
    LocalMux I__9864 (
            .O(N__46330),
            .I(N__46322));
    Odrv4 I__9863 (
            .O(N__46327),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_12));
    Odrv4 I__9862 (
            .O(N__46322),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_12));
    InMux I__9861 (
            .O(N__46317),
            .I(N__46314));
    LocalMux I__9860 (
            .O(N__46314),
            .I(N__46311));
    Span4Mux_h I__9859 (
            .O(N__46311),
            .I(N__46308));
    Span4Mux_h I__9858 (
            .O(N__46308),
            .I(N__46303));
    InMux I__9857 (
            .O(N__46307),
            .I(N__46298));
    InMux I__9856 (
            .O(N__46306),
            .I(N__46298));
    Odrv4 I__9855 (
            .O(N__46303),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_21));
    LocalMux I__9854 (
            .O(N__46298),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_21));
    CascadeMux I__9853 (
            .O(N__46293),
            .I(N__46290));
    InMux I__9852 (
            .O(N__46290),
            .I(N__46287));
    LocalMux I__9851 (
            .O(N__46287),
            .I(N__46284));
    Span4Mux_h I__9850 (
            .O(N__46284),
            .I(N__46281));
    Span4Mux_h I__9849 (
            .O(N__46281),
            .I(N__46278));
    Span4Mux_h I__9848 (
            .O(N__46278),
            .I(N__46275));
    Odrv4 I__9847 (
            .O(N__46275),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_30));
    InMux I__9846 (
            .O(N__46272),
            .I(N__46267));
    InMux I__9845 (
            .O(N__46271),
            .I(N__46264));
    InMux I__9844 (
            .O(N__46270),
            .I(N__46261));
    LocalMux I__9843 (
            .O(N__46267),
            .I(N__46258));
    LocalMux I__9842 (
            .O(N__46264),
            .I(N__46255));
    LocalMux I__9841 (
            .O(N__46261),
            .I(N__46252));
    Span4Mux_v I__9840 (
            .O(N__46258),
            .I(N__46249));
    Span4Mux_h I__9839 (
            .O(N__46255),
            .I(N__46246));
    Span4Mux_h I__9838 (
            .O(N__46252),
            .I(N__46243));
    Span4Mux_h I__9837 (
            .O(N__46249),
            .I(N__46240));
    Span4Mux_h I__9836 (
            .O(N__46246),
            .I(N__46237));
    Span4Mux_h I__9835 (
            .O(N__46243),
            .I(N__46234));
    Odrv4 I__9834 (
            .O(N__46240),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_13));
    Odrv4 I__9833 (
            .O(N__46237),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_13));
    Odrv4 I__9832 (
            .O(N__46234),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_13));
    CascadeMux I__9831 (
            .O(N__46227),
            .I(N__46224));
    InMux I__9830 (
            .O(N__46224),
            .I(N__46221));
    LocalMux I__9829 (
            .O(N__46221),
            .I(N__46218));
    Span12Mux_v I__9828 (
            .O(N__46218),
            .I(N__46215));
    Odrv12 I__9827 (
            .O(N__46215),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_31));
    InMux I__9826 (
            .O(N__46212),
            .I(N__46208));
    InMux I__9825 (
            .O(N__46211),
            .I(N__46205));
    LocalMux I__9824 (
            .O(N__46208),
            .I(N__46202));
    LocalMux I__9823 (
            .O(N__46205),
            .I(N__46199));
    Span4Mux_h I__9822 (
            .O(N__46202),
            .I(N__46195));
    Span4Mux_h I__9821 (
            .O(N__46199),
            .I(N__46192));
    InMux I__9820 (
            .O(N__46198),
            .I(N__46189));
    Span4Mux_h I__9819 (
            .O(N__46195),
            .I(N__46186));
    Span4Mux_h I__9818 (
            .O(N__46192),
            .I(N__46183));
    LocalMux I__9817 (
            .O(N__46189),
            .I(N__46180));
    Odrv4 I__9816 (
            .O(N__46186),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_15));
    Odrv4 I__9815 (
            .O(N__46183),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_15));
    Odrv12 I__9814 (
            .O(N__46180),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_15));
    InMux I__9813 (
            .O(N__46173),
            .I(N__46169));
    CascadeMux I__9812 (
            .O(N__46172),
            .I(N__46166));
    LocalMux I__9811 (
            .O(N__46169),
            .I(N__46163));
    InMux I__9810 (
            .O(N__46166),
            .I(N__46160));
    Span4Mux_v I__9809 (
            .O(N__46163),
            .I(N__46154));
    LocalMux I__9808 (
            .O(N__46160),
            .I(N__46154));
    CascadeMux I__9807 (
            .O(N__46159),
            .I(N__46151));
    Span4Mux_v I__9806 (
            .O(N__46154),
            .I(N__46148));
    InMux I__9805 (
            .O(N__46151),
            .I(N__46145));
    Span4Mux_h I__9804 (
            .O(N__46148),
            .I(N__46142));
    LocalMux I__9803 (
            .O(N__46145),
            .I(N__46137));
    Span4Mux_h I__9802 (
            .O(N__46142),
            .I(N__46137));
    Odrv4 I__9801 (
            .O(N__46137),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_13));
    InMux I__9800 (
            .O(N__46134),
            .I(N__46131));
    LocalMux I__9799 (
            .O(N__46131),
            .I(N__46128));
    Span4Mux_h I__9798 (
            .O(N__46128),
            .I(N__46125));
    Span4Mux_h I__9797 (
            .O(N__46125),
            .I(N__46122));
    Span4Mux_h I__9796 (
            .O(N__46122),
            .I(N__46119));
    Odrv4 I__9795 (
            .O(N__46119),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_31));
    InMux I__9794 (
            .O(N__46116),
            .I(N__46112));
    InMux I__9793 (
            .O(N__46115),
            .I(N__46109));
    LocalMux I__9792 (
            .O(N__46112),
            .I(N__46106));
    LocalMux I__9791 (
            .O(N__46109),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11 ));
    Odrv4 I__9790 (
            .O(N__46106),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11 ));
    InMux I__9789 (
            .O(N__46101),
            .I(N__46098));
    LocalMux I__9788 (
            .O(N__46098),
            .I(N__46095));
    Span4Mux_h I__9787 (
            .O(N__46095),
            .I(N__46092));
    Odrv4 I__9786 (
            .O(N__46092),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_11 ));
    CascadeMux I__9785 (
            .O(N__46089),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_21_cascade_ ));
    InMux I__9784 (
            .O(N__46086),
            .I(N__46083));
    LocalMux I__9783 (
            .O(N__46083),
            .I(N__46080));
    Span4Mux_h I__9782 (
            .O(N__46080),
            .I(N__46077));
    Odrv4 I__9781 (
            .O(N__46077),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LHZ0Z5 ));
    InMux I__9780 (
            .O(N__46074),
            .I(N__46071));
    LocalMux I__9779 (
            .O(N__46071),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_21 ));
    CascadeMux I__9778 (
            .O(N__46068),
            .I(N__46065));
    InMux I__9777 (
            .O(N__46065),
            .I(N__46061));
    InMux I__9776 (
            .O(N__46064),
            .I(N__46047));
    LocalMux I__9775 (
            .O(N__46061),
            .I(N__46038));
    InMux I__9774 (
            .O(N__46060),
            .I(N__46035));
    InMux I__9773 (
            .O(N__46059),
            .I(N__46032));
    InMux I__9772 (
            .O(N__46058),
            .I(N__46027));
    InMux I__9771 (
            .O(N__46057),
            .I(N__46027));
    InMux I__9770 (
            .O(N__46056),
            .I(N__46014));
    InMux I__9769 (
            .O(N__46055),
            .I(N__46014));
    InMux I__9768 (
            .O(N__46054),
            .I(N__46014));
    InMux I__9767 (
            .O(N__46053),
            .I(N__46014));
    InMux I__9766 (
            .O(N__46052),
            .I(N__46014));
    InMux I__9765 (
            .O(N__46051),
            .I(N__46014));
    InMux I__9764 (
            .O(N__46050),
            .I(N__46010));
    LocalMux I__9763 (
            .O(N__46047),
            .I(N__46007));
    InMux I__9762 (
            .O(N__46046),
            .I(N__45996));
    InMux I__9761 (
            .O(N__46045),
            .I(N__45996));
    InMux I__9760 (
            .O(N__46044),
            .I(N__45996));
    InMux I__9759 (
            .O(N__46043),
            .I(N__45996));
    InMux I__9758 (
            .O(N__46042),
            .I(N__45996));
    CascadeMux I__9757 (
            .O(N__46041),
            .I(N__45993));
    Span4Mux_h I__9756 (
            .O(N__46038),
            .I(N__45984));
    LocalMux I__9755 (
            .O(N__46035),
            .I(N__45984));
    LocalMux I__9754 (
            .O(N__46032),
            .I(N__45977));
    LocalMux I__9753 (
            .O(N__46027),
            .I(N__45977));
    LocalMux I__9752 (
            .O(N__46014),
            .I(N__45977));
    InMux I__9751 (
            .O(N__46013),
            .I(N__45974));
    LocalMux I__9750 (
            .O(N__46010),
            .I(N__45967));
    Span4Mux_v I__9749 (
            .O(N__46007),
            .I(N__45967));
    LocalMux I__9748 (
            .O(N__45996),
            .I(N__45967));
    InMux I__9747 (
            .O(N__45993),
            .I(N__45962));
    InMux I__9746 (
            .O(N__45992),
            .I(N__45962));
    InMux I__9745 (
            .O(N__45991),
            .I(N__45959));
    InMux I__9744 (
            .O(N__45990),
            .I(N__45954));
    InMux I__9743 (
            .O(N__45989),
            .I(N__45954));
    Span4Mux_h I__9742 (
            .O(N__45984),
            .I(N__45949));
    Span4Mux_v I__9741 (
            .O(N__45977),
            .I(N__45949));
    LocalMux I__9740 (
            .O(N__45974),
            .I(N__45944));
    Span4Mux_h I__9739 (
            .O(N__45967),
            .I(N__45944));
    LocalMux I__9738 (
            .O(N__45962),
            .I(N__45941));
    LocalMux I__9737 (
            .O(N__45959),
            .I(N__45934));
    LocalMux I__9736 (
            .O(N__45954),
            .I(N__45934));
    Span4Mux_h I__9735 (
            .O(N__45949),
            .I(N__45934));
    Span4Mux_h I__9734 (
            .O(N__45944),
            .I(N__45931));
    Span4Mux_v I__9733 (
            .O(N__45941),
            .I(N__45926));
    Span4Mux_h I__9732 (
            .O(N__45934),
            .I(N__45926));
    Odrv4 I__9731 (
            .O(N__45931),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0 ));
    Odrv4 I__9730 (
            .O(N__45926),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0 ));
    CascadeMux I__9729 (
            .O(N__45921),
            .I(N__45916));
    CascadeMux I__9728 (
            .O(N__45920),
            .I(N__45912));
    CascadeMux I__9727 (
            .O(N__45919),
            .I(N__45909));
    InMux I__9726 (
            .O(N__45916),
            .I(N__45899));
    CascadeMux I__9725 (
            .O(N__45915),
            .I(N__45896));
    InMux I__9724 (
            .O(N__45912),
            .I(N__45879));
    InMux I__9723 (
            .O(N__45909),
            .I(N__45879));
    InMux I__9722 (
            .O(N__45908),
            .I(N__45879));
    InMux I__9721 (
            .O(N__45907),
            .I(N__45879));
    InMux I__9720 (
            .O(N__45906),
            .I(N__45879));
    InMux I__9719 (
            .O(N__45905),
            .I(N__45879));
    InMux I__9718 (
            .O(N__45904),
            .I(N__45879));
    InMux I__9717 (
            .O(N__45903),
            .I(N__45879));
    InMux I__9716 (
            .O(N__45902),
            .I(N__45876));
    LocalMux I__9715 (
            .O(N__45899),
            .I(N__45863));
    InMux I__9714 (
            .O(N__45896),
            .I(N__45860));
    LocalMux I__9713 (
            .O(N__45879),
            .I(N__45857));
    LocalMux I__9712 (
            .O(N__45876),
            .I(N__45854));
    InMux I__9711 (
            .O(N__45875),
            .I(N__45843));
    InMux I__9710 (
            .O(N__45874),
            .I(N__45843));
    InMux I__9709 (
            .O(N__45873),
            .I(N__45843));
    InMux I__9708 (
            .O(N__45872),
            .I(N__45843));
    InMux I__9707 (
            .O(N__45871),
            .I(N__45843));
    CascadeMux I__9706 (
            .O(N__45870),
            .I(N__45839));
    InMux I__9705 (
            .O(N__45869),
            .I(N__45836));
    CascadeMux I__9704 (
            .O(N__45868),
            .I(N__45833));
    InMux I__9703 (
            .O(N__45867),
            .I(N__45826));
    InMux I__9702 (
            .O(N__45866),
            .I(N__45826));
    Span4Mux_v I__9701 (
            .O(N__45863),
            .I(N__45819));
    LocalMux I__9700 (
            .O(N__45860),
            .I(N__45819));
    Span4Mux_v I__9699 (
            .O(N__45857),
            .I(N__45819));
    Span4Mux_v I__9698 (
            .O(N__45854),
            .I(N__45814));
    LocalMux I__9697 (
            .O(N__45843),
            .I(N__45814));
    InMux I__9696 (
            .O(N__45842),
            .I(N__45811));
    InMux I__9695 (
            .O(N__45839),
            .I(N__45808));
    LocalMux I__9694 (
            .O(N__45836),
            .I(N__45805));
    InMux I__9693 (
            .O(N__45833),
            .I(N__45798));
    InMux I__9692 (
            .O(N__45832),
            .I(N__45798));
    InMux I__9691 (
            .O(N__45831),
            .I(N__45798));
    LocalMux I__9690 (
            .O(N__45826),
            .I(N__45795));
    Span4Mux_h I__9689 (
            .O(N__45819),
            .I(N__45788));
    Span4Mux_h I__9688 (
            .O(N__45814),
            .I(N__45788));
    LocalMux I__9687 (
            .O(N__45811),
            .I(N__45788));
    LocalMux I__9686 (
            .O(N__45808),
            .I(N__45781));
    Sp12to4 I__9685 (
            .O(N__45805),
            .I(N__45781));
    LocalMux I__9684 (
            .O(N__45798),
            .I(N__45781));
    Span4Mux_v I__9683 (
            .O(N__45795),
            .I(N__45776));
    Span4Mux_h I__9682 (
            .O(N__45788),
            .I(N__45776));
    Span12Mux_h I__9681 (
            .O(N__45781),
            .I(N__45773));
    Odrv4 I__9680 (
            .O(N__45776),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271 ));
    Odrv12 I__9679 (
            .O(N__45773),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271 ));
    CascadeMux I__9678 (
            .O(N__45768),
            .I(N__45765));
    InMux I__9677 (
            .O(N__45765),
            .I(N__45760));
    InMux I__9676 (
            .O(N__45764),
            .I(N__45755));
    InMux I__9675 (
            .O(N__45763),
            .I(N__45755));
    LocalMux I__9674 (
            .O(N__45760),
            .I(N__45752));
    LocalMux I__9673 (
            .O(N__45755),
            .I(N__45749));
    Odrv4 I__9672 (
            .O(N__45752),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_21));
    Odrv4 I__9671 (
            .O(N__45749),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_21));
    InMux I__9670 (
            .O(N__45744),
            .I(N__45739));
    CascadeMux I__9669 (
            .O(N__45743),
            .I(N__45736));
    InMux I__9668 (
            .O(N__45742),
            .I(N__45733));
    LocalMux I__9667 (
            .O(N__45739),
            .I(N__45730));
    InMux I__9666 (
            .O(N__45736),
            .I(N__45727));
    LocalMux I__9665 (
            .O(N__45733),
            .I(N__45724));
    Span4Mux_h I__9664 (
            .O(N__45730),
            .I(N__45719));
    LocalMux I__9663 (
            .O(N__45727),
            .I(N__45719));
    Span4Mux_v I__9662 (
            .O(N__45724),
            .I(N__45714));
    Span4Mux_v I__9661 (
            .O(N__45719),
            .I(N__45714));
    Odrv4 I__9660 (
            .O(N__45714),
            .I(cemf_module_64ch_ctrl_inst1_data_config_21));
    CascadeMux I__9659 (
            .O(N__45711),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_21_cascade_ ));
    InMux I__9658 (
            .O(N__45708),
            .I(N__45705));
    LocalMux I__9657 (
            .O(N__45705),
            .I(N__45702));
    Odrv12 I__9656 (
            .O(N__45702),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDDZ0Z7 ));
    InMux I__9655 (
            .O(N__45699),
            .I(N__45696));
    LocalMux I__9654 (
            .O(N__45696),
            .I(N__45693));
    Span4Mux_v I__9653 (
            .O(N__45693),
            .I(N__45688));
    InMux I__9652 (
            .O(N__45692),
            .I(N__45683));
    InMux I__9651 (
            .O(N__45691),
            .I(N__45683));
    Odrv4 I__9650 (
            .O(N__45688),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_21));
    LocalMux I__9649 (
            .O(N__45683),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_21));
    InMux I__9648 (
            .O(N__45678),
            .I(N__45675));
    LocalMux I__9647 (
            .O(N__45675),
            .I(N__45671));
    CascadeMux I__9646 (
            .O(N__45674),
            .I(N__45667));
    Span4Mux_h I__9645 (
            .O(N__45671),
            .I(N__45664));
    InMux I__9644 (
            .O(N__45670),
            .I(N__45661));
    InMux I__9643 (
            .O(N__45667),
            .I(N__45658));
    Odrv4 I__9642 (
            .O(N__45664),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_21));
    LocalMux I__9641 (
            .O(N__45661),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_21));
    LocalMux I__9640 (
            .O(N__45658),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_21));
    InMux I__9639 (
            .O(N__45651),
            .I(N__45648));
    LocalMux I__9638 (
            .O(N__45648),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_21 ));
    CascadeMux I__9637 (
            .O(N__45645),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_17_cascade_ ));
    CascadeMux I__9636 (
            .O(N__45642),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029DZ0Z7_cascade_ ));
    InMux I__9635 (
            .O(N__45639),
            .I(N__45636));
    LocalMux I__9634 (
            .O(N__45636),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17 ));
    CascadeMux I__9633 (
            .O(N__45633),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17_cascade_ ));
    InMux I__9632 (
            .O(N__45630),
            .I(N__45627));
    LocalMux I__9631 (
            .O(N__45627),
            .I(N__45624));
    Sp12to4 I__9630 (
            .O(N__45624),
            .I(N__45621));
    Odrv12 I__9629 (
            .O(N__45621),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_16 ));
    CascadeMux I__9628 (
            .O(N__45618),
            .I(N__45614));
    InMux I__9627 (
            .O(N__45617),
            .I(N__45610));
    InMux I__9626 (
            .O(N__45614),
            .I(N__45605));
    InMux I__9625 (
            .O(N__45613),
            .I(N__45605));
    LocalMux I__9624 (
            .O(N__45610),
            .I(N__45602));
    LocalMux I__9623 (
            .O(N__45605),
            .I(N__45599));
    Odrv12 I__9622 (
            .O(N__45602),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_17));
    Odrv4 I__9621 (
            .O(N__45599),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_17));
    InMux I__9620 (
            .O(N__45594),
            .I(N__45591));
    LocalMux I__9619 (
            .O(N__45591),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_17 ));
    InMux I__9618 (
            .O(N__45588),
            .I(N__45585));
    LocalMux I__9617 (
            .O(N__45585),
            .I(N__45582));
    Span4Mux_h I__9616 (
            .O(N__45582),
            .I(N__45579));
    Sp12to4 I__9615 (
            .O(N__45579),
            .I(N__45576));
    Odrv12 I__9614 (
            .O(N__45576),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_3Z0Z_26 ));
    CEMux I__9613 (
            .O(N__45573),
            .I(N__45552));
    CEMux I__9612 (
            .O(N__45572),
            .I(N__45552));
    CEMux I__9611 (
            .O(N__45571),
            .I(N__45552));
    CEMux I__9610 (
            .O(N__45570),
            .I(N__45552));
    CEMux I__9609 (
            .O(N__45569),
            .I(N__45552));
    CEMux I__9608 (
            .O(N__45568),
            .I(N__45552));
    CEMux I__9607 (
            .O(N__45567),
            .I(N__45552));
    GlobalMux I__9606 (
            .O(N__45552),
            .I(N__45549));
    gio2CtrlBuf I__9605 (
            .O(N__45549),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g ));
    InMux I__9604 (
            .O(N__45546),
            .I(N__45543));
    LocalMux I__9603 (
            .O(N__45543),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_15 ));
    InMux I__9602 (
            .O(N__45540),
            .I(N__45537));
    LocalMux I__9601 (
            .O(N__45537),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_16 ));
    InMux I__9600 (
            .O(N__45534),
            .I(N__45531));
    LocalMux I__9599 (
            .O(N__45531),
            .I(N__45526));
    InMux I__9598 (
            .O(N__45530),
            .I(N__45523));
    InMux I__9597 (
            .O(N__45529),
            .I(N__45520));
    Odrv12 I__9596 (
            .O(N__45526),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_7));
    LocalMux I__9595 (
            .O(N__45523),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_7));
    LocalMux I__9594 (
            .O(N__45520),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_7));
    InMux I__9593 (
            .O(N__45513),
            .I(N__45510));
    LocalMux I__9592 (
            .O(N__45510),
            .I(N__45507));
    Span12Mux_v I__9591 (
            .O(N__45507),
            .I(N__45504));
    Odrv12 I__9590 (
            .O(N__45504),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_7 ));
    CascadeMux I__9589 (
            .O(N__45501),
            .I(\serializer_mod_inst.un22_next_state_1_cascade_ ));
    InMux I__9588 (
            .O(N__45498),
            .I(N__45495));
    LocalMux I__9587 (
            .O(N__45495),
            .I(N__45492));
    Span4Mux_h I__9586 (
            .O(N__45492),
            .I(N__45489));
    Odrv4 I__9585 (
            .O(N__45489),
            .I(\serializer_mod_inst.un22_next_state ));
    InMux I__9584 (
            .O(N__45486),
            .I(N__45482));
    InMux I__9583 (
            .O(N__45485),
            .I(N__45479));
    LocalMux I__9582 (
            .O(N__45482),
            .I(N__45476));
    LocalMux I__9581 (
            .O(N__45479),
            .I(N__45473));
    Span4Mux_v I__9580 (
            .O(N__45476),
            .I(N__45470));
    Span4Mux_v I__9579 (
            .O(N__45473),
            .I(N__45466));
    Span4Mux_v I__9578 (
            .O(N__45470),
            .I(N__45438));
    InMux I__9577 (
            .O(N__45469),
            .I(N__45435));
    Span4Mux_v I__9576 (
            .O(N__45466),
            .I(N__45432));
    CascadeMux I__9575 (
            .O(N__45465),
            .I(N__45429));
    CascadeMux I__9574 (
            .O(N__45464),
            .I(N__45423));
    CascadeMux I__9573 (
            .O(N__45463),
            .I(N__45419));
    CascadeMux I__9572 (
            .O(N__45462),
            .I(N__45412));
    InMux I__9571 (
            .O(N__45461),
            .I(N__45397));
    InMux I__9570 (
            .O(N__45460),
            .I(N__45397));
    InMux I__9569 (
            .O(N__45459),
            .I(N__45392));
    InMux I__9568 (
            .O(N__45458),
            .I(N__45392));
    InMux I__9567 (
            .O(N__45457),
            .I(N__45385));
    InMux I__9566 (
            .O(N__45456),
            .I(N__45382));
    InMux I__9565 (
            .O(N__45455),
            .I(N__45373));
    InMux I__9564 (
            .O(N__45454),
            .I(N__45373));
    InMux I__9563 (
            .O(N__45453),
            .I(N__45373));
    InMux I__9562 (
            .O(N__45452),
            .I(N__45373));
    InMux I__9561 (
            .O(N__45451),
            .I(N__45364));
    InMux I__9560 (
            .O(N__45450),
            .I(N__45364));
    InMux I__9559 (
            .O(N__45449),
            .I(N__45364));
    InMux I__9558 (
            .O(N__45448),
            .I(N__45364));
    InMux I__9557 (
            .O(N__45447),
            .I(N__45361));
    InMux I__9556 (
            .O(N__45446),
            .I(N__45354));
    InMux I__9555 (
            .O(N__45445),
            .I(N__45349));
    InMux I__9554 (
            .O(N__45444),
            .I(N__45349));
    InMux I__9553 (
            .O(N__45443),
            .I(N__45346));
    InMux I__9552 (
            .O(N__45442),
            .I(N__45341));
    InMux I__9551 (
            .O(N__45441),
            .I(N__45341));
    Span4Mux_h I__9550 (
            .O(N__45438),
            .I(N__45336));
    LocalMux I__9549 (
            .O(N__45435),
            .I(N__45336));
    Span4Mux_v I__9548 (
            .O(N__45432),
            .I(N__45333));
    InMux I__9547 (
            .O(N__45429),
            .I(N__45326));
    InMux I__9546 (
            .O(N__45428),
            .I(N__45326));
    InMux I__9545 (
            .O(N__45427),
            .I(N__45326));
    InMux I__9544 (
            .O(N__45426),
            .I(N__45319));
    InMux I__9543 (
            .O(N__45423),
            .I(N__45319));
    InMux I__9542 (
            .O(N__45422),
            .I(N__45319));
    InMux I__9541 (
            .O(N__45419),
            .I(N__45310));
    InMux I__9540 (
            .O(N__45418),
            .I(N__45310));
    InMux I__9539 (
            .O(N__45417),
            .I(N__45310));
    InMux I__9538 (
            .O(N__45416),
            .I(N__45310));
    InMux I__9537 (
            .O(N__45415),
            .I(N__45303));
    InMux I__9536 (
            .O(N__45412),
            .I(N__45303));
    InMux I__9535 (
            .O(N__45411),
            .I(N__45303));
    InMux I__9534 (
            .O(N__45410),
            .I(N__45294));
    InMux I__9533 (
            .O(N__45409),
            .I(N__45294));
    InMux I__9532 (
            .O(N__45408),
            .I(N__45294));
    InMux I__9531 (
            .O(N__45407),
            .I(N__45294));
    InMux I__9530 (
            .O(N__45406),
            .I(N__45285));
    InMux I__9529 (
            .O(N__45405),
            .I(N__45285));
    InMux I__9528 (
            .O(N__45404),
            .I(N__45285));
    InMux I__9527 (
            .O(N__45403),
            .I(N__45285));
    InMux I__9526 (
            .O(N__45402),
            .I(N__45282));
    LocalMux I__9525 (
            .O(N__45397),
            .I(N__45277));
    LocalMux I__9524 (
            .O(N__45392),
            .I(N__45277));
    InMux I__9523 (
            .O(N__45391),
            .I(N__45274));
    InMux I__9522 (
            .O(N__45390),
            .I(N__45271));
    InMux I__9521 (
            .O(N__45389),
            .I(N__45266));
    InMux I__9520 (
            .O(N__45388),
            .I(N__45266));
    LocalMux I__9519 (
            .O(N__45385),
            .I(N__45263));
    LocalMux I__9518 (
            .O(N__45382),
            .I(N__45254));
    LocalMux I__9517 (
            .O(N__45373),
            .I(N__45254));
    LocalMux I__9516 (
            .O(N__45364),
            .I(N__45254));
    LocalMux I__9515 (
            .O(N__45361),
            .I(N__45254));
    InMux I__9514 (
            .O(N__45360),
            .I(N__45251));
    InMux I__9513 (
            .O(N__45359),
            .I(N__45248));
    CascadeMux I__9512 (
            .O(N__45358),
            .I(N__45236));
    CascadeMux I__9511 (
            .O(N__45357),
            .I(N__45233));
    LocalMux I__9510 (
            .O(N__45354),
            .I(N__45229));
    LocalMux I__9509 (
            .O(N__45349),
            .I(N__45222));
    LocalMux I__9508 (
            .O(N__45346),
            .I(N__45222));
    LocalMux I__9507 (
            .O(N__45341),
            .I(N__45222));
    Span4Mux_h I__9506 (
            .O(N__45336),
            .I(N__45205));
    Span4Mux_h I__9505 (
            .O(N__45333),
            .I(N__45205));
    LocalMux I__9504 (
            .O(N__45326),
            .I(N__45205));
    LocalMux I__9503 (
            .O(N__45319),
            .I(N__45205));
    LocalMux I__9502 (
            .O(N__45310),
            .I(N__45205));
    LocalMux I__9501 (
            .O(N__45303),
            .I(N__45205));
    LocalMux I__9500 (
            .O(N__45294),
            .I(N__45205));
    LocalMux I__9499 (
            .O(N__45285),
            .I(N__45205));
    LocalMux I__9498 (
            .O(N__45282),
            .I(N__45202));
    Span4Mux_v I__9497 (
            .O(N__45277),
            .I(N__45194));
    LocalMux I__9496 (
            .O(N__45274),
            .I(N__45194));
    LocalMux I__9495 (
            .O(N__45271),
            .I(N__45194));
    LocalMux I__9494 (
            .O(N__45266),
            .I(N__45191));
    Span4Mux_v I__9493 (
            .O(N__45263),
            .I(N__45182));
    Span4Mux_v I__9492 (
            .O(N__45254),
            .I(N__45182));
    LocalMux I__9491 (
            .O(N__45251),
            .I(N__45182));
    LocalMux I__9490 (
            .O(N__45248),
            .I(N__45182));
    InMux I__9489 (
            .O(N__45247),
            .I(N__45179));
    InMux I__9488 (
            .O(N__45246),
            .I(N__45169));
    InMux I__9487 (
            .O(N__45245),
            .I(N__45169));
    InMux I__9486 (
            .O(N__45244),
            .I(N__45162));
    InMux I__9485 (
            .O(N__45243),
            .I(N__45162));
    InMux I__9484 (
            .O(N__45242),
            .I(N__45162));
    InMux I__9483 (
            .O(N__45241),
            .I(N__45155));
    InMux I__9482 (
            .O(N__45240),
            .I(N__45155));
    InMux I__9481 (
            .O(N__45239),
            .I(N__45155));
    InMux I__9480 (
            .O(N__45236),
            .I(N__45148));
    InMux I__9479 (
            .O(N__45233),
            .I(N__45148));
    InMux I__9478 (
            .O(N__45232),
            .I(N__45148));
    Span4Mux_v I__9477 (
            .O(N__45229),
            .I(N__45139));
    Span4Mux_v I__9476 (
            .O(N__45222),
            .I(N__45139));
    Span4Mux_v I__9475 (
            .O(N__45205),
            .I(N__45139));
    Span4Mux_v I__9474 (
            .O(N__45202),
            .I(N__45139));
    InMux I__9473 (
            .O(N__45201),
            .I(N__45136));
    Span4Mux_h I__9472 (
            .O(N__45194),
            .I(N__45127));
    Span4Mux_v I__9471 (
            .O(N__45191),
            .I(N__45127));
    Span4Mux_h I__9470 (
            .O(N__45182),
            .I(N__45127));
    LocalMux I__9469 (
            .O(N__45179),
            .I(N__45127));
    InMux I__9468 (
            .O(N__45178),
            .I(N__45120));
    InMux I__9467 (
            .O(N__45177),
            .I(N__45120));
    InMux I__9466 (
            .O(N__45176),
            .I(N__45120));
    InMux I__9465 (
            .O(N__45175),
            .I(N__45117));
    InMux I__9464 (
            .O(N__45174),
            .I(N__45114));
    LocalMux I__9463 (
            .O(N__45169),
            .I(N__45101));
    LocalMux I__9462 (
            .O(N__45162),
            .I(N__45101));
    LocalMux I__9461 (
            .O(N__45155),
            .I(N__45101));
    LocalMux I__9460 (
            .O(N__45148),
            .I(N__45101));
    Sp12to4 I__9459 (
            .O(N__45139),
            .I(N__45101));
    LocalMux I__9458 (
            .O(N__45136),
            .I(N__45101));
    Odrv4 I__9457 (
            .O(N__45127),
            .I(\serializer_mod_inst.current_stateZ0Z_1 ));
    LocalMux I__9456 (
            .O(N__45120),
            .I(\serializer_mod_inst.current_stateZ0Z_1 ));
    LocalMux I__9455 (
            .O(N__45117),
            .I(\serializer_mod_inst.current_stateZ0Z_1 ));
    LocalMux I__9454 (
            .O(N__45114),
            .I(\serializer_mod_inst.current_stateZ0Z_1 ));
    Odrv12 I__9453 (
            .O(N__45101),
            .I(\serializer_mod_inst.current_stateZ0Z_1 ));
    InMux I__9452 (
            .O(N__45090),
            .I(N__45061));
    InMux I__9451 (
            .O(N__45089),
            .I(N__45054));
    InMux I__9450 (
            .O(N__45088),
            .I(N__45036));
    InMux I__9449 (
            .O(N__45087),
            .I(N__45023));
    InMux I__9448 (
            .O(N__45086),
            .I(N__45020));
    InMux I__9447 (
            .O(N__45085),
            .I(N__45013));
    InMux I__9446 (
            .O(N__45084),
            .I(N__45013));
    InMux I__9445 (
            .O(N__45083),
            .I(N__45013));
    InMux I__9444 (
            .O(N__45082),
            .I(N__45010));
    InMux I__9443 (
            .O(N__45081),
            .I(N__44999));
    InMux I__9442 (
            .O(N__45080),
            .I(N__44999));
    InMux I__9441 (
            .O(N__45079),
            .I(N__44999));
    InMux I__9440 (
            .O(N__45078),
            .I(N__44999));
    InMux I__9439 (
            .O(N__45077),
            .I(N__44999));
    InMux I__9438 (
            .O(N__45076),
            .I(N__44992));
    InMux I__9437 (
            .O(N__45075),
            .I(N__44992));
    InMux I__9436 (
            .O(N__45074),
            .I(N__44992));
    InMux I__9435 (
            .O(N__45073),
            .I(N__44983));
    InMux I__9434 (
            .O(N__45072),
            .I(N__44983));
    InMux I__9433 (
            .O(N__45071),
            .I(N__44983));
    InMux I__9432 (
            .O(N__45070),
            .I(N__44983));
    InMux I__9431 (
            .O(N__45069),
            .I(N__44974));
    InMux I__9430 (
            .O(N__45068),
            .I(N__44974));
    InMux I__9429 (
            .O(N__45067),
            .I(N__44974));
    InMux I__9428 (
            .O(N__45066),
            .I(N__44974));
    InMux I__9427 (
            .O(N__45065),
            .I(N__44971));
    InMux I__9426 (
            .O(N__45064),
            .I(N__44968));
    LocalMux I__9425 (
            .O(N__45061),
            .I(N__44965));
    InMux I__9424 (
            .O(N__45060),
            .I(N__44961));
    InMux I__9423 (
            .O(N__45059),
            .I(N__44956));
    InMux I__9422 (
            .O(N__45058),
            .I(N__44956));
    InMux I__9421 (
            .O(N__45057),
            .I(N__44953));
    LocalMux I__9420 (
            .O(N__45054),
            .I(N__44950));
    InMux I__9419 (
            .O(N__45053),
            .I(N__44943));
    InMux I__9418 (
            .O(N__45052),
            .I(N__44943));
    InMux I__9417 (
            .O(N__45051),
            .I(N__44936));
    InMux I__9416 (
            .O(N__45050),
            .I(N__44936));
    InMux I__9415 (
            .O(N__45049),
            .I(N__44936));
    InMux I__9414 (
            .O(N__45048),
            .I(N__44931));
    InMux I__9413 (
            .O(N__45047),
            .I(N__44931));
    InMux I__9412 (
            .O(N__45046),
            .I(N__44926));
    InMux I__9411 (
            .O(N__45045),
            .I(N__44923));
    InMux I__9410 (
            .O(N__45044),
            .I(N__44914));
    InMux I__9409 (
            .O(N__45043),
            .I(N__44914));
    InMux I__9408 (
            .O(N__45042),
            .I(N__44914));
    InMux I__9407 (
            .O(N__45041),
            .I(N__44914));
    InMux I__9406 (
            .O(N__45040),
            .I(N__44909));
    InMux I__9405 (
            .O(N__45039),
            .I(N__44909));
    LocalMux I__9404 (
            .O(N__45036),
            .I(N__44906));
    InMux I__9403 (
            .O(N__45035),
            .I(N__44903));
    InMux I__9402 (
            .O(N__45034),
            .I(N__44889));
    InMux I__9401 (
            .O(N__45033),
            .I(N__44889));
    InMux I__9400 (
            .O(N__45032),
            .I(N__44882));
    InMux I__9399 (
            .O(N__45031),
            .I(N__44882));
    InMux I__9398 (
            .O(N__45030),
            .I(N__44882));
    InMux I__9397 (
            .O(N__45029),
            .I(N__44873));
    InMux I__9396 (
            .O(N__45028),
            .I(N__44873));
    InMux I__9395 (
            .O(N__45027),
            .I(N__44873));
    InMux I__9394 (
            .O(N__45026),
            .I(N__44873));
    LocalMux I__9393 (
            .O(N__45023),
            .I(N__44870));
    LocalMux I__9392 (
            .O(N__45020),
            .I(N__44853));
    LocalMux I__9391 (
            .O(N__45013),
            .I(N__44853));
    LocalMux I__9390 (
            .O(N__45010),
            .I(N__44853));
    LocalMux I__9389 (
            .O(N__44999),
            .I(N__44853));
    LocalMux I__9388 (
            .O(N__44992),
            .I(N__44853));
    LocalMux I__9387 (
            .O(N__44983),
            .I(N__44853));
    LocalMux I__9386 (
            .O(N__44974),
            .I(N__44853));
    LocalMux I__9385 (
            .O(N__44971),
            .I(N__44853));
    LocalMux I__9384 (
            .O(N__44968),
            .I(N__44850));
    Span4Mux_v I__9383 (
            .O(N__44965),
            .I(N__44847));
    InMux I__9382 (
            .O(N__44964),
            .I(N__44844));
    LocalMux I__9381 (
            .O(N__44961),
            .I(N__44835));
    LocalMux I__9380 (
            .O(N__44956),
            .I(N__44835));
    LocalMux I__9379 (
            .O(N__44953),
            .I(N__44835));
    Span4Mux_h I__9378 (
            .O(N__44950),
            .I(N__44835));
    InMux I__9377 (
            .O(N__44949),
            .I(N__44832));
    InMux I__9376 (
            .O(N__44948),
            .I(N__44829));
    LocalMux I__9375 (
            .O(N__44943),
            .I(N__44822));
    LocalMux I__9374 (
            .O(N__44936),
            .I(N__44822));
    LocalMux I__9373 (
            .O(N__44931),
            .I(N__44822));
    InMux I__9372 (
            .O(N__44930),
            .I(N__44817));
    InMux I__9371 (
            .O(N__44929),
            .I(N__44817));
    LocalMux I__9370 (
            .O(N__44926),
            .I(N__44804));
    LocalMux I__9369 (
            .O(N__44923),
            .I(N__44804));
    LocalMux I__9368 (
            .O(N__44914),
            .I(N__44804));
    LocalMux I__9367 (
            .O(N__44909),
            .I(N__44804));
    Span4Mux_v I__9366 (
            .O(N__44906),
            .I(N__44804));
    LocalMux I__9365 (
            .O(N__44903),
            .I(N__44804));
    InMux I__9364 (
            .O(N__44902),
            .I(N__44801));
    InMux I__9363 (
            .O(N__44901),
            .I(N__44796));
    InMux I__9362 (
            .O(N__44900),
            .I(N__44796));
    InMux I__9361 (
            .O(N__44899),
            .I(N__44793));
    InMux I__9360 (
            .O(N__44898),
            .I(N__44788));
    InMux I__9359 (
            .O(N__44897),
            .I(N__44788));
    InMux I__9358 (
            .O(N__44896),
            .I(N__44781));
    InMux I__9357 (
            .O(N__44895),
            .I(N__44781));
    InMux I__9356 (
            .O(N__44894),
            .I(N__44781));
    LocalMux I__9355 (
            .O(N__44889),
            .I(N__44776));
    LocalMux I__9354 (
            .O(N__44882),
            .I(N__44776));
    LocalMux I__9353 (
            .O(N__44873),
            .I(N__44771));
    Span12Mux_h I__9352 (
            .O(N__44870),
            .I(N__44771));
    Span4Mux_v I__9351 (
            .O(N__44853),
            .I(N__44766));
    Span4Mux_v I__9350 (
            .O(N__44850),
            .I(N__44766));
    Span4Mux_v I__9349 (
            .O(N__44847),
            .I(N__44763));
    LocalMux I__9348 (
            .O(N__44844),
            .I(N__44758));
    Span4Mux_v I__9347 (
            .O(N__44835),
            .I(N__44758));
    LocalMux I__9346 (
            .O(N__44832),
            .I(N__44751));
    LocalMux I__9345 (
            .O(N__44829),
            .I(N__44751));
    Span4Mux_v I__9344 (
            .O(N__44822),
            .I(N__44751));
    LocalMux I__9343 (
            .O(N__44817),
            .I(N__44746));
    Span4Mux_v I__9342 (
            .O(N__44804),
            .I(N__44746));
    LocalMux I__9341 (
            .O(N__44801),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    LocalMux I__9340 (
            .O(N__44796),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    LocalMux I__9339 (
            .O(N__44793),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    LocalMux I__9338 (
            .O(N__44788),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    LocalMux I__9337 (
            .O(N__44781),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv4 I__9336 (
            .O(N__44776),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv12 I__9335 (
            .O(N__44771),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv4 I__9334 (
            .O(N__44766),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv4 I__9333 (
            .O(N__44763),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv4 I__9332 (
            .O(N__44758),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv4 I__9331 (
            .O(N__44751),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    Odrv4 I__9330 (
            .O(N__44746),
            .I(\serializer_mod_inst.current_stateZ0Z_0 ));
    CascadeMux I__9329 (
            .O(N__44721),
            .I(N__44718));
    InMux I__9328 (
            .O(N__44718),
            .I(N__44715));
    LocalMux I__9327 (
            .O(N__44715),
            .I(N__44712));
    Span4Mux_h I__9326 (
            .O(N__44712),
            .I(N__44709));
    Odrv4 I__9325 (
            .O(N__44709),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_0 ));
    InMux I__9324 (
            .O(N__44706),
            .I(N__44703));
    LocalMux I__9323 (
            .O(N__44703),
            .I(N__44700));
    Span4Mux_h I__9322 (
            .O(N__44700),
            .I(N__44697));
    Span4Mux_h I__9321 (
            .O(N__44697),
            .I(N__44694));
    Odrv4 I__9320 (
            .O(N__44694),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_0 ));
    InMux I__9319 (
            .O(N__44691),
            .I(N__44688));
    LocalMux I__9318 (
            .O(N__44688),
            .I(N__44685));
    Span12Mux_v I__9317 (
            .O(N__44685),
            .I(N__44682));
    Span12Mux_h I__9316 (
            .O(N__44682),
            .I(N__44679));
    Odrv12 I__9315 (
            .O(N__44679),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_0));
    InMux I__9314 (
            .O(N__44676),
            .I(N__44672));
    InMux I__9313 (
            .O(N__44675),
            .I(N__44669));
    LocalMux I__9312 (
            .O(N__44672),
            .I(N__44666));
    LocalMux I__9311 (
            .O(N__44669),
            .I(N__44654));
    Span4Mux_h I__9310 (
            .O(N__44666),
            .I(N__44651));
    CascadeMux I__9309 (
            .O(N__44665),
            .I(N__44648));
    InMux I__9308 (
            .O(N__44664),
            .I(N__44644));
    InMux I__9307 (
            .O(N__44663),
            .I(N__44641));
    CascadeMux I__9306 (
            .O(N__44662),
            .I(N__44636));
    InMux I__9305 (
            .O(N__44661),
            .I(N__44632));
    CascadeMux I__9304 (
            .O(N__44660),
            .I(N__44629));
    CascadeMux I__9303 (
            .O(N__44659),
            .I(N__44625));
    InMux I__9302 (
            .O(N__44658),
            .I(N__44621));
    InMux I__9301 (
            .O(N__44657),
            .I(N__44618));
    Span4Mux_h I__9300 (
            .O(N__44654),
            .I(N__44609));
    Span4Mux_h I__9299 (
            .O(N__44651),
            .I(N__44609));
    InMux I__9298 (
            .O(N__44648),
            .I(N__44606));
    CascadeMux I__9297 (
            .O(N__44647),
            .I(N__44603));
    LocalMux I__9296 (
            .O(N__44644),
            .I(N__44598));
    LocalMux I__9295 (
            .O(N__44641),
            .I(N__44598));
    InMux I__9294 (
            .O(N__44640),
            .I(N__44593));
    InMux I__9293 (
            .O(N__44639),
            .I(N__44593));
    InMux I__9292 (
            .O(N__44636),
            .I(N__44585));
    InMux I__9291 (
            .O(N__44635),
            .I(N__44585));
    LocalMux I__9290 (
            .O(N__44632),
            .I(N__44582));
    InMux I__9289 (
            .O(N__44629),
            .I(N__44577));
    InMux I__9288 (
            .O(N__44628),
            .I(N__44577));
    InMux I__9287 (
            .O(N__44625),
            .I(N__44572));
    InMux I__9286 (
            .O(N__44624),
            .I(N__44572));
    LocalMux I__9285 (
            .O(N__44621),
            .I(N__44567));
    LocalMux I__9284 (
            .O(N__44618),
            .I(N__44567));
    InMux I__9283 (
            .O(N__44617),
            .I(N__44564));
    InMux I__9282 (
            .O(N__44616),
            .I(N__44557));
    InMux I__9281 (
            .O(N__44615),
            .I(N__44557));
    InMux I__9280 (
            .O(N__44614),
            .I(N__44557));
    Span4Mux_h I__9279 (
            .O(N__44609),
            .I(N__44552));
    LocalMux I__9278 (
            .O(N__44606),
            .I(N__44552));
    InMux I__9277 (
            .O(N__44603),
            .I(N__44549));
    Sp12to4 I__9276 (
            .O(N__44598),
            .I(N__44542));
    LocalMux I__9275 (
            .O(N__44593),
            .I(N__44542));
    CascadeMux I__9274 (
            .O(N__44592),
            .I(N__44538));
    CascadeMux I__9273 (
            .O(N__44591),
            .I(N__44535));
    InMux I__9272 (
            .O(N__44590),
            .I(N__44530));
    LocalMux I__9271 (
            .O(N__44585),
            .I(N__44527));
    Span4Mux_v I__9270 (
            .O(N__44582),
            .I(N__44518));
    LocalMux I__9269 (
            .O(N__44577),
            .I(N__44518));
    LocalMux I__9268 (
            .O(N__44572),
            .I(N__44518));
    Span4Mux_h I__9267 (
            .O(N__44567),
            .I(N__44518));
    LocalMux I__9266 (
            .O(N__44564),
            .I(N__44515));
    LocalMux I__9265 (
            .O(N__44557),
            .I(N__44510));
    Span4Mux_h I__9264 (
            .O(N__44552),
            .I(N__44510));
    LocalMux I__9263 (
            .O(N__44549),
            .I(N__44505));
    InMux I__9262 (
            .O(N__44548),
            .I(N__44500));
    InMux I__9261 (
            .O(N__44547),
            .I(N__44500));
    Span12Mux_s11_v I__9260 (
            .O(N__44542),
            .I(N__44497));
    InMux I__9259 (
            .O(N__44541),
            .I(N__44486));
    InMux I__9258 (
            .O(N__44538),
            .I(N__44486));
    InMux I__9257 (
            .O(N__44535),
            .I(N__44486));
    InMux I__9256 (
            .O(N__44534),
            .I(N__44486));
    InMux I__9255 (
            .O(N__44533),
            .I(N__44486));
    LocalMux I__9254 (
            .O(N__44530),
            .I(N__44479));
    Span4Mux_v I__9253 (
            .O(N__44527),
            .I(N__44479));
    Span4Mux_h I__9252 (
            .O(N__44518),
            .I(N__44479));
    Span4Mux_v I__9251 (
            .O(N__44515),
            .I(N__44474));
    Span4Mux_v I__9250 (
            .O(N__44510),
            .I(N__44474));
    InMux I__9249 (
            .O(N__44509),
            .I(N__44469));
    InMux I__9248 (
            .O(N__44508),
            .I(N__44469));
    Odrv12 I__9247 (
            .O(N__44505),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    LocalMux I__9246 (
            .O(N__44500),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    Odrv12 I__9245 (
            .O(N__44497),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    LocalMux I__9244 (
            .O(N__44486),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    Odrv4 I__9243 (
            .O(N__44479),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    Odrv4 I__9242 (
            .O(N__44474),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    LocalMux I__9241 (
            .O(N__44469),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ));
    CascadeMux I__9240 (
            .O(N__44454),
            .I(N__44451));
    InMux I__9239 (
            .O(N__44451),
            .I(N__44448));
    LocalMux I__9238 (
            .O(N__44448),
            .I(N__44445));
    Span4Mux_h I__9237 (
            .O(N__44445),
            .I(N__44442));
    Sp12to4 I__9236 (
            .O(N__44442),
            .I(N__44439));
    Span12Mux_v I__9235 (
            .O(N__44439),
            .I(N__44436));
    Odrv12 I__9234 (
            .O(N__44436),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_0 ));
    InMux I__9233 (
            .O(N__44433),
            .I(N__44428));
    InMux I__9232 (
            .O(N__44432),
            .I(N__44422));
    InMux I__9231 (
            .O(N__44431),
            .I(N__44422));
    LocalMux I__9230 (
            .O(N__44428),
            .I(N__44419));
    InMux I__9229 (
            .O(N__44427),
            .I(N__44415));
    LocalMux I__9228 (
            .O(N__44422),
            .I(N__44410));
    Span4Mux_h I__9227 (
            .O(N__44419),
            .I(N__44403));
    InMux I__9226 (
            .O(N__44418),
            .I(N__44400));
    LocalMux I__9225 (
            .O(N__44415),
            .I(N__44397));
    InMux I__9224 (
            .O(N__44414),
            .I(N__44394));
    InMux I__9223 (
            .O(N__44413),
            .I(N__44391));
    Span4Mux_h I__9222 (
            .O(N__44410),
            .I(N__44388));
    InMux I__9221 (
            .O(N__44409),
            .I(N__44383));
    InMux I__9220 (
            .O(N__44408),
            .I(N__44383));
    InMux I__9219 (
            .O(N__44407),
            .I(N__44378));
    InMux I__9218 (
            .O(N__44406),
            .I(N__44378));
    Span4Mux_h I__9217 (
            .O(N__44403),
            .I(N__44373));
    LocalMux I__9216 (
            .O(N__44400),
            .I(N__44373));
    Span4Mux_h I__9215 (
            .O(N__44397),
            .I(N__44360));
    LocalMux I__9214 (
            .O(N__44394),
            .I(N__44360));
    LocalMux I__9213 (
            .O(N__44391),
            .I(N__44360));
    Span4Mux_h I__9212 (
            .O(N__44388),
            .I(N__44355));
    LocalMux I__9211 (
            .O(N__44383),
            .I(N__44355));
    LocalMux I__9210 (
            .O(N__44378),
            .I(N__44350));
    Span4Mux_h I__9209 (
            .O(N__44373),
            .I(N__44350));
    InMux I__9208 (
            .O(N__44372),
            .I(N__44343));
    InMux I__9207 (
            .O(N__44371),
            .I(N__44343));
    InMux I__9206 (
            .O(N__44370),
            .I(N__44343));
    InMux I__9205 (
            .O(N__44369),
            .I(N__44340));
    InMux I__9204 (
            .O(N__44368),
            .I(N__44335));
    InMux I__9203 (
            .O(N__44367),
            .I(N__44335));
    Span4Mux_h I__9202 (
            .O(N__44360),
            .I(N__44323));
    Span4Mux_h I__9201 (
            .O(N__44355),
            .I(N__44320));
    Span4Mux_v I__9200 (
            .O(N__44350),
            .I(N__44315));
    LocalMux I__9199 (
            .O(N__44343),
            .I(N__44315));
    LocalMux I__9198 (
            .O(N__44340),
            .I(N__44310));
    LocalMux I__9197 (
            .O(N__44335),
            .I(N__44310));
    InMux I__9196 (
            .O(N__44334),
            .I(N__44305));
    InMux I__9195 (
            .O(N__44333),
            .I(N__44305));
    InMux I__9194 (
            .O(N__44332),
            .I(N__44300));
    InMux I__9193 (
            .O(N__44331),
            .I(N__44300));
    InMux I__9192 (
            .O(N__44330),
            .I(N__44289));
    InMux I__9191 (
            .O(N__44329),
            .I(N__44289));
    InMux I__9190 (
            .O(N__44328),
            .I(N__44289));
    InMux I__9189 (
            .O(N__44327),
            .I(N__44289));
    InMux I__9188 (
            .O(N__44326),
            .I(N__44289));
    Odrv4 I__9187 (
            .O(N__44323),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    Odrv4 I__9186 (
            .O(N__44320),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    Odrv4 I__9185 (
            .O(N__44315),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    Odrv12 I__9184 (
            .O(N__44310),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    LocalMux I__9183 (
            .O(N__44305),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    LocalMux I__9182 (
            .O(N__44300),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    LocalMux I__9181 (
            .O(N__44289),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ));
    InMux I__9180 (
            .O(N__44274),
            .I(N__44271));
    LocalMux I__9179 (
            .O(N__44271),
            .I(N__44268));
    Span4Mux_h I__9178 (
            .O(N__44268),
            .I(N__44265));
    Span4Mux_v I__9177 (
            .O(N__44265),
            .I(N__44262));
    Span4Mux_h I__9176 (
            .O(N__44262),
            .I(N__44259));
    Span4Mux_h I__9175 (
            .O(N__44259),
            .I(N__44256));
    Odrv4 I__9174 (
            .O(N__44256),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_940 ));
    CascadeMux I__9173 (
            .O(N__44253),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_cascade_ ));
    InMux I__9172 (
            .O(N__44250),
            .I(N__44247));
    LocalMux I__9171 (
            .O(N__44247),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_0 ));
    InMux I__9170 (
            .O(N__44244),
            .I(N__44241));
    LocalMux I__9169 (
            .O(N__44241),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_0 ));
    CascadeMux I__9168 (
            .O(N__44238),
            .I(N__44235));
    InMux I__9167 (
            .O(N__44235),
            .I(N__44232));
    LocalMux I__9166 (
            .O(N__44232),
            .I(N__44229));
    Span4Mux_v I__9165 (
            .O(N__44229),
            .I(N__44226));
    Span4Mux_h I__9164 (
            .O(N__44226),
            .I(N__44223));
    Odrv4 I__9163 (
            .O(N__44223),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_25));
    InMux I__9162 (
            .O(N__44220),
            .I(N__44217));
    LocalMux I__9161 (
            .O(N__44217),
            .I(\serializer_mod_inst.shift_regZ0Z_29 ));
    InMux I__9160 (
            .O(N__44214),
            .I(N__44211));
    LocalMux I__9159 (
            .O(N__44211),
            .I(N__44208));
    Odrv12 I__9158 (
            .O(N__44208),
            .I(\serializer_mod_inst.shift_regZ0Z_30 ));
    InMux I__9157 (
            .O(N__44205),
            .I(N__44202));
    LocalMux I__9156 (
            .O(N__44202),
            .I(\serializer_mod_inst.shift_regZ0Z_62 ));
    InMux I__9155 (
            .O(N__44199),
            .I(N__44196));
    LocalMux I__9154 (
            .O(N__44196),
            .I(\serializer_mod_inst.shift_regZ0Z_63 ));
    InMux I__9153 (
            .O(N__44193),
            .I(N__44190));
    LocalMux I__9152 (
            .O(N__44190),
            .I(\serializer_mod_inst.shift_regZ0Z_58 ));
    InMux I__9151 (
            .O(N__44187),
            .I(N__44184));
    LocalMux I__9150 (
            .O(N__44184),
            .I(\serializer_mod_inst.shift_regZ0Z_59 ));
    InMux I__9149 (
            .O(N__44181),
            .I(N__44178));
    LocalMux I__9148 (
            .O(N__44178),
            .I(\serializer_mod_inst.shift_regZ0Z_60 ));
    InMux I__9147 (
            .O(N__44175),
            .I(N__44172));
    LocalMux I__9146 (
            .O(N__44172),
            .I(\serializer_mod_inst.shift_regZ0Z_61 ));
    InMux I__9145 (
            .O(N__44169),
            .I(N__44166));
    LocalMux I__9144 (
            .O(N__44166),
            .I(N__44163));
    Span4Mux_h I__9143 (
            .O(N__44163),
            .I(N__44160));
    Odrv4 I__9142 (
            .O(N__44160),
            .I(\serializer_mod_inst.shift_regZ0Z_56 ));
    InMux I__9141 (
            .O(N__44157),
            .I(N__44154));
    LocalMux I__9140 (
            .O(N__44154),
            .I(\serializer_mod_inst.shift_regZ0Z_57 ));
    CascadeMux I__9139 (
            .O(N__44151),
            .I(N__44148));
    InMux I__9138 (
            .O(N__44148),
            .I(N__44145));
    LocalMux I__9137 (
            .O(N__44145),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_3 ));
    InMux I__9136 (
            .O(N__44142),
            .I(N__44135));
    InMux I__9135 (
            .O(N__44141),
            .I(N__44135));
    InMux I__9134 (
            .O(N__44140),
            .I(N__44132));
    LocalMux I__9133 (
            .O(N__44135),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0 ));
    LocalMux I__9132 (
            .O(N__44132),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0 ));
    CascadeMux I__9131 (
            .O(N__44127),
            .I(N__44124));
    InMux I__9130 (
            .O(N__44124),
            .I(N__44121));
    LocalMux I__9129 (
            .O(N__44121),
            .I(N__44118));
    Sp12to4 I__9128 (
            .O(N__44118),
            .I(N__44115));
    Span12Mux_s8_h I__9127 (
            .O(N__44115),
            .I(N__44112));
    Span12Mux_v I__9126 (
            .O(N__44112),
            .I(N__44109));
    Odrv12 I__9125 (
            .O(N__44109),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_1 ));
    CEMux I__9124 (
            .O(N__44106),
            .I(N__44102));
    CEMux I__9123 (
            .O(N__44105),
            .I(N__44099));
    LocalMux I__9122 (
            .O(N__44102),
            .I(N__44096));
    LocalMux I__9121 (
            .O(N__44099),
            .I(N__44093));
    Span4Mux_h I__9120 (
            .O(N__44096),
            .I(N__44089));
    Span4Mux_v I__9119 (
            .O(N__44093),
            .I(N__44085));
    CEMux I__9118 (
            .O(N__44092),
            .I(N__44082));
    Span4Mux_v I__9117 (
            .O(N__44089),
            .I(N__44079));
    CEMux I__9116 (
            .O(N__44088),
            .I(N__44076));
    Span4Mux_h I__9115 (
            .O(N__44085),
            .I(N__44071));
    LocalMux I__9114 (
            .O(N__44082),
            .I(N__44071));
    Span4Mux_v I__9113 (
            .O(N__44079),
            .I(N__44068));
    LocalMux I__9112 (
            .O(N__44076),
            .I(N__44065));
    Span4Mux_h I__9111 (
            .O(N__44071),
            .I(N__44062));
    Span4Mux_v I__9110 (
            .O(N__44068),
            .I(N__44058));
    Span4Mux_v I__9109 (
            .O(N__44065),
            .I(N__44055));
    Sp12to4 I__9108 (
            .O(N__44062),
            .I(N__44052));
    CEMux I__9107 (
            .O(N__44061),
            .I(N__44049));
    Span4Mux_h I__9106 (
            .O(N__44058),
            .I(N__44046));
    Span4Mux_h I__9105 (
            .O(N__44055),
            .I(N__44043));
    Span12Mux_v I__9104 (
            .O(N__44052),
            .I(N__44040));
    LocalMux I__9103 (
            .O(N__44049),
            .I(N__44035));
    Span4Mux_h I__9102 (
            .O(N__44046),
            .I(N__44035));
    Sp12to4 I__9101 (
            .O(N__44043),
            .I(N__44030));
    Span12Mux_h I__9100 (
            .O(N__44040),
            .I(N__44030));
    Odrv4 I__9099 (
            .O(N__44035),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0 ));
    Odrv12 I__9098 (
            .O(N__44030),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0 ));
    InMux I__9097 (
            .O(N__44025),
            .I(N__44022));
    LocalMux I__9096 (
            .O(N__44022),
            .I(\serializer_mod_inst.shift_regZ0Z_64 ));
    InMux I__9095 (
            .O(N__44019),
            .I(N__44016));
    LocalMux I__9094 (
            .O(N__44016),
            .I(N__44013));
    Span4Mux_h I__9093 (
            .O(N__44013),
            .I(N__44010));
    Odrv4 I__9092 (
            .O(N__44010),
            .I(\serializer_mod_inst.shift_regZ0Z_65 ));
    InMux I__9091 (
            .O(N__44007),
            .I(N__44004));
    LocalMux I__9090 (
            .O(N__44004),
            .I(N__44000));
    InMux I__9089 (
            .O(N__44003),
            .I(N__43997));
    Span4Mux_h I__9088 (
            .O(N__44000),
            .I(N__43994));
    LocalMux I__9087 (
            .O(N__43997),
            .I(N__43991));
    Span4Mux_v I__9086 (
            .O(N__43994),
            .I(N__43988));
    Span4Mux_h I__9085 (
            .O(N__43991),
            .I(N__43985));
    Span4Mux_v I__9084 (
            .O(N__43988),
            .I(N__43982));
    Span4Mux_v I__9083 (
            .O(N__43985),
            .I(N__43979));
    Odrv4 I__9082 (
            .O(N__43982),
            .I(\serializer_mod_inst.shift_regZ0Z_128 ));
    Odrv4 I__9081 (
            .O(N__43979),
            .I(\serializer_mod_inst.shift_regZ0Z_128 ));
    InMux I__9080 (
            .O(N__43974),
            .I(N__43971));
    LocalMux I__9079 (
            .O(N__43971),
            .I(\serializer_mod_inst.shift_regZ0Z_126 ));
    InMux I__9078 (
            .O(N__43968),
            .I(N__43965));
    LocalMux I__9077 (
            .O(N__43965),
            .I(\serializer_mod_inst.shift_regZ0Z_127 ));
    InMux I__9076 (
            .O(N__43962),
            .I(N__43959));
    LocalMux I__9075 (
            .O(N__43959),
            .I(\serializer_mod_inst.shift_regZ0Z_28 ));
    InMux I__9074 (
            .O(N__43956),
            .I(N__43951));
    InMux I__9073 (
            .O(N__43955),
            .I(N__43948));
    InMux I__9072 (
            .O(N__43954),
            .I(N__43945));
    LocalMux I__9071 (
            .O(N__43951),
            .I(N__43942));
    LocalMux I__9070 (
            .O(N__43948),
            .I(N__43939));
    LocalMux I__9069 (
            .O(N__43945),
            .I(N__43933));
    Span4Mux_v I__9068 (
            .O(N__43942),
            .I(N__43933));
    Span4Mux_h I__9067 (
            .O(N__43939),
            .I(N__43928));
    InMux I__9066 (
            .O(N__43938),
            .I(N__43925));
    Sp12to4 I__9065 (
            .O(N__43933),
            .I(N__43922));
    InMux I__9064 (
            .O(N__43932),
            .I(N__43917));
    InMux I__9063 (
            .O(N__43931),
            .I(N__43917));
    Span4Mux_h I__9062 (
            .O(N__43928),
            .I(N__43914));
    LocalMux I__9061 (
            .O(N__43925),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13 ));
    Odrv12 I__9060 (
            .O(N__43922),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13 ));
    LocalMux I__9059 (
            .O(N__43917),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13 ));
    Odrv4 I__9058 (
            .O(N__43914),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13 ));
    InMux I__9057 (
            .O(N__43905),
            .I(N__43898));
    InMux I__9056 (
            .O(N__43904),
            .I(N__43891));
    InMux I__9055 (
            .O(N__43903),
            .I(N__43891));
    InMux I__9054 (
            .O(N__43902),
            .I(N__43891));
    CascadeMux I__9053 (
            .O(N__43901),
            .I(N__43888));
    LocalMux I__9052 (
            .O(N__43898),
            .I(N__43882));
    LocalMux I__9051 (
            .O(N__43891),
            .I(N__43879));
    InMux I__9050 (
            .O(N__43888),
            .I(N__43874));
    InMux I__9049 (
            .O(N__43887),
            .I(N__43874));
    InMux I__9048 (
            .O(N__43886),
            .I(N__43869));
    InMux I__9047 (
            .O(N__43885),
            .I(N__43869));
    Span4Mux_v I__9046 (
            .O(N__43882),
            .I(N__43866));
    Odrv4 I__9045 (
            .O(N__43879),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3 ));
    LocalMux I__9044 (
            .O(N__43874),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3 ));
    LocalMux I__9043 (
            .O(N__43869),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3 ));
    Odrv4 I__9042 (
            .O(N__43866),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3 ));
    InMux I__9041 (
            .O(N__43857),
            .I(N__43854));
    LocalMux I__9040 (
            .O(N__43854),
            .I(N__43849));
    InMux I__9039 (
            .O(N__43853),
            .I(N__43844));
    InMux I__9038 (
            .O(N__43852),
            .I(N__43844));
    Span4Mux_v I__9037 (
            .O(N__43849),
            .I(N__43841));
    LocalMux I__9036 (
            .O(N__43844),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_300_6 ));
    Odrv4 I__9035 (
            .O(N__43841),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_300_6 ));
    InMux I__9034 (
            .O(N__43836),
            .I(N__43833));
    LocalMux I__9033 (
            .O(N__43833),
            .I(N__43830));
    Span4Mux_v I__9032 (
            .O(N__43830),
            .I(N__43825));
    InMux I__9031 (
            .O(N__43829),
            .I(N__43822));
    InMux I__9030 (
            .O(N__43828),
            .I(N__43819));
    Span4Mux_h I__9029 (
            .O(N__43825),
            .I(N__43814));
    LocalMux I__9028 (
            .O(N__43822),
            .I(N__43814));
    LocalMux I__9027 (
            .O(N__43819),
            .I(N__43810));
    Span4Mux_h I__9026 (
            .O(N__43814),
            .I(N__43807));
    InMux I__9025 (
            .O(N__43813),
            .I(N__43804));
    Span4Mux_v I__9024 (
            .O(N__43810),
            .I(N__43799));
    Span4Mux_v I__9023 (
            .O(N__43807),
            .I(N__43799));
    LocalMux I__9022 (
            .O(N__43804),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2 ));
    Odrv4 I__9021 (
            .O(N__43799),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2 ));
    InMux I__9020 (
            .O(N__43794),
            .I(N__43791));
    LocalMux I__9019 (
            .O(N__43791),
            .I(N__43786));
    InMux I__9018 (
            .O(N__43790),
            .I(N__43781));
    InMux I__9017 (
            .O(N__43789),
            .I(N__43781));
    Span4Mux_h I__9016 (
            .O(N__43786),
            .I(N__43778));
    LocalMux I__9015 (
            .O(N__43781),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1425_1 ));
    Odrv4 I__9014 (
            .O(N__43778),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1425_1 ));
    InMux I__9013 (
            .O(N__43773),
            .I(N__43770));
    LocalMux I__9012 (
            .O(N__43770),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_0 ));
    InMux I__9011 (
            .O(N__43767),
            .I(N__43764));
    LocalMux I__9010 (
            .O(N__43764),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_1 ));
    InMux I__9009 (
            .O(N__43761),
            .I(N__43758));
    LocalMux I__9008 (
            .O(N__43758),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_0 ));
    InMux I__9007 (
            .O(N__43755),
            .I(N__43752));
    LocalMux I__9006 (
            .O(N__43752),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_1 ));
    CascadeMux I__9005 (
            .O(N__43749),
            .I(N__43743));
    CascadeMux I__9004 (
            .O(N__43748),
            .I(N__43740));
    InMux I__9003 (
            .O(N__43747),
            .I(N__43734));
    InMux I__9002 (
            .O(N__43746),
            .I(N__43734));
    InMux I__9001 (
            .O(N__43743),
            .I(N__43728));
    InMux I__9000 (
            .O(N__43740),
            .I(N__43728));
    CEMux I__8999 (
            .O(N__43739),
            .I(N__43725));
    LocalMux I__8998 (
            .O(N__43734),
            .I(N__43722));
    CascadeMux I__8997 (
            .O(N__43733),
            .I(N__43717));
    LocalMux I__8996 (
            .O(N__43728),
            .I(N__43712));
    LocalMux I__8995 (
            .O(N__43725),
            .I(N__43712));
    Span4Mux_h I__8994 (
            .O(N__43722),
            .I(N__43709));
    InMux I__8993 (
            .O(N__43721),
            .I(N__43704));
    InMux I__8992 (
            .O(N__43720),
            .I(N__43704));
    InMux I__8991 (
            .O(N__43717),
            .I(N__43701));
    Span4Mux_h I__8990 (
            .O(N__43712),
            .I(N__43698));
    Span4Mux_h I__8989 (
            .O(N__43709),
            .I(N__43695));
    LocalMux I__8988 (
            .O(N__43704),
            .I(\I2C_top_level_inst1.s_load_addr0 ));
    LocalMux I__8987 (
            .O(N__43701),
            .I(\I2C_top_level_inst1.s_load_addr0 ));
    Odrv4 I__8986 (
            .O(N__43698),
            .I(\I2C_top_level_inst1.s_load_addr0 ));
    Odrv4 I__8985 (
            .O(N__43695),
            .I(\I2C_top_level_inst1.s_load_addr0 ));
    CascadeMux I__8984 (
            .O(N__43686),
            .I(N__43683));
    InMux I__8983 (
            .O(N__43683),
            .I(N__43680));
    LocalMux I__8982 (
            .O(N__43680),
            .I(N__43677));
    Span4Mux_h I__8981 (
            .O(N__43677),
            .I(N__43674));
    Odrv4 I__8980 (
            .O(N__43674),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_6_0_0 ));
    InMux I__8979 (
            .O(N__43671),
            .I(N__43666));
    InMux I__8978 (
            .O(N__43670),
            .I(N__43659));
    InMux I__8977 (
            .O(N__43669),
            .I(N__43659));
    LocalMux I__8976 (
            .O(N__43666),
            .I(N__43656));
    InMux I__8975 (
            .O(N__43665),
            .I(N__43651));
    InMux I__8974 (
            .O(N__43664),
            .I(N__43651));
    LocalMux I__8973 (
            .O(N__43659),
            .I(N__43648));
    Span4Mux_h I__8972 (
            .O(N__43656),
            .I(N__43645));
    LocalMux I__8971 (
            .O(N__43651),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0 ));
    Odrv12 I__8970 (
            .O(N__43648),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0 ));
    Odrv4 I__8969 (
            .O(N__43645),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0 ));
    CascadeMux I__8968 (
            .O(N__43638),
            .I(N__43635));
    InMux I__8967 (
            .O(N__43635),
            .I(N__43632));
    LocalMux I__8966 (
            .O(N__43632),
            .I(N__43629));
    Odrv12 I__8965 (
            .O(N__43629),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1378 ));
    CascadeMux I__8964 (
            .O(N__43626),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_1676_cascade_ ));
    InMux I__8963 (
            .O(N__43623),
            .I(N__43620));
    LocalMux I__8962 (
            .O(N__43620),
            .I(N__43616));
    InMux I__8961 (
            .O(N__43619),
            .I(N__43613));
    Span4Mux_h I__8960 (
            .O(N__43616),
            .I(N__43609));
    LocalMux I__8959 (
            .O(N__43613),
            .I(N__43606));
    CascadeMux I__8958 (
            .O(N__43612),
            .I(N__43603));
    Span4Mux_v I__8957 (
            .O(N__43609),
            .I(N__43600));
    Span4Mux_h I__8956 (
            .O(N__43606),
            .I(N__43597));
    InMux I__8955 (
            .O(N__43603),
            .I(N__43594));
    Odrv4 I__8954 (
            .O(N__43600),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21));
    Odrv4 I__8953 (
            .O(N__43597),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21));
    LocalMux I__8952 (
            .O(N__43594),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21));
    CascadeMux I__8951 (
            .O(N__43587),
            .I(c_state_RNIEVJ7_22_cascade_));
    InMux I__8950 (
            .O(N__43584),
            .I(N__43566));
    CascadeMux I__8949 (
            .O(N__43583),
            .I(N__43563));
    CascadeMux I__8948 (
            .O(N__43582),
            .I(N__43556));
    CascadeMux I__8947 (
            .O(N__43581),
            .I(N__43553));
    CascadeMux I__8946 (
            .O(N__43580),
            .I(N__43550));
    CascadeMux I__8945 (
            .O(N__43579),
            .I(N__43546));
    CascadeMux I__8944 (
            .O(N__43578),
            .I(N__43542));
    InMux I__8943 (
            .O(N__43577),
            .I(N__43537));
    CascadeMux I__8942 (
            .O(N__43576),
            .I(N__43534));
    CascadeMux I__8941 (
            .O(N__43575),
            .I(N__43530));
    CascadeMux I__8940 (
            .O(N__43574),
            .I(N__43526));
    CascadeMux I__8939 (
            .O(N__43573),
            .I(N__43523));
    CascadeMux I__8938 (
            .O(N__43572),
            .I(N__43520));
    CascadeMux I__8937 (
            .O(N__43571),
            .I(N__43515));
    InMux I__8936 (
            .O(N__43570),
            .I(N__43508));
    CascadeMux I__8935 (
            .O(N__43569),
            .I(N__43505));
    LocalMux I__8934 (
            .O(N__43566),
            .I(N__43502));
    InMux I__8933 (
            .O(N__43563),
            .I(N__43499));
    CascadeMux I__8932 (
            .O(N__43562),
            .I(N__43496));
    CascadeMux I__8931 (
            .O(N__43561),
            .I(N__43493));
    CascadeMux I__8930 (
            .O(N__43560),
            .I(N__43488));
    CascadeMux I__8929 (
            .O(N__43559),
            .I(N__43484));
    InMux I__8928 (
            .O(N__43556),
            .I(N__43481));
    InMux I__8927 (
            .O(N__43553),
            .I(N__43478));
    InMux I__8926 (
            .O(N__43550),
            .I(N__43463));
    InMux I__8925 (
            .O(N__43549),
            .I(N__43463));
    InMux I__8924 (
            .O(N__43546),
            .I(N__43463));
    InMux I__8923 (
            .O(N__43545),
            .I(N__43463));
    InMux I__8922 (
            .O(N__43542),
            .I(N__43463));
    InMux I__8921 (
            .O(N__43541),
            .I(N__43463));
    InMux I__8920 (
            .O(N__43540),
            .I(N__43463));
    LocalMux I__8919 (
            .O(N__43537),
            .I(N__43460));
    InMux I__8918 (
            .O(N__43534),
            .I(N__43455));
    InMux I__8917 (
            .O(N__43533),
            .I(N__43455));
    InMux I__8916 (
            .O(N__43530),
            .I(N__43452));
    InMux I__8915 (
            .O(N__43529),
            .I(N__43437));
    InMux I__8914 (
            .O(N__43526),
            .I(N__43437));
    InMux I__8913 (
            .O(N__43523),
            .I(N__43437));
    InMux I__8912 (
            .O(N__43520),
            .I(N__43437));
    InMux I__8911 (
            .O(N__43519),
            .I(N__43437));
    InMux I__8910 (
            .O(N__43518),
            .I(N__43437));
    InMux I__8909 (
            .O(N__43515),
            .I(N__43437));
    CascadeMux I__8908 (
            .O(N__43514),
            .I(N__43432));
    InMux I__8907 (
            .O(N__43513),
            .I(N__43428));
    InMux I__8906 (
            .O(N__43512),
            .I(N__43423));
    InMux I__8905 (
            .O(N__43511),
            .I(N__43423));
    LocalMux I__8904 (
            .O(N__43508),
            .I(N__43420));
    InMux I__8903 (
            .O(N__43505),
            .I(N__43417));
    Span4Mux_h I__8902 (
            .O(N__43502),
            .I(N__43412));
    LocalMux I__8901 (
            .O(N__43499),
            .I(N__43412));
    InMux I__8900 (
            .O(N__43496),
            .I(N__43397));
    InMux I__8899 (
            .O(N__43493),
            .I(N__43397));
    InMux I__8898 (
            .O(N__43492),
            .I(N__43397));
    InMux I__8897 (
            .O(N__43491),
            .I(N__43397));
    InMux I__8896 (
            .O(N__43488),
            .I(N__43397));
    InMux I__8895 (
            .O(N__43487),
            .I(N__43397));
    InMux I__8894 (
            .O(N__43484),
            .I(N__43397));
    LocalMux I__8893 (
            .O(N__43481),
            .I(N__43392));
    LocalMux I__8892 (
            .O(N__43478),
            .I(N__43392));
    LocalMux I__8891 (
            .O(N__43463),
            .I(N__43389));
    Span4Mux_h I__8890 (
            .O(N__43460),
            .I(N__43384));
    LocalMux I__8889 (
            .O(N__43455),
            .I(N__43384));
    LocalMux I__8888 (
            .O(N__43452),
            .I(N__43381));
    LocalMux I__8887 (
            .O(N__43437),
            .I(N__43378));
    InMux I__8886 (
            .O(N__43436),
            .I(N__43371));
    InMux I__8885 (
            .O(N__43435),
            .I(N__43371));
    InMux I__8884 (
            .O(N__43432),
            .I(N__43371));
    CascadeMux I__8883 (
            .O(N__43431),
            .I(N__43367));
    LocalMux I__8882 (
            .O(N__43428),
            .I(N__43362));
    LocalMux I__8881 (
            .O(N__43423),
            .I(N__43359));
    Span4Mux_v I__8880 (
            .O(N__43420),
            .I(N__43356));
    LocalMux I__8879 (
            .O(N__43417),
            .I(N__43351));
    Span4Mux_v I__8878 (
            .O(N__43412),
            .I(N__43351));
    LocalMux I__8877 (
            .O(N__43397),
            .I(N__43342));
    Span4Mux_v I__8876 (
            .O(N__43392),
            .I(N__43342));
    Span4Mux_v I__8875 (
            .O(N__43389),
            .I(N__43342));
    Span4Mux_v I__8874 (
            .O(N__43384),
            .I(N__43342));
    Span4Mux_h I__8873 (
            .O(N__43381),
            .I(N__43335));
    Span4Mux_v I__8872 (
            .O(N__43378),
            .I(N__43335));
    LocalMux I__8871 (
            .O(N__43371),
            .I(N__43335));
    InMux I__8870 (
            .O(N__43370),
            .I(N__43330));
    InMux I__8869 (
            .O(N__43367),
            .I(N__43330));
    InMux I__8868 (
            .O(N__43366),
            .I(N__43325));
    InMux I__8867 (
            .O(N__43365),
            .I(N__43325));
    Span12Mux_v I__8866 (
            .O(N__43362),
            .I(N__43322));
    Span4Mux_v I__8865 (
            .O(N__43359),
            .I(N__43315));
    Span4Mux_h I__8864 (
            .O(N__43356),
            .I(N__43315));
    Span4Mux_v I__8863 (
            .O(N__43351),
            .I(N__43315));
    Span4Mux_h I__8862 (
            .O(N__43342),
            .I(N__43310));
    Span4Mux_v I__8861 (
            .O(N__43335),
            .I(N__43310));
    LocalMux I__8860 (
            .O(N__43330),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ));
    LocalMux I__8859 (
            .O(N__43325),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ));
    Odrv12 I__8858 (
            .O(N__43322),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ));
    Odrv4 I__8857 (
            .O(N__43315),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ));
    Odrv4 I__8856 (
            .O(N__43310),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ));
    CascadeMux I__8855 (
            .O(N__43299),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_77_cascade_ ));
    IoInMux I__8854 (
            .O(N__43296),
            .I(N__43293));
    LocalMux I__8853 (
            .O(N__43293),
            .I(N__43290));
    Span4Mux_s1_h I__8852 (
            .O(N__43290),
            .I(N__43287));
    Span4Mux_v I__8851 (
            .O(N__43287),
            .I(N__43284));
    Span4Mux_h I__8850 (
            .O(N__43284),
            .I(N__43281));
    Span4Mux_h I__8849 (
            .O(N__43281),
            .I(N__43278));
    Odrv4 I__8848 (
            .O(N__43278),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0 ));
    InMux I__8847 (
            .O(N__43275),
            .I(N__43272));
    LocalMux I__8846 (
            .O(N__43272),
            .I(N__43269));
    Span4Mux_v I__8845 (
            .O(N__43269),
            .I(N__43265));
    InMux I__8844 (
            .O(N__43268),
            .I(N__43262));
    Odrv4 I__8843 (
            .O(N__43265),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13 ));
    LocalMux I__8842 (
            .O(N__43262),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13 ));
    InMux I__8841 (
            .O(N__43257),
            .I(N__43254));
    LocalMux I__8840 (
            .O(N__43254),
            .I(N__43251));
    Span4Mux_v I__8839 (
            .O(N__43251),
            .I(N__43248));
    Odrv4 I__8838 (
            .O(N__43248),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_13 ));
    InMux I__8837 (
            .O(N__43245),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12 ));
    InMux I__8836 (
            .O(N__43242),
            .I(N__43239));
    LocalMux I__8835 (
            .O(N__43239),
            .I(N__43236));
    Span4Mux_v I__8834 (
            .O(N__43236),
            .I(N__43232));
    InMux I__8833 (
            .O(N__43235),
            .I(N__43229));
    Odrv4 I__8832 (
            .O(N__43232),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14 ));
    LocalMux I__8831 (
            .O(N__43229),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14 ));
    InMux I__8830 (
            .O(N__43224),
            .I(N__43221));
    LocalMux I__8829 (
            .O(N__43221),
            .I(N__43218));
    Span4Mux_h I__8828 (
            .O(N__43218),
            .I(N__43215));
    Odrv4 I__8827 (
            .O(N__43215),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_14 ));
    InMux I__8826 (
            .O(N__43212),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13 ));
    InMux I__8825 (
            .O(N__43209),
            .I(N__43206));
    LocalMux I__8824 (
            .O(N__43206),
            .I(N__43202));
    CascadeMux I__8823 (
            .O(N__43205),
            .I(N__43199));
    Span4Mux_h I__8822 (
            .O(N__43202),
            .I(N__43196));
    InMux I__8821 (
            .O(N__43199),
            .I(N__43193));
    Odrv4 I__8820 (
            .O(N__43196),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15 ));
    LocalMux I__8819 (
            .O(N__43193),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15 ));
    InMux I__8818 (
            .O(N__43188),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_14 ));
    InMux I__8817 (
            .O(N__43185),
            .I(N__43182));
    LocalMux I__8816 (
            .O(N__43182),
            .I(N__43179));
    Span4Mux_h I__8815 (
            .O(N__43179),
            .I(N__43176));
    Odrv4 I__8814 (
            .O(N__43176),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_15 ));
    InMux I__8813 (
            .O(N__43173),
            .I(N__43170));
    LocalMux I__8812 (
            .O(N__43170),
            .I(N__43167));
    Span4Mux_h I__8811 (
            .O(N__43167),
            .I(N__43164));
    Span4Mux_v I__8810 (
            .O(N__43164),
            .I(N__43161));
    Odrv4 I__8809 (
            .O(N__43161),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_103_0 ));
    InMux I__8808 (
            .O(N__43158),
            .I(N__43155));
    LocalMux I__8807 (
            .O(N__43155),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_1 ));
    InMux I__8806 (
            .O(N__43152),
            .I(N__43149));
    LocalMux I__8805 (
            .O(N__43149),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_0 ));
    InMux I__8804 (
            .O(N__43146),
            .I(N__43143));
    LocalMux I__8803 (
            .O(N__43143),
            .I(N__43139));
    CascadeMux I__8802 (
            .O(N__43142),
            .I(N__43136));
    Span4Mux_h I__8801 (
            .O(N__43139),
            .I(N__43131));
    InMux I__8800 (
            .O(N__43136),
            .I(N__43124));
    InMux I__8799 (
            .O(N__43135),
            .I(N__43124));
    InMux I__8798 (
            .O(N__43134),
            .I(N__43124));
    Odrv4 I__8797 (
            .O(N__43131),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5));
    LocalMux I__8796 (
            .O(N__43124),
            .I(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5));
    CascadeMux I__8795 (
            .O(N__43119),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_291_cascade_ ));
    InMux I__8794 (
            .O(N__43116),
            .I(N__43113));
    LocalMux I__8793 (
            .O(N__43113),
            .I(N__43110));
    Span4Mux_h I__8792 (
            .O(N__43110),
            .I(N__43107));
    Odrv4 I__8791 (
            .O(N__43107),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_5 ));
    InMux I__8790 (
            .O(N__43104),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4 ));
    InMux I__8789 (
            .O(N__43101),
            .I(N__43098));
    LocalMux I__8788 (
            .O(N__43098),
            .I(N__43095));
    Span4Mux_h I__8787 (
            .O(N__43095),
            .I(N__43092));
    Odrv4 I__8786 (
            .O(N__43092),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_6 ));
    InMux I__8785 (
            .O(N__43089),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5 ));
    InMux I__8784 (
            .O(N__43086),
            .I(N__43083));
    LocalMux I__8783 (
            .O(N__43083),
            .I(N__43080));
    Span4Mux_h I__8782 (
            .O(N__43080),
            .I(N__43077));
    Odrv4 I__8781 (
            .O(N__43077),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_7 ));
    InMux I__8780 (
            .O(N__43074),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6 ));
    InMux I__8779 (
            .O(N__43071),
            .I(bfn_20_18_0_));
    InMux I__8778 (
            .O(N__43068),
            .I(N__43065));
    LocalMux I__8777 (
            .O(N__43065),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_9 ));
    InMux I__8776 (
            .O(N__43062),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8 ));
    InMux I__8775 (
            .O(N__43059),
            .I(N__43056));
    LocalMux I__8774 (
            .O(N__43056),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_10 ));
    InMux I__8773 (
            .O(N__43053),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9 ));
    InMux I__8772 (
            .O(N__43050),
            .I(N__43047));
    LocalMux I__8771 (
            .O(N__43047),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_11 ));
    InMux I__8770 (
            .O(N__43044),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10 ));
    InMux I__8769 (
            .O(N__43041),
            .I(N__43038));
    LocalMux I__8768 (
            .O(N__43038),
            .I(N__43035));
    Span4Mux_h I__8767 (
            .O(N__43035),
            .I(N__43031));
    InMux I__8766 (
            .O(N__43034),
            .I(N__43028));
    Odrv4 I__8765 (
            .O(N__43031),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12 ));
    LocalMux I__8764 (
            .O(N__43028),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12 ));
    InMux I__8763 (
            .O(N__43023),
            .I(N__43020));
    LocalMux I__8762 (
            .O(N__43020),
            .I(N__43017));
    Span4Mux_v I__8761 (
            .O(N__43017),
            .I(N__43014));
    Span4Mux_h I__8760 (
            .O(N__43014),
            .I(N__43011));
    Odrv4 I__8759 (
            .O(N__43011),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_12 ));
    InMux I__8758 (
            .O(N__43008),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11 ));
    InMux I__8757 (
            .O(N__43005),
            .I(N__43000));
    CascadeMux I__8756 (
            .O(N__43004),
            .I(N__42997));
    CascadeMux I__8755 (
            .O(N__43003),
            .I(N__42994));
    LocalMux I__8754 (
            .O(N__43000),
            .I(N__42991));
    InMux I__8753 (
            .O(N__42997),
            .I(N__42986));
    InMux I__8752 (
            .O(N__42994),
            .I(N__42986));
    Span12Mux_h I__8751 (
            .O(N__42991),
            .I(N__42983));
    LocalMux I__8750 (
            .O(N__42986),
            .I(N__42980));
    Odrv12 I__8749 (
            .O(N__42983),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_2));
    Odrv4 I__8748 (
            .O(N__42980),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_2));
    InMux I__8747 (
            .O(N__42975),
            .I(N__42972));
    LocalMux I__8746 (
            .O(N__42972),
            .I(N__42969));
    Span4Mux_v I__8745 (
            .O(N__42969),
            .I(N__42966));
    Span4Mux_v I__8744 (
            .O(N__42966),
            .I(N__42961));
    InMux I__8743 (
            .O(N__42965),
            .I(N__42956));
    InMux I__8742 (
            .O(N__42964),
            .I(N__42956));
    Odrv4 I__8741 (
            .O(N__42961),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_2));
    LocalMux I__8740 (
            .O(N__42956),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_2));
    InMux I__8739 (
            .O(N__42951),
            .I(N__42948));
    LocalMux I__8738 (
            .O(N__42948),
            .I(N__42945));
    Span4Mux_h I__8737 (
            .O(N__42945),
            .I(N__42941));
    CascadeMux I__8736 (
            .O(N__42944),
            .I(N__42937));
    Span4Mux_v I__8735 (
            .O(N__42941),
            .I(N__42934));
    InMux I__8734 (
            .O(N__42940),
            .I(N__42931));
    InMux I__8733 (
            .O(N__42937),
            .I(N__42928));
    Odrv4 I__8732 (
            .O(N__42934),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_11));
    LocalMux I__8731 (
            .O(N__42931),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_11));
    LocalMux I__8730 (
            .O(N__42928),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_11));
    InMux I__8729 (
            .O(N__42921),
            .I(N__42918));
    LocalMux I__8728 (
            .O(N__42918),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_11 ));
    InMux I__8727 (
            .O(N__42915),
            .I(N__42912));
    LocalMux I__8726 (
            .O(N__42912),
            .I(N__42909));
    Span4Mux_v I__8725 (
            .O(N__42909),
            .I(N__42906));
    Span4Mux_h I__8724 (
            .O(N__42906),
            .I(N__42901));
    InMux I__8723 (
            .O(N__42905),
            .I(N__42898));
    InMux I__8722 (
            .O(N__42904),
            .I(N__42895));
    Odrv4 I__8721 (
            .O(N__42901),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_11));
    LocalMux I__8720 (
            .O(N__42898),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_11));
    LocalMux I__8719 (
            .O(N__42895),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_11));
    InMux I__8718 (
            .O(N__42888),
            .I(N__42885));
    LocalMux I__8717 (
            .O(N__42885),
            .I(N__42882));
    Span4Mux_h I__8716 (
            .O(N__42882),
            .I(N__42879));
    Span4Mux_v I__8715 (
            .O(N__42879),
            .I(N__42876));
    Odrv4 I__8714 (
            .O(N__42876),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_1 ));
    InMux I__8713 (
            .O(N__42873),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0 ));
    InMux I__8712 (
            .O(N__42870),
            .I(N__42867));
    LocalMux I__8711 (
            .O(N__42867),
            .I(N__42864));
    Span4Mux_v I__8710 (
            .O(N__42864),
            .I(N__42861));
    Span4Mux_v I__8709 (
            .O(N__42861),
            .I(N__42858));
    Odrv4 I__8708 (
            .O(N__42858),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_2 ));
    InMux I__8707 (
            .O(N__42855),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1 ));
    InMux I__8706 (
            .O(N__42852),
            .I(N__42849));
    LocalMux I__8705 (
            .O(N__42849),
            .I(N__42846));
    Span4Mux_v I__8704 (
            .O(N__42846),
            .I(N__42843));
    Odrv4 I__8703 (
            .O(N__42843),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_CO ));
    InMux I__8702 (
            .O(N__42840),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2 ));
    InMux I__8701 (
            .O(N__42837),
            .I(N__42834));
    LocalMux I__8700 (
            .O(N__42834),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_4 ));
    InMux I__8699 (
            .O(N__42831),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3 ));
    CascadeMux I__8698 (
            .O(N__42828),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238DZ0Z7_cascade_ ));
    InMux I__8697 (
            .O(N__42825),
            .I(N__42822));
    LocalMux I__8696 (
            .O(N__42822),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_11 ));
    InMux I__8695 (
            .O(N__42819),
            .I(N__42816));
    LocalMux I__8694 (
            .O(N__42816),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_13 ));
    InMux I__8693 (
            .O(N__42813),
            .I(N__42809));
    InMux I__8692 (
            .O(N__42812),
            .I(N__42806));
    LocalMux I__8691 (
            .O(N__42809),
            .I(N__42803));
    LocalMux I__8690 (
            .O(N__42806),
            .I(N__42800));
    Span4Mux_h I__8689 (
            .O(N__42803),
            .I(N__42797));
    Span4Mux_h I__8688 (
            .O(N__42800),
            .I(N__42794));
    Span4Mux_v I__8687 (
            .O(N__42797),
            .I(N__42790));
    Span4Mux_h I__8686 (
            .O(N__42794),
            .I(N__42787));
    InMux I__8685 (
            .O(N__42793),
            .I(N__42784));
    Odrv4 I__8684 (
            .O(N__42790),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_13));
    Odrv4 I__8683 (
            .O(N__42787),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_13));
    LocalMux I__8682 (
            .O(N__42784),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_13));
    InMux I__8681 (
            .O(N__42777),
            .I(N__42774));
    LocalMux I__8680 (
            .O(N__42774),
            .I(N__42771));
    Span4Mux_h I__8679 (
            .O(N__42771),
            .I(N__42768));
    Odrv4 I__8678 (
            .O(N__42768),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_23 ));
    InMux I__8677 (
            .O(N__42765),
            .I(N__42762));
    LocalMux I__8676 (
            .O(N__42762),
            .I(N__42759));
    Span4Mux_h I__8675 (
            .O(N__42759),
            .I(N__42755));
    CascadeMux I__8674 (
            .O(N__42758),
            .I(N__42752));
    Span4Mux_v I__8673 (
            .O(N__42755),
            .I(N__42748));
    InMux I__8672 (
            .O(N__42752),
            .I(N__42743));
    InMux I__8671 (
            .O(N__42751),
            .I(N__42743));
    Odrv4 I__8670 (
            .O(N__42748),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_10));
    LocalMux I__8669 (
            .O(N__42743),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_10));
    InMux I__8668 (
            .O(N__42738),
            .I(N__42735));
    LocalMux I__8667 (
            .O(N__42735),
            .I(N__42732));
    Span4Mux_v I__8666 (
            .O(N__42732),
            .I(N__42729));
    Span4Mux_h I__8665 (
            .O(N__42729),
            .I(N__42725));
    CascadeMux I__8664 (
            .O(N__42728),
            .I(N__42721));
    Span4Mux_v I__8663 (
            .O(N__42725),
            .I(N__42718));
    InMux I__8662 (
            .O(N__42724),
            .I(N__42715));
    InMux I__8661 (
            .O(N__42721),
            .I(N__42712));
    Odrv4 I__8660 (
            .O(N__42718),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_10));
    LocalMux I__8659 (
            .O(N__42715),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_10));
    LocalMux I__8658 (
            .O(N__42712),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_10));
    InMux I__8657 (
            .O(N__42705),
            .I(N__42702));
    LocalMux I__8656 (
            .O(N__42702),
            .I(N__42698));
    CascadeMux I__8655 (
            .O(N__42701),
            .I(N__42694));
    Span4Mux_h I__8654 (
            .O(N__42698),
            .I(N__42691));
    InMux I__8653 (
            .O(N__42697),
            .I(N__42686));
    InMux I__8652 (
            .O(N__42694),
            .I(N__42686));
    Odrv4 I__8651 (
            .O(N__42691),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_12));
    LocalMux I__8650 (
            .O(N__42686),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_12));
    InMux I__8649 (
            .O(N__42681),
            .I(N__42678));
    LocalMux I__8648 (
            .O(N__42678),
            .I(N__42675));
    Span4Mux_v I__8647 (
            .O(N__42675),
            .I(N__42671));
    CascadeMux I__8646 (
            .O(N__42674),
            .I(N__42667));
    Span4Mux_v I__8645 (
            .O(N__42671),
            .I(N__42664));
    InMux I__8644 (
            .O(N__42670),
            .I(N__42661));
    InMux I__8643 (
            .O(N__42667),
            .I(N__42658));
    Span4Mux_h I__8642 (
            .O(N__42664),
            .I(N__42655));
    LocalMux I__8641 (
            .O(N__42661),
            .I(N__42650));
    LocalMux I__8640 (
            .O(N__42658),
            .I(N__42650));
    Odrv4 I__8639 (
            .O(N__42655),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_22));
    Odrv4 I__8638 (
            .O(N__42650),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_22));
    CascadeMux I__8637 (
            .O(N__42645),
            .I(N__42640));
    CascadeMux I__8636 (
            .O(N__42644),
            .I(N__42637));
    InMux I__8635 (
            .O(N__42643),
            .I(N__42634));
    InMux I__8634 (
            .O(N__42640),
            .I(N__42629));
    InMux I__8633 (
            .O(N__42637),
            .I(N__42629));
    LocalMux I__8632 (
            .O(N__42634),
            .I(N__42626));
    LocalMux I__8631 (
            .O(N__42629),
            .I(N__42623));
    Span4Mux_h I__8630 (
            .O(N__42626),
            .I(N__42620));
    Span4Mux_h I__8629 (
            .O(N__42623),
            .I(N__42617));
    Odrv4 I__8628 (
            .O(N__42620),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_14));
    Odrv4 I__8627 (
            .O(N__42617),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_14));
    InMux I__8626 (
            .O(N__42612),
            .I(N__42609));
    LocalMux I__8625 (
            .O(N__42609),
            .I(N__42605));
    CascadeMux I__8624 (
            .O(N__42608),
            .I(N__42601));
    Span4Mux_h I__8623 (
            .O(N__42605),
            .I(N__42598));
    InMux I__8622 (
            .O(N__42604),
            .I(N__42593));
    InMux I__8621 (
            .O(N__42601),
            .I(N__42593));
    Span4Mux_v I__8620 (
            .O(N__42598),
            .I(N__42590));
    LocalMux I__8619 (
            .O(N__42593),
            .I(N__42587));
    Odrv4 I__8618 (
            .O(N__42590),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_15));
    Odrv4 I__8617 (
            .O(N__42587),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_15));
    InMux I__8616 (
            .O(N__42582),
            .I(N__42579));
    LocalMux I__8615 (
            .O(N__42579),
            .I(N__42574));
    InMux I__8614 (
            .O(N__42578),
            .I(N__42569));
    InMux I__8613 (
            .O(N__42577),
            .I(N__42569));
    Span12Mux_v I__8612 (
            .O(N__42574),
            .I(N__42566));
    LocalMux I__8611 (
            .O(N__42569),
            .I(N__42563));
    Odrv12 I__8610 (
            .O(N__42566),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_16));
    Odrv4 I__8609 (
            .O(N__42563),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_16));
    InMux I__8608 (
            .O(N__42558),
            .I(N__42555));
    LocalMux I__8607 (
            .O(N__42555),
            .I(N__42551));
    InMux I__8606 (
            .O(N__42554),
            .I(N__42547));
    Span4Mux_v I__8605 (
            .O(N__42551),
            .I(N__42544));
    InMux I__8604 (
            .O(N__42550),
            .I(N__42541));
    LocalMux I__8603 (
            .O(N__42547),
            .I(N__42538));
    Span4Mux_h I__8602 (
            .O(N__42544),
            .I(N__42531));
    LocalMux I__8601 (
            .O(N__42541),
            .I(N__42531));
    Span4Mux_v I__8600 (
            .O(N__42538),
            .I(N__42531));
    Odrv4 I__8599 (
            .O(N__42531),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_11));
    CascadeMux I__8598 (
            .O(N__42528),
            .I(N__42524));
    InMux I__8597 (
            .O(N__42527),
            .I(N__42521));
    InMux I__8596 (
            .O(N__42524),
            .I(N__42518));
    LocalMux I__8595 (
            .O(N__42521),
            .I(N__42515));
    LocalMux I__8594 (
            .O(N__42518),
            .I(N__42511));
    Span4Mux_h I__8593 (
            .O(N__42515),
            .I(N__42508));
    InMux I__8592 (
            .O(N__42514),
            .I(N__42505));
    Span4Mux_v I__8591 (
            .O(N__42511),
            .I(N__42502));
    Span4Mux_v I__8590 (
            .O(N__42508),
            .I(N__42497));
    LocalMux I__8589 (
            .O(N__42505),
            .I(N__42497));
    Span4Mux_h I__8588 (
            .O(N__42502),
            .I(N__42494));
    Odrv4 I__8587 (
            .O(N__42497),
            .I(cemf_module_64ch_ctrl_inst1_data_config_11));
    Odrv4 I__8586 (
            .O(N__42494),
            .I(cemf_module_64ch_ctrl_inst1_data_config_11));
    CascadeMux I__8585 (
            .O(N__42489),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_11_cascade_ ));
    InMux I__8584 (
            .O(N__42486),
            .I(N__42483));
    LocalMux I__8583 (
            .O(N__42483),
            .I(N__42478));
    InMux I__8582 (
            .O(N__42482),
            .I(N__42475));
    CascadeMux I__8581 (
            .O(N__42481),
            .I(N__42472));
    Span4Mux_v I__8580 (
            .O(N__42478),
            .I(N__42467));
    LocalMux I__8579 (
            .O(N__42475),
            .I(N__42467));
    InMux I__8578 (
            .O(N__42472),
            .I(N__42464));
    Span4Mux_h I__8577 (
            .O(N__42467),
            .I(N__42461));
    LocalMux I__8576 (
            .O(N__42464),
            .I(N__42458));
    Span4Mux_h I__8575 (
            .O(N__42461),
            .I(N__42455));
    Span12Mux_v I__8574 (
            .O(N__42458),
            .I(N__42452));
    Odrv4 I__8573 (
            .O(N__42455),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_4));
    Odrv12 I__8572 (
            .O(N__42452),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_4));
    InMux I__8571 (
            .O(N__42447),
            .I(N__42440));
    InMux I__8570 (
            .O(N__42446),
            .I(N__42440));
    CascadeMux I__8569 (
            .O(N__42445),
            .I(N__42437));
    LocalMux I__8568 (
            .O(N__42440),
            .I(N__42434));
    InMux I__8567 (
            .O(N__42437),
            .I(N__42431));
    Span4Mux_h I__8566 (
            .O(N__42434),
            .I(N__42428));
    LocalMux I__8565 (
            .O(N__42431),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_20));
    Odrv4 I__8564 (
            .O(N__42428),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_20));
    InMux I__8563 (
            .O(N__42423),
            .I(N__42420));
    LocalMux I__8562 (
            .O(N__42420),
            .I(N__42416));
    CascadeMux I__8561 (
            .O(N__42419),
            .I(N__42413));
    Span4Mux_v I__8560 (
            .O(N__42416),
            .I(N__42409));
    InMux I__8559 (
            .O(N__42413),
            .I(N__42404));
    InMux I__8558 (
            .O(N__42412),
            .I(N__42404));
    Sp12to4 I__8557 (
            .O(N__42409),
            .I(N__42399));
    LocalMux I__8556 (
            .O(N__42404),
            .I(N__42399));
    Odrv12 I__8555 (
            .O(N__42399),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_20));
    InMux I__8554 (
            .O(N__42396),
            .I(N__42393));
    LocalMux I__8553 (
            .O(N__42393),
            .I(N__42390));
    Odrv12 I__8552 (
            .O(N__42390),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_15 ));
    CascadeMux I__8551 (
            .O(N__42387),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_15_cascade_ ));
    CascadeMux I__8550 (
            .O(N__42384),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8DZ0Z7_cascade_ ));
    InMux I__8549 (
            .O(N__42381),
            .I(N__42378));
    LocalMux I__8548 (
            .O(N__42378),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15 ));
    InMux I__8547 (
            .O(N__42375),
            .I(N__42372));
    LocalMux I__8546 (
            .O(N__42372),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_14 ));
    CascadeMux I__8545 (
            .O(N__42369),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15_cascade_ ));
    CascadeMux I__8544 (
            .O(N__42366),
            .I(N__42363));
    InMux I__8543 (
            .O(N__42363),
            .I(N__42360));
    LocalMux I__8542 (
            .O(N__42360),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_16 ));
    CascadeMux I__8541 (
            .O(N__42357),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8DZ0Z7_cascade_ ));
    InMux I__8540 (
            .O(N__42354),
            .I(N__42351));
    LocalMux I__8539 (
            .O(N__42351),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16 ));
    CascadeMux I__8538 (
            .O(N__42348),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16_cascade_ ));
    InMux I__8537 (
            .O(N__42345),
            .I(N__42342));
    LocalMux I__8536 (
            .O(N__42342),
            .I(N__42339));
    Odrv4 I__8535 (
            .O(N__42339),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_15 ));
    InMux I__8534 (
            .O(N__42336),
            .I(N__42333));
    LocalMux I__8533 (
            .O(N__42333),
            .I(N__42330));
    Odrv12 I__8532 (
            .O(N__42330),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_16 ));
    InMux I__8531 (
            .O(N__42327),
            .I(N__42324));
    LocalMux I__8530 (
            .O(N__42324),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_16 ));
    CascadeMux I__8529 (
            .O(N__42321),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_16_cascade_ ));
    InMux I__8528 (
            .O(N__42318),
            .I(N__42315));
    LocalMux I__8527 (
            .O(N__42315),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_16 ));
    InMux I__8526 (
            .O(N__42312),
            .I(N__42309));
    LocalMux I__8525 (
            .O(N__42309),
            .I(N__42306));
    Span4Mux_h I__8524 (
            .O(N__42306),
            .I(N__42303));
    Span4Mux_h I__8523 (
            .O(N__42303),
            .I(N__42300));
    Span4Mux_v I__8522 (
            .O(N__42300),
            .I(N__42297));
    Span4Mux_h I__8521 (
            .O(N__42297),
            .I(N__42294));
    Odrv4 I__8520 (
            .O(N__42294),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_24));
    InMux I__8519 (
            .O(N__42291),
            .I(N__42288));
    LocalMux I__8518 (
            .O(N__42288),
            .I(N__42285));
    Span4Mux_h I__8517 (
            .O(N__42285),
            .I(N__42282));
    Odrv4 I__8516 (
            .O(N__42282),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_24 ));
    InMux I__8515 (
            .O(N__42279),
            .I(N__42274));
    InMux I__8514 (
            .O(N__42278),
            .I(N__42269));
    InMux I__8513 (
            .O(N__42277),
            .I(N__42269));
    LocalMux I__8512 (
            .O(N__42274),
            .I(N__42266));
    LocalMux I__8511 (
            .O(N__42269),
            .I(N__42263));
    Span12Mux_h I__8510 (
            .O(N__42266),
            .I(N__42260));
    Span4Mux_v I__8509 (
            .O(N__42263),
            .I(N__42257));
    Odrv12 I__8508 (
            .O(N__42260),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_22));
    Odrv4 I__8507 (
            .O(N__42257),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_22));
    InMux I__8506 (
            .O(N__42252),
            .I(N__42249));
    LocalMux I__8505 (
            .O(N__42249),
            .I(N__42244));
    InMux I__8504 (
            .O(N__42248),
            .I(N__42239));
    InMux I__8503 (
            .O(N__42247),
            .I(N__42239));
    Span4Mux_h I__8502 (
            .O(N__42244),
            .I(N__42236));
    LocalMux I__8501 (
            .O(N__42239),
            .I(N__42233));
    Span4Mux_h I__8500 (
            .O(N__42236),
            .I(N__42230));
    Span4Mux_h I__8499 (
            .O(N__42233),
            .I(N__42227));
    Span4Mux_h I__8498 (
            .O(N__42230),
            .I(N__42224));
    Span4Mux_h I__8497 (
            .O(N__42227),
            .I(N__42221));
    Odrv4 I__8496 (
            .O(N__42224),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_4));
    Odrv4 I__8495 (
            .O(N__42221),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_4));
    InMux I__8494 (
            .O(N__42216),
            .I(N__42213));
    LocalMux I__8493 (
            .O(N__42213),
            .I(N__42209));
    InMux I__8492 (
            .O(N__42212),
            .I(N__42205));
    Span4Mux_h I__8491 (
            .O(N__42209),
            .I(N__42202));
    InMux I__8490 (
            .O(N__42208),
            .I(N__42199));
    LocalMux I__8489 (
            .O(N__42205),
            .I(N__42196));
    Sp12to4 I__8488 (
            .O(N__42202),
            .I(N__42191));
    LocalMux I__8487 (
            .O(N__42199),
            .I(N__42191));
    Span4Mux_h I__8486 (
            .O(N__42196),
            .I(N__42188));
    Span12Mux_v I__8485 (
            .O(N__42191),
            .I(N__42185));
    Span4Mux_h I__8484 (
            .O(N__42188),
            .I(N__42182));
    Odrv12 I__8483 (
            .O(N__42185),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_5));
    Odrv4 I__8482 (
            .O(N__42182),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_5));
    InMux I__8481 (
            .O(N__42177),
            .I(N__42172));
    CascadeMux I__8480 (
            .O(N__42176),
            .I(N__42169));
    InMux I__8479 (
            .O(N__42175),
            .I(N__42166));
    LocalMux I__8478 (
            .O(N__42172),
            .I(N__42163));
    InMux I__8477 (
            .O(N__42169),
            .I(N__42160));
    LocalMux I__8476 (
            .O(N__42166),
            .I(N__42153));
    Span4Mux_v I__8475 (
            .O(N__42163),
            .I(N__42153));
    LocalMux I__8474 (
            .O(N__42160),
            .I(N__42153));
    Span4Mux_h I__8473 (
            .O(N__42153),
            .I(N__42150));
    Span4Mux_h I__8472 (
            .O(N__42150),
            .I(N__42147));
    Odrv4 I__8471 (
            .O(N__42147),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_6));
    InMux I__8470 (
            .O(N__42144),
            .I(N__42141));
    LocalMux I__8469 (
            .O(N__42141),
            .I(N__42138));
    Span4Mux_v I__8468 (
            .O(N__42138),
            .I(N__42135));
    Span4Mux_v I__8467 (
            .O(N__42135),
            .I(N__42132));
    Sp12to4 I__8466 (
            .O(N__42132),
            .I(N__42129));
    Odrv12 I__8465 (
            .O(N__42129),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_27));
    CascadeMux I__8464 (
            .O(N__42126),
            .I(N__42123));
    InMux I__8463 (
            .O(N__42123),
            .I(N__42120));
    LocalMux I__8462 (
            .O(N__42120),
            .I(N__42117));
    Span4Mux_v I__8461 (
            .O(N__42117),
            .I(N__42114));
    Sp12to4 I__8460 (
            .O(N__42114),
            .I(N__42111));
    Span12Mux_h I__8459 (
            .O(N__42111),
            .I(N__42108));
    Odrv12 I__8458 (
            .O(N__42108),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_27));
    CascadeMux I__8457 (
            .O(N__42105),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_27_cascade_ ));
    InMux I__8456 (
            .O(N__42102),
            .I(N__42099));
    LocalMux I__8455 (
            .O(N__42099),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_27 ));
    InMux I__8454 (
            .O(N__42096),
            .I(N__42093));
    LocalMux I__8453 (
            .O(N__42093),
            .I(N__42090));
    Span4Mux_h I__8452 (
            .O(N__42090),
            .I(N__42087));
    Odrv4 I__8451 (
            .O(N__42087),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_27 ));
    CascadeMux I__8450 (
            .O(N__42084),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_27_cascade_ ));
    InMux I__8449 (
            .O(N__42081),
            .I(N__42078));
    LocalMux I__8448 (
            .O(N__42078),
            .I(N__42075));
    Odrv12 I__8447 (
            .O(N__42075),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_654 ));
    InMux I__8446 (
            .O(N__42072),
            .I(N__42069));
    LocalMux I__8445 (
            .O(N__42069),
            .I(N__42066));
    Span12Mux_h I__8444 (
            .O(N__42066),
            .I(N__42063));
    Odrv12 I__8443 (
            .O(N__42063),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_27 ));
    InMux I__8442 (
            .O(N__42060),
            .I(N__42057));
    LocalMux I__8441 (
            .O(N__42057),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_27 ));
    InMux I__8440 (
            .O(N__42054),
            .I(N__42051));
    LocalMux I__8439 (
            .O(N__42051),
            .I(N__42048));
    Span4Mux_v I__8438 (
            .O(N__42048),
            .I(N__42045));
    Sp12to4 I__8437 (
            .O(N__42045),
            .I(N__42042));
    Span12Mux_h I__8436 (
            .O(N__42042),
            .I(N__42039));
    Odrv12 I__8435 (
            .O(N__42039),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_16));
    CascadeMux I__8434 (
            .O(N__42036),
            .I(N__42033));
    InMux I__8433 (
            .O(N__42033),
            .I(N__42030));
    LocalMux I__8432 (
            .O(N__42030),
            .I(N__42027));
    Span4Mux_v I__8431 (
            .O(N__42027),
            .I(N__42024));
    Span4Mux_h I__8430 (
            .O(N__42024),
            .I(N__42021));
    Sp12to4 I__8429 (
            .O(N__42021),
            .I(N__42018));
    Odrv12 I__8428 (
            .O(N__42018),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_16));
    CascadeMux I__8427 (
            .O(N__42015),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_16_cascade_ ));
    InMux I__8426 (
            .O(N__42012),
            .I(N__42007));
    CascadeMux I__8425 (
            .O(N__42011),
            .I(N__42004));
    CascadeMux I__8424 (
            .O(N__42010),
            .I(N__42001));
    LocalMux I__8423 (
            .O(N__42007),
            .I(N__41998));
    InMux I__8422 (
            .O(N__42004),
            .I(N__41993));
    InMux I__8421 (
            .O(N__42001),
            .I(N__41993));
    Odrv4 I__8420 (
            .O(N__41998),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_16));
    LocalMux I__8419 (
            .O(N__41993),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_16));
    InMux I__8418 (
            .O(N__41988),
            .I(N__41985));
    LocalMux I__8417 (
            .O(N__41985),
            .I(N__41982));
    Span12Mux_s10_v I__8416 (
            .O(N__41982),
            .I(N__41979));
    Span12Mux_v I__8415 (
            .O(N__41979),
            .I(N__41976));
    Span12Mux_h I__8414 (
            .O(N__41976),
            .I(N__41973));
    Odrv12 I__8413 (
            .O(N__41973),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_16));
    InMux I__8412 (
            .O(N__41970),
            .I(N__41967));
    LocalMux I__8411 (
            .O(N__41967),
            .I(N__41964));
    Span4Mux_h I__8410 (
            .O(N__41964),
            .I(N__41961));
    Span4Mux_v I__8409 (
            .O(N__41961),
            .I(N__41958));
    Span4Mux_h I__8408 (
            .O(N__41958),
            .I(N__41955));
    Odrv4 I__8407 (
            .O(N__41955),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_764 ));
    CascadeMux I__8406 (
            .O(N__41952),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_16_cascade_ ));
    InMux I__8405 (
            .O(N__41949),
            .I(N__41946));
    LocalMux I__8404 (
            .O(N__41946),
            .I(\serializer_mod_inst.shift_regZ0Z_27 ));
    InMux I__8403 (
            .O(N__41943),
            .I(N__41940));
    LocalMux I__8402 (
            .O(N__41940),
            .I(\serializer_mod_inst.shift_regZ0Z_22 ));
    InMux I__8401 (
            .O(N__41937),
            .I(N__41934));
    LocalMux I__8400 (
            .O(N__41934),
            .I(\serializer_mod_inst.shift_regZ0Z_23 ));
    InMux I__8399 (
            .O(N__41931),
            .I(N__41928));
    LocalMux I__8398 (
            .O(N__41928),
            .I(N__41925));
    Odrv4 I__8397 (
            .O(N__41925),
            .I(\serializer_mod_inst.shift_regZ0Z_108 ));
    InMux I__8396 (
            .O(N__41922),
            .I(N__41919));
    LocalMux I__8395 (
            .O(N__41919),
            .I(N__41916));
    Odrv12 I__8394 (
            .O(N__41916),
            .I(\serializer_mod_inst.shift_regZ0Z_109 ));
    InMux I__8393 (
            .O(N__41913),
            .I(N__41910));
    LocalMux I__8392 (
            .O(N__41910),
            .I(N__41907));
    Odrv4 I__8391 (
            .O(N__41907),
            .I(\serializer_mod_inst.shift_regZ0Z_19 ));
    InMux I__8390 (
            .O(N__41904),
            .I(N__41901));
    LocalMux I__8389 (
            .O(N__41901),
            .I(\serializer_mod_inst.shift_regZ0Z_20 ));
    InMux I__8388 (
            .O(N__41898),
            .I(N__41895));
    LocalMux I__8387 (
            .O(N__41895),
            .I(\serializer_mod_inst.shift_regZ0Z_24 ));
    InMux I__8386 (
            .O(N__41892),
            .I(N__41889));
    LocalMux I__8385 (
            .O(N__41889),
            .I(\serializer_mod_inst.shift_regZ0Z_124 ));
    InMux I__8384 (
            .O(N__41886),
            .I(N__41883));
    LocalMux I__8383 (
            .O(N__41883),
            .I(N__41880));
    Odrv4 I__8382 (
            .O(N__41880),
            .I(\serializer_mod_inst.shift_regZ0Z_125 ));
    InMux I__8381 (
            .O(N__41877),
            .I(N__41874));
    LocalMux I__8380 (
            .O(N__41874),
            .I(N__41871));
    Span4Mux_v I__8379 (
            .O(N__41871),
            .I(N__41868));
    Odrv4 I__8378 (
            .O(N__41868),
            .I(\serializer_mod_inst.shift_regZ0Z_122 ));
    InMux I__8377 (
            .O(N__41865),
            .I(N__41862));
    LocalMux I__8376 (
            .O(N__41862),
            .I(\serializer_mod_inst.shift_regZ0Z_123 ));
    InMux I__8375 (
            .O(N__41859),
            .I(N__41856));
    LocalMux I__8374 (
            .O(N__41856),
            .I(\serializer_mod_inst.shift_regZ0Z_25 ));
    InMux I__8373 (
            .O(N__41853),
            .I(N__41850));
    LocalMux I__8372 (
            .O(N__41850),
            .I(\serializer_mod_inst.shift_regZ0Z_26 ));
    InMux I__8371 (
            .O(N__41847),
            .I(N__41844));
    LocalMux I__8370 (
            .O(N__41844),
            .I(N__41841));
    Odrv12 I__8369 (
            .O(N__41841),
            .I(\serializer_mod_inst.shift_regZ0Z_6 ));
    InMux I__8368 (
            .O(N__41838),
            .I(N__41835));
    LocalMux I__8367 (
            .O(N__41835),
            .I(\serializer_mod_inst.shift_regZ0Z_5 ));
    InMux I__8366 (
            .O(N__41832),
            .I(N__41829));
    LocalMux I__8365 (
            .O(N__41829),
            .I(\serializer_mod_inst.shift_regZ0Z_2 ));
    InMux I__8364 (
            .O(N__41826),
            .I(N__41823));
    LocalMux I__8363 (
            .O(N__41823),
            .I(\serializer_mod_inst.shift_regZ0Z_3 ));
    InMux I__8362 (
            .O(N__41820),
            .I(N__41817));
    LocalMux I__8361 (
            .O(N__41817),
            .I(\serializer_mod_inst.shift_regZ0Z_4 ));
    InMux I__8360 (
            .O(N__41814),
            .I(N__41811));
    LocalMux I__8359 (
            .O(N__41811),
            .I(\serializer_mod_inst.shift_regZ0Z_21 ));
    InMux I__8358 (
            .O(N__41808),
            .I(N__41803));
    InMux I__8357 (
            .O(N__41807),
            .I(N__41800));
    InMux I__8356 (
            .O(N__41806),
            .I(N__41797));
    LocalMux I__8355 (
            .O(N__41803),
            .I(N__41791));
    LocalMux I__8354 (
            .O(N__41800),
            .I(N__41791));
    LocalMux I__8353 (
            .O(N__41797),
            .I(N__41788));
    InMux I__8352 (
            .O(N__41796),
            .I(N__41783));
    Span12Mux_v I__8351 (
            .O(N__41791),
            .I(N__41778));
    Span12Mux_v I__8350 (
            .O(N__41788),
            .I(N__41778));
    InMux I__8349 (
            .O(N__41787),
            .I(N__41773));
    InMux I__8348 (
            .O(N__41786),
            .I(N__41773));
    LocalMux I__8347 (
            .O(N__41783),
            .I(\I2C_top_level_inst1.s_data_ireg_5 ));
    Odrv12 I__8346 (
            .O(N__41778),
            .I(\I2C_top_level_inst1.s_data_ireg_5 ));
    LocalMux I__8345 (
            .O(N__41773),
            .I(\I2C_top_level_inst1.s_data_ireg_5 ));
    CascadeMux I__8344 (
            .O(N__41766),
            .I(N__41763));
    InMux I__8343 (
            .O(N__41763),
            .I(N__41760));
    LocalMux I__8342 (
            .O(N__41760),
            .I(\I2C_top_level_inst1.s_addr0_o_5 ));
    InMux I__8341 (
            .O(N__41757),
            .I(N__41754));
    LocalMux I__8340 (
            .O(N__41754),
            .I(N__41749));
    InMux I__8339 (
            .O(N__41753),
            .I(N__41746));
    InMux I__8338 (
            .O(N__41752),
            .I(N__41743));
    Span4Mux_v I__8337 (
            .O(N__41749),
            .I(N__41740));
    LocalMux I__8336 (
            .O(N__41746),
            .I(N__41735));
    LocalMux I__8335 (
            .O(N__41743),
            .I(N__41735));
    Span4Mux_h I__8334 (
            .O(N__41740),
            .I(N__41730));
    Span4Mux_v I__8333 (
            .O(N__41735),
            .I(N__41726));
    InMux I__8332 (
            .O(N__41734),
            .I(N__41723));
    InMux I__8331 (
            .O(N__41733),
            .I(N__41720));
    Span4Mux_h I__8330 (
            .O(N__41730),
            .I(N__41717));
    InMux I__8329 (
            .O(N__41729),
            .I(N__41714));
    Odrv4 I__8328 (
            .O(N__41726),
            .I(\I2C_top_level_inst1.s_data_ireg_6 ));
    LocalMux I__8327 (
            .O(N__41723),
            .I(\I2C_top_level_inst1.s_data_ireg_6 ));
    LocalMux I__8326 (
            .O(N__41720),
            .I(\I2C_top_level_inst1.s_data_ireg_6 ));
    Odrv4 I__8325 (
            .O(N__41717),
            .I(\I2C_top_level_inst1.s_data_ireg_6 ));
    LocalMux I__8324 (
            .O(N__41714),
            .I(\I2C_top_level_inst1.s_data_ireg_6 ));
    CascadeMux I__8323 (
            .O(N__41703),
            .I(N__41700));
    InMux I__8322 (
            .O(N__41700),
            .I(N__41697));
    LocalMux I__8321 (
            .O(N__41697),
            .I(N__41694));
    Odrv4 I__8320 (
            .O(N__41694),
            .I(\I2C_top_level_inst1.s_addr0_o_6 ));
    InMux I__8319 (
            .O(N__41691),
            .I(N__41685));
    InMux I__8318 (
            .O(N__41690),
            .I(N__41682));
    InMux I__8317 (
            .O(N__41689),
            .I(N__41679));
    InMux I__8316 (
            .O(N__41688),
            .I(N__41676));
    LocalMux I__8315 (
            .O(N__41685),
            .I(N__41671));
    LocalMux I__8314 (
            .O(N__41682),
            .I(N__41671));
    LocalMux I__8313 (
            .O(N__41679),
            .I(N__41668));
    LocalMux I__8312 (
            .O(N__41676),
            .I(N__41665));
    Span4Mux_v I__8311 (
            .O(N__41671),
            .I(N__41662));
    Span4Mux_v I__8310 (
            .O(N__41668),
            .I(N__41659));
    Span4Mux_h I__8309 (
            .O(N__41665),
            .I(N__41655));
    Span4Mux_h I__8308 (
            .O(N__41662),
            .I(N__41652));
    Sp12to4 I__8307 (
            .O(N__41659),
            .I(N__41649));
    CascadeMux I__8306 (
            .O(N__41658),
            .I(N__41646));
    Span4Mux_h I__8305 (
            .O(N__41655),
            .I(N__41643));
    Sp12to4 I__8304 (
            .O(N__41652),
            .I(N__41638));
    Span12Mux_h I__8303 (
            .O(N__41649),
            .I(N__41638));
    InMux I__8302 (
            .O(N__41646),
            .I(N__41635));
    Odrv4 I__8301 (
            .O(N__41643),
            .I(\I2C_top_level_inst1.s_data_ireg_7 ));
    Odrv12 I__8300 (
            .O(N__41638),
            .I(\I2C_top_level_inst1.s_data_ireg_7 ));
    LocalMux I__8299 (
            .O(N__41635),
            .I(\I2C_top_level_inst1.s_data_ireg_7 ));
    CascadeMux I__8298 (
            .O(N__41628),
            .I(N__41625));
    InMux I__8297 (
            .O(N__41625),
            .I(N__41622));
    LocalMux I__8296 (
            .O(N__41622),
            .I(\I2C_top_level_inst1.s_addr0_o_7 ));
    InMux I__8295 (
            .O(N__41619),
            .I(N__41616));
    LocalMux I__8294 (
            .O(N__41616),
            .I(N__41613));
    Span4Mux_h I__8293 (
            .O(N__41613),
            .I(N__41610));
    Span4Mux_v I__8292 (
            .O(N__41610),
            .I(N__41606));
    InMux I__8291 (
            .O(N__41609),
            .I(N__41603));
    Odrv4 I__8290 (
            .O(N__41606),
            .I(N_396));
    LocalMux I__8289 (
            .O(N__41603),
            .I(N_396));
    CascadeMux I__8288 (
            .O(N__41598),
            .I(N__41595));
    InMux I__8287 (
            .O(N__41595),
            .I(N__41592));
    LocalMux I__8286 (
            .O(N__41592),
            .I(N__41589));
    Span12Mux_h I__8285 (
            .O(N__41589),
            .I(N__41586));
    Odrv12 I__8284 (
            .O(N__41586),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_3 ));
    CascadeMux I__8283 (
            .O(N__41583),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_4_cascade_ ));
    CascadeMux I__8282 (
            .O(N__41580),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNOZ0Z_0_cascade_ ));
    InMux I__8281 (
            .O(N__41577),
            .I(N__41571));
    InMux I__8280 (
            .O(N__41576),
            .I(N__41564));
    InMux I__8279 (
            .O(N__41575),
            .I(N__41564));
    InMux I__8278 (
            .O(N__41574),
            .I(N__41564));
    LocalMux I__8277 (
            .O(N__41571),
            .I(N__41560));
    LocalMux I__8276 (
            .O(N__41564),
            .I(N__41557));
    InMux I__8275 (
            .O(N__41563),
            .I(N__41554));
    Span4Mux_h I__8274 (
            .O(N__41560),
            .I(N__41551));
    Span4Mux_h I__8273 (
            .O(N__41557),
            .I(N__41548));
    LocalMux I__8272 (
            .O(N__41554),
            .I(\I2C_top_level_inst1.s_no_restart ));
    Odrv4 I__8271 (
            .O(N__41551),
            .I(\I2C_top_level_inst1.s_no_restart ));
    Odrv4 I__8270 (
            .O(N__41548),
            .I(\I2C_top_level_inst1.s_no_restart ));
    InMux I__8269 (
            .O(N__41541),
            .I(N__41538));
    LocalMux I__8268 (
            .O(N__41538),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_1 ));
    InMux I__8267 (
            .O(N__41535),
            .I(N__41532));
    LocalMux I__8266 (
            .O(N__41532),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_304_0 ));
    CascadeMux I__8265 (
            .O(N__41529),
            .I(N__41526));
    InMux I__8264 (
            .O(N__41526),
            .I(N__41523));
    LocalMux I__8263 (
            .O(N__41523),
            .I(N__41518));
    InMux I__8262 (
            .O(N__41522),
            .I(N__41512));
    InMux I__8261 (
            .O(N__41521),
            .I(N__41512));
    Span4Mux_v I__8260 (
            .O(N__41518),
            .I(N__41509));
    CascadeMux I__8259 (
            .O(N__41517),
            .I(N__41506));
    LocalMux I__8258 (
            .O(N__41512),
            .I(N__41503));
    Span4Mux_h I__8257 (
            .O(N__41509),
            .I(N__41500));
    InMux I__8256 (
            .O(N__41506),
            .I(N__41497));
    Span4Mux_h I__8255 (
            .O(N__41503),
            .I(N__41494));
    Odrv4 I__8254 (
            .O(N__41500),
            .I(\I2C_top_level_inst1.s_ack ));
    LocalMux I__8253 (
            .O(N__41497),
            .I(\I2C_top_level_inst1.s_ack ));
    Odrv4 I__8252 (
            .O(N__41494),
            .I(\I2C_top_level_inst1.s_ack ));
    CascadeMux I__8251 (
            .O(N__41487),
            .I(N__41484));
    InMux I__8250 (
            .O(N__41484),
            .I(N__41481));
    LocalMux I__8249 (
            .O(N__41481),
            .I(N__41478));
    Span4Mux_v I__8248 (
            .O(N__41478),
            .I(N__41475));
    Span4Mux_h I__8247 (
            .O(N__41475),
            .I(N__41472));
    Odrv4 I__8246 (
            .O(N__41472),
            .I(\I2C_top_level_inst1.s_addr1_o_4 ));
    CascadeMux I__8245 (
            .O(N__41469),
            .I(N__41466));
    InMux I__8244 (
            .O(N__41466),
            .I(N__41463));
    LocalMux I__8243 (
            .O(N__41463),
            .I(N__41460));
    Span4Mux_h I__8242 (
            .O(N__41460),
            .I(N__41457));
    Odrv4 I__8241 (
            .O(N__41457),
            .I(\I2C_top_level_inst1.s_addr1_o_5 ));
    CascadeMux I__8240 (
            .O(N__41454),
            .I(N__41451));
    InMux I__8239 (
            .O(N__41451),
            .I(N__41448));
    LocalMux I__8238 (
            .O(N__41448),
            .I(N__41445));
    Span4Mux_h I__8237 (
            .O(N__41445),
            .I(N__41442));
    Odrv4 I__8236 (
            .O(N__41442),
            .I(\I2C_top_level_inst1.s_addr1_o_6 ));
    CascadeMux I__8235 (
            .O(N__41439),
            .I(N__41436));
    InMux I__8234 (
            .O(N__41436),
            .I(N__41433));
    LocalMux I__8233 (
            .O(N__41433),
            .I(N__41430));
    Span4Mux_v I__8232 (
            .O(N__41430),
            .I(N__41427));
    Odrv4 I__8231 (
            .O(N__41427),
            .I(\I2C_top_level_inst1.s_addr1_o_7 ));
    InMux I__8230 (
            .O(N__41424),
            .I(N__41421));
    LocalMux I__8229 (
            .O(N__41421),
            .I(N__41417));
    CEMux I__8228 (
            .O(N__41420),
            .I(N__41414));
    Span4Mux_h I__8227 (
            .O(N__41417),
            .I(N__41410));
    LocalMux I__8226 (
            .O(N__41414),
            .I(N__41407));
    InMux I__8225 (
            .O(N__41413),
            .I(N__41403));
    Sp12to4 I__8224 (
            .O(N__41410),
            .I(N__41400));
    Span4Mux_h I__8223 (
            .O(N__41407),
            .I(N__41397));
    InMux I__8222 (
            .O(N__41406),
            .I(N__41394));
    LocalMux I__8221 (
            .O(N__41403),
            .I(\I2C_top_level_inst1.s_load_addr1 ));
    Odrv12 I__8220 (
            .O(N__41400),
            .I(\I2C_top_level_inst1.s_load_addr1 ));
    Odrv4 I__8219 (
            .O(N__41397),
            .I(\I2C_top_level_inst1.s_load_addr1 ));
    LocalMux I__8218 (
            .O(N__41394),
            .I(\I2C_top_level_inst1.s_load_addr1 ));
    InMux I__8217 (
            .O(N__41385),
            .I(N__41382));
    LocalMux I__8216 (
            .O(N__41382),
            .I(\I2C_top_level_inst1.s_addr0_o_3 ));
    InMux I__8215 (
            .O(N__41379),
            .I(N__41372));
    InMux I__8214 (
            .O(N__41378),
            .I(N__41369));
    InMux I__8213 (
            .O(N__41377),
            .I(N__41366));
    InMux I__8212 (
            .O(N__41376),
            .I(N__41363));
    InMux I__8211 (
            .O(N__41375),
            .I(N__41360));
    LocalMux I__8210 (
            .O(N__41372),
            .I(N__41355));
    LocalMux I__8209 (
            .O(N__41369),
            .I(N__41355));
    LocalMux I__8208 (
            .O(N__41366),
            .I(N__41352));
    LocalMux I__8207 (
            .O(N__41363),
            .I(N__41349));
    LocalMux I__8206 (
            .O(N__41360),
            .I(N__41343));
    Span4Mux_v I__8205 (
            .O(N__41355),
            .I(N__41343));
    Span4Mux_h I__8204 (
            .O(N__41352),
            .I(N__41338));
    Span4Mux_v I__8203 (
            .O(N__41349),
            .I(N__41338));
    InMux I__8202 (
            .O(N__41348),
            .I(N__41335));
    Odrv4 I__8201 (
            .O(N__41343),
            .I(\I2C_top_level_inst1.s_data_ireg_4 ));
    Odrv4 I__8200 (
            .O(N__41338),
            .I(\I2C_top_level_inst1.s_data_ireg_4 ));
    LocalMux I__8199 (
            .O(N__41335),
            .I(\I2C_top_level_inst1.s_data_ireg_4 ));
    CascadeMux I__8198 (
            .O(N__41328),
            .I(N__41325));
    InMux I__8197 (
            .O(N__41325),
            .I(N__41322));
    LocalMux I__8196 (
            .O(N__41322),
            .I(N__41319));
    Odrv4 I__8195 (
            .O(N__41319),
            .I(\I2C_top_level_inst1.s_addr0_o_4 ));
    CascadeMux I__8194 (
            .O(N__41316),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0_cascade_ ));
    CascadeMux I__8193 (
            .O(N__41313),
            .I(N__41310));
    InMux I__8192 (
            .O(N__41310),
            .I(N__41307));
    LocalMux I__8191 (
            .O(N__41307),
            .I(\I2C_top_level_inst1.s_addr1_o_1 ));
    InMux I__8190 (
            .O(N__41304),
            .I(N__41301));
    LocalMux I__8189 (
            .O(N__41301),
            .I(\I2C_top_level_inst1.s_addr1_o_2 ));
    InMux I__8188 (
            .O(N__41298),
            .I(N__41295));
    LocalMux I__8187 (
            .O(N__41295),
            .I(\I2C_top_level_inst1.s_addr1_o_3 ));
    InMux I__8186 (
            .O(N__41292),
            .I(N__41289));
    LocalMux I__8185 (
            .O(N__41289),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11 ));
    CascadeMux I__8184 (
            .O(N__41286),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11_cascade_ ));
    InMux I__8183 (
            .O(N__41283),
            .I(N__41280));
    LocalMux I__8182 (
            .O(N__41280),
            .I(N__41277));
    Odrv12 I__8181 (
            .O(N__41277),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_12 ));
    CascadeMux I__8180 (
            .O(N__41274),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GHZ0Z5_cascade_ ));
    InMux I__8179 (
            .O(N__41271),
            .I(N__41268));
    LocalMux I__8178 (
            .O(N__41268),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12 ));
    InMux I__8177 (
            .O(N__41265),
            .I(N__41262));
    LocalMux I__8176 (
            .O(N__41262),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_11 ));
    CascadeMux I__8175 (
            .O(N__41259),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12_cascade_ ));
    InMux I__8174 (
            .O(N__41256),
            .I(N__41253));
    LocalMux I__8173 (
            .O(N__41253),
            .I(N__41250));
    Span4Mux_v I__8172 (
            .O(N__41250),
            .I(N__41247));
    Span4Mux_h I__8171 (
            .O(N__41247),
            .I(N__41244));
    Span4Mux_h I__8170 (
            .O(N__41244),
            .I(N__41241));
    Odrv4 I__8169 (
            .O(N__41241),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_12 ));
    CascadeMux I__8168 (
            .O(N__41238),
            .I(N__41235));
    InMux I__8167 (
            .O(N__41235),
            .I(N__41231));
    InMux I__8166 (
            .O(N__41234),
            .I(N__41228));
    LocalMux I__8165 (
            .O(N__41231),
            .I(N__41225));
    LocalMux I__8164 (
            .O(N__41228),
            .I(N__41222));
    Span4Mux_v I__8163 (
            .O(N__41225),
            .I(N__41218));
    Span4Mux_v I__8162 (
            .O(N__41222),
            .I(N__41215));
    InMux I__8161 (
            .O(N__41221),
            .I(N__41212));
    Span4Mux_h I__8160 (
            .O(N__41218),
            .I(N__41209));
    Odrv4 I__8159 (
            .O(N__41215),
            .I(cemf_module_64ch_ctrl_inst1_data_config_12));
    LocalMux I__8158 (
            .O(N__41212),
            .I(cemf_module_64ch_ctrl_inst1_data_config_12));
    Odrv4 I__8157 (
            .O(N__41209),
            .I(cemf_module_64ch_ctrl_inst1_data_config_12));
    InMux I__8156 (
            .O(N__41202),
            .I(N__41198));
    InMux I__8155 (
            .O(N__41201),
            .I(N__41194));
    LocalMux I__8154 (
            .O(N__41198),
            .I(N__41191));
    CascadeMux I__8153 (
            .O(N__41197),
            .I(N__41188));
    LocalMux I__8152 (
            .O(N__41194),
            .I(N__41185));
    Span4Mux_h I__8151 (
            .O(N__41191),
            .I(N__41182));
    InMux I__8150 (
            .O(N__41188),
            .I(N__41179));
    Span4Mux_v I__8149 (
            .O(N__41185),
            .I(N__41176));
    Odrv4 I__8148 (
            .O(N__41182),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_12));
    LocalMux I__8147 (
            .O(N__41179),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_12));
    Odrv4 I__8146 (
            .O(N__41176),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_12));
    CascadeMux I__8145 (
            .O(N__41169),
            .I(N__41166));
    InMux I__8144 (
            .O(N__41166),
            .I(N__41163));
    LocalMux I__8143 (
            .O(N__41163),
            .I(N__41160));
    Odrv4 I__8142 (
            .O(N__41160),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_12 ));
    CascadeMux I__8141 (
            .O(N__41157),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_11_cascade_ ));
    InMux I__8140 (
            .O(N__41154),
            .I(N__41151));
    LocalMux I__8139 (
            .O(N__41151),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFHZ0Z5 ));
    CascadeMux I__8138 (
            .O(N__41148),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13_cascade_ ));
    InMux I__8137 (
            .O(N__41145),
            .I(N__41142));
    LocalMux I__8136 (
            .O(N__41142),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_12 ));
    InMux I__8135 (
            .O(N__41139),
            .I(N__41136));
    LocalMux I__8134 (
            .O(N__41136),
            .I(N__41133));
    Span4Mux_h I__8133 (
            .O(N__41133),
            .I(N__41130));
    Odrv4 I__8132 (
            .O(N__41130),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_13 ));
    InMux I__8131 (
            .O(N__41127),
            .I(N__41122));
    CascadeMux I__8130 (
            .O(N__41126),
            .I(N__41119));
    CascadeMux I__8129 (
            .O(N__41125),
            .I(N__41116));
    LocalMux I__8128 (
            .O(N__41122),
            .I(N__41113));
    InMux I__8127 (
            .O(N__41119),
            .I(N__41110));
    InMux I__8126 (
            .O(N__41116),
            .I(N__41107));
    Span4Mux_v I__8125 (
            .O(N__41113),
            .I(N__41104));
    LocalMux I__8124 (
            .O(N__41110),
            .I(N__41101));
    LocalMux I__8123 (
            .O(N__41107),
            .I(N__41098));
    Span4Mux_h I__8122 (
            .O(N__41104),
            .I(N__41093));
    Span4Mux_v I__8121 (
            .O(N__41101),
            .I(N__41093));
    Odrv12 I__8120 (
            .O(N__41098),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_5));
    Odrv4 I__8119 (
            .O(N__41093),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_5));
    CascadeMux I__8118 (
            .O(N__41088),
            .I(N__41084));
    InMux I__8117 (
            .O(N__41087),
            .I(N__41078));
    InMux I__8116 (
            .O(N__41084),
            .I(N__41078));
    InMux I__8115 (
            .O(N__41083),
            .I(N__41075));
    LocalMux I__8114 (
            .O(N__41078),
            .I(N__41072));
    LocalMux I__8113 (
            .O(N__41075),
            .I(N__41067));
    Span4Mux_v I__8112 (
            .O(N__41072),
            .I(N__41067));
    Span4Mux_v I__8111 (
            .O(N__41067),
            .I(N__41064));
    Span4Mux_h I__8110 (
            .O(N__41064),
            .I(N__41061));
    Odrv4 I__8109 (
            .O(N__41061),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_6));
    InMux I__8108 (
            .O(N__41058),
            .I(N__41055));
    LocalMux I__8107 (
            .O(N__41055),
            .I(N__41050));
    CascadeMux I__8106 (
            .O(N__41054),
            .I(N__41047));
    CascadeMux I__8105 (
            .O(N__41053),
            .I(N__41044));
    Span12Mux_v I__8104 (
            .O(N__41050),
            .I(N__41041));
    InMux I__8103 (
            .O(N__41047),
            .I(N__41038));
    InMux I__8102 (
            .O(N__41044),
            .I(N__41035));
    Span12Mux_h I__8101 (
            .O(N__41041),
            .I(N__41028));
    LocalMux I__8100 (
            .O(N__41038),
            .I(N__41028));
    LocalMux I__8099 (
            .O(N__41035),
            .I(N__41028));
    Odrv12 I__8098 (
            .O(N__41028),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_7));
    InMux I__8097 (
            .O(N__41025),
            .I(N__41022));
    LocalMux I__8096 (
            .O(N__41022),
            .I(N__41017));
    CascadeMux I__8095 (
            .O(N__41021),
            .I(N__41014));
    CascadeMux I__8094 (
            .O(N__41020),
            .I(N__41011));
    Span4Mux_h I__8093 (
            .O(N__41017),
            .I(N__41008));
    InMux I__8092 (
            .O(N__41014),
            .I(N__41005));
    InMux I__8091 (
            .O(N__41011),
            .I(N__41002));
    Span4Mux_h I__8090 (
            .O(N__41008),
            .I(N__40997));
    LocalMux I__8089 (
            .O(N__41005),
            .I(N__40997));
    LocalMux I__8088 (
            .O(N__41002),
            .I(N__40994));
    Span4Mux_v I__8087 (
            .O(N__40997),
            .I(N__40991));
    Odrv4 I__8086 (
            .O(N__40994),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_8));
    Odrv4 I__8085 (
            .O(N__40991),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_8));
    InMux I__8084 (
            .O(N__40986),
            .I(N__40982));
    InMux I__8083 (
            .O(N__40985),
            .I(N__40979));
    LocalMux I__8082 (
            .O(N__40982),
            .I(N__40974));
    LocalMux I__8081 (
            .O(N__40979),
            .I(N__40974));
    Span4Mux_h I__8080 (
            .O(N__40974),
            .I(N__40970));
    InMux I__8079 (
            .O(N__40973),
            .I(N__40967));
    Odrv4 I__8078 (
            .O(N__40970),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_20));
    LocalMux I__8077 (
            .O(N__40967),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_20));
    CascadeMux I__8076 (
            .O(N__40962),
            .I(N__40958));
    InMux I__8075 (
            .O(N__40961),
            .I(N__40954));
    InMux I__8074 (
            .O(N__40958),
            .I(N__40949));
    InMux I__8073 (
            .O(N__40957),
            .I(N__40949));
    LocalMux I__8072 (
            .O(N__40954),
            .I(N__40946));
    LocalMux I__8071 (
            .O(N__40949),
            .I(N__40943));
    Span4Mux_v I__8070 (
            .O(N__40946),
            .I(N__40938));
    Span4Mux_h I__8069 (
            .O(N__40943),
            .I(N__40938));
    Odrv4 I__8068 (
            .O(N__40938),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_12));
    CascadeMux I__8067 (
            .O(N__40935),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_0_12_cascade_ ));
    InMux I__8066 (
            .O(N__40932),
            .I(N__40929));
    LocalMux I__8065 (
            .O(N__40929),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_2_12 ));
    CascadeMux I__8064 (
            .O(N__40926),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_0_i_12_cascade_ ));
    InMux I__8063 (
            .O(N__40923),
            .I(N__40920));
    LocalMux I__8062 (
            .O(N__40920),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12 ));
    CascadeMux I__8061 (
            .O(N__40917),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12_cascade_ ));
    InMux I__8060 (
            .O(N__40914),
            .I(N__40911));
    LocalMux I__8059 (
            .O(N__40911),
            .I(N__40908));
    Span4Mux_h I__8058 (
            .O(N__40908),
            .I(N__40905));
    Span4Mux_v I__8057 (
            .O(N__40905),
            .I(N__40902));
    Span4Mux_h I__8056 (
            .O(N__40902),
            .I(N__40899));
    Odrv4 I__8055 (
            .O(N__40899),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_13 ));
    CascadeMux I__8054 (
            .O(N__40896),
            .I(N__40893));
    InMux I__8053 (
            .O(N__40893),
            .I(N__40889));
    CascadeMux I__8052 (
            .O(N__40892),
            .I(N__40885));
    LocalMux I__8051 (
            .O(N__40889),
            .I(N__40882));
    InMux I__8050 (
            .O(N__40888),
            .I(N__40879));
    InMux I__8049 (
            .O(N__40885),
            .I(N__40876));
    Span4Mux_v I__8048 (
            .O(N__40882),
            .I(N__40871));
    LocalMux I__8047 (
            .O(N__40879),
            .I(N__40871));
    LocalMux I__8046 (
            .O(N__40876),
            .I(N__40868));
    Span4Mux_h I__8045 (
            .O(N__40871),
            .I(N__40865));
    Odrv12 I__8044 (
            .O(N__40868),
            .I(cemf_module_64ch_ctrl_inst1_data_config_13));
    Odrv4 I__8043 (
            .O(N__40865),
            .I(cemf_module_64ch_ctrl_inst1_data_config_13));
    CascadeMux I__8042 (
            .O(N__40860),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8DZ0Z7_cascade_ ));
    InMux I__8041 (
            .O(N__40857),
            .I(N__40854));
    LocalMux I__8040 (
            .O(N__40854),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13 ));
    InMux I__8039 (
            .O(N__40851),
            .I(N__40848));
    LocalMux I__8038 (
            .O(N__40848),
            .I(N__40845));
    Odrv4 I__8037 (
            .O(N__40845),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8DZ0Z7 ));
    InMux I__8036 (
            .O(N__40842),
            .I(N__40839));
    LocalMux I__8035 (
            .O(N__40839),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14 ));
    CascadeMux I__8034 (
            .O(N__40836),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14_cascade_ ));
    InMux I__8033 (
            .O(N__40833),
            .I(N__40830));
    LocalMux I__8032 (
            .O(N__40830),
            .I(N__40827));
    Span4Mux_h I__8031 (
            .O(N__40827),
            .I(N__40824));
    Span4Mux_v I__8030 (
            .O(N__40824),
            .I(N__40819));
    InMux I__8029 (
            .O(N__40823),
            .I(N__40816));
    InMux I__8028 (
            .O(N__40822),
            .I(N__40813));
    Odrv4 I__8027 (
            .O(N__40819),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_8));
    LocalMux I__8026 (
            .O(N__40816),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_8));
    LocalMux I__8025 (
            .O(N__40813),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_8));
    InMux I__8024 (
            .O(N__40806),
            .I(N__40803));
    LocalMux I__8023 (
            .O(N__40803),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_8 ));
    InMux I__8022 (
            .O(N__40800),
            .I(N__40797));
    LocalMux I__8021 (
            .O(N__40797),
            .I(N__40794));
    Odrv4 I__8020 (
            .O(N__40794),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_20 ));
    InMux I__8019 (
            .O(N__40791),
            .I(N__40788));
    LocalMux I__8018 (
            .O(N__40788),
            .I(N__40785));
    Odrv12 I__8017 (
            .O(N__40785),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_3 ));
    InMux I__8016 (
            .O(N__40782),
            .I(N__40779));
    LocalMux I__8015 (
            .O(N__40779),
            .I(N__40776));
    Odrv4 I__8014 (
            .O(N__40776),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_8 ));
    CascadeMux I__8013 (
            .O(N__40773),
            .I(N__40770));
    InMux I__8012 (
            .O(N__40770),
            .I(N__40767));
    LocalMux I__8011 (
            .O(N__40767),
            .I(N__40763));
    InMux I__8010 (
            .O(N__40766),
            .I(N__40760));
    Span4Mux_v I__8009 (
            .O(N__40763),
            .I(N__40754));
    LocalMux I__8008 (
            .O(N__40760),
            .I(N__40754));
    InMux I__8007 (
            .O(N__40759),
            .I(N__40751));
    Span4Mux_h I__8006 (
            .O(N__40754),
            .I(N__40748));
    LocalMux I__8005 (
            .O(N__40751),
            .I(N__40745));
    Span4Mux_v I__8004 (
            .O(N__40748),
            .I(N__40742));
    Span4Mux_h I__8003 (
            .O(N__40745),
            .I(N__40739));
    Sp12to4 I__8002 (
            .O(N__40742),
            .I(N__40736));
    Odrv4 I__8001 (
            .O(N__40739),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_8));
    Odrv12 I__8000 (
            .O(N__40736),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_8));
    InMux I__7999 (
            .O(N__40731),
            .I(N__40728));
    LocalMux I__7998 (
            .O(N__40728),
            .I(N__40725));
    Span4Mux_h I__7997 (
            .O(N__40725),
            .I(N__40722));
    Span4Mux_h I__7996 (
            .O(N__40722),
            .I(N__40718));
    InMux I__7995 (
            .O(N__40721),
            .I(N__40714));
    Span4Mux_v I__7994 (
            .O(N__40718),
            .I(N__40711));
    InMux I__7993 (
            .O(N__40717),
            .I(N__40708));
    LocalMux I__7992 (
            .O(N__40714),
            .I(N__40705));
    Odrv4 I__7991 (
            .O(N__40711),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_8));
    LocalMux I__7990 (
            .O(N__40708),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_8));
    Odrv4 I__7989 (
            .O(N__40705),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_8));
    InMux I__7988 (
            .O(N__40698),
            .I(N__40693));
    InMux I__7987 (
            .O(N__40697),
            .I(N__40690));
    InMux I__7986 (
            .O(N__40696),
            .I(N__40687));
    LocalMux I__7985 (
            .O(N__40693),
            .I(N__40684));
    LocalMux I__7984 (
            .O(N__40690),
            .I(N__40681));
    LocalMux I__7983 (
            .O(N__40687),
            .I(N__40678));
    Span4Mux_h I__7982 (
            .O(N__40684),
            .I(N__40675));
    Span4Mux_h I__7981 (
            .O(N__40681),
            .I(N__40672));
    Span4Mux_h I__7980 (
            .O(N__40678),
            .I(N__40669));
    Span4Mux_v I__7979 (
            .O(N__40675),
            .I(N__40666));
    Span4Mux_h I__7978 (
            .O(N__40672),
            .I(N__40663));
    Span4Mux_h I__7977 (
            .O(N__40669),
            .I(N__40660));
    Odrv4 I__7976 (
            .O(N__40666),
            .I(cemf_module_64ch_ctrl_inst1_data_config_8));
    Odrv4 I__7975 (
            .O(N__40663),
            .I(cemf_module_64ch_ctrl_inst1_data_config_8));
    Odrv4 I__7974 (
            .O(N__40660),
            .I(cemf_module_64ch_ctrl_inst1_data_config_8));
    CascadeMux I__7973 (
            .O(N__40653),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_8_cascade_ ));
    CascadeMux I__7972 (
            .O(N__40650),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SLZ0Z7_cascade_ ));
    InMux I__7971 (
            .O(N__40647),
            .I(N__40644));
    LocalMux I__7970 (
            .O(N__40644),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8 ));
    InMux I__7969 (
            .O(N__40641),
            .I(N__40638));
    LocalMux I__7968 (
            .O(N__40638),
            .I(N__40635));
    Span4Mux_v I__7967 (
            .O(N__40635),
            .I(N__40632));
    Span4Mux_h I__7966 (
            .O(N__40632),
            .I(N__40629));
    Odrv4 I__7965 (
            .O(N__40629),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_7 ));
    CascadeMux I__7964 (
            .O(N__40626),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8_cascade_ ));
    CascadeMux I__7963 (
            .O(N__40623),
            .I(N__40620));
    InMux I__7962 (
            .O(N__40620),
            .I(N__40617));
    LocalMux I__7961 (
            .O(N__40617),
            .I(N__40614));
    Span4Mux_h I__7960 (
            .O(N__40614),
            .I(N__40611));
    Span4Mux_h I__7959 (
            .O(N__40611),
            .I(N__40608));
    Sp12to4 I__7958 (
            .O(N__40608),
            .I(N__40605));
    Odrv12 I__7957 (
            .O(N__40605),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_28));
    InMux I__7956 (
            .O(N__40602),
            .I(N__40599));
    LocalMux I__7955 (
            .O(N__40599),
            .I(N__40596));
    Span4Mux_v I__7954 (
            .O(N__40596),
            .I(N__40593));
    Span4Mux_v I__7953 (
            .O(N__40593),
            .I(N__40590));
    Sp12to4 I__7952 (
            .O(N__40590),
            .I(N__40587));
    Odrv12 I__7951 (
            .O(N__40587),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_1Z0Z_26 ));
    CascadeMux I__7950 (
            .O(N__40584),
            .I(N__40581));
    InMux I__7949 (
            .O(N__40581),
            .I(N__40578));
    LocalMux I__7948 (
            .O(N__40578),
            .I(N__40575));
    Span4Mux_h I__7947 (
            .O(N__40575),
            .I(N__40572));
    Odrv4 I__7946 (
            .O(N__40572),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_27));
    InMux I__7945 (
            .O(N__40569),
            .I(N__40566));
    LocalMux I__7944 (
            .O(N__40566),
            .I(N__40563));
    Odrv4 I__7943 (
            .O(N__40563),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_7 ));
    InMux I__7942 (
            .O(N__40560),
            .I(N__40557));
    LocalMux I__7941 (
            .O(N__40557),
            .I(N__40554));
    Odrv12 I__7940 (
            .O(N__40554),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_7 ));
    InMux I__7939 (
            .O(N__40551),
            .I(N__40548));
    LocalMux I__7938 (
            .O(N__40548),
            .I(N__40545));
    Span12Mux_h I__7937 (
            .O(N__40545),
            .I(N__40540));
    InMux I__7936 (
            .O(N__40544),
            .I(N__40535));
    InMux I__7935 (
            .O(N__40543),
            .I(N__40535));
    Odrv12 I__7934 (
            .O(N__40540),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_7));
    LocalMux I__7933 (
            .O(N__40535),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_7));
    CascadeMux I__7932 (
            .O(N__40530),
            .I(N__40526));
    InMux I__7931 (
            .O(N__40529),
            .I(N__40523));
    InMux I__7930 (
            .O(N__40526),
            .I(N__40520));
    LocalMux I__7929 (
            .O(N__40523),
            .I(N__40517));
    LocalMux I__7928 (
            .O(N__40520),
            .I(N__40514));
    Span4Mux_h I__7927 (
            .O(N__40517),
            .I(N__40511));
    Span4Mux_h I__7926 (
            .O(N__40514),
            .I(N__40507));
    Span4Mux_h I__7925 (
            .O(N__40511),
            .I(N__40504));
    InMux I__7924 (
            .O(N__40510),
            .I(N__40501));
    Span4Mux_h I__7923 (
            .O(N__40507),
            .I(N__40498));
    Odrv4 I__7922 (
            .O(N__40504),
            .I(cemf_module_64ch_ctrl_inst1_data_config_7));
    LocalMux I__7921 (
            .O(N__40501),
            .I(cemf_module_64ch_ctrl_inst1_data_config_7));
    Odrv4 I__7920 (
            .O(N__40498),
            .I(cemf_module_64ch_ctrl_inst1_data_config_7));
    CascadeMux I__7919 (
            .O(N__40491),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_8_cascade_ ));
    CascadeMux I__7918 (
            .O(N__40488),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3QZ0Z5_cascade_ ));
    InMux I__7917 (
            .O(N__40485),
            .I(N__40482));
    LocalMux I__7916 (
            .O(N__40482),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8 ));
    CascadeMux I__7915 (
            .O(N__40479),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8_cascade_ ));
    CascadeMux I__7914 (
            .O(N__40476),
            .I(N__40473));
    InMux I__7913 (
            .O(N__40473),
            .I(N__40470));
    LocalMux I__7912 (
            .O(N__40470),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_7 ));
    CascadeMux I__7911 (
            .O(N__40467),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3QZ0Z5_cascade_ ));
    InMux I__7910 (
            .O(N__40464),
            .I(N__40461));
    LocalMux I__7909 (
            .O(N__40461),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7 ));
    InMux I__7908 (
            .O(N__40458),
            .I(N__40455));
    LocalMux I__7907 (
            .O(N__40455),
            .I(N__40452));
    Span12Mux_v I__7906 (
            .O(N__40452),
            .I(N__40449));
    Odrv12 I__7905 (
            .O(N__40449),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_6 ));
    CascadeMux I__7904 (
            .O(N__40446),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7_cascade_ ));
    InMux I__7903 (
            .O(N__40443),
            .I(N__40440));
    LocalMux I__7902 (
            .O(N__40440),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_7 ));
    CascadeMux I__7901 (
            .O(N__40437),
            .I(N__40434));
    InMux I__7900 (
            .O(N__40434),
            .I(N__40431));
    LocalMux I__7899 (
            .O(N__40431),
            .I(N__40428));
    Span4Mux_v I__7898 (
            .O(N__40428),
            .I(N__40425));
    Odrv4 I__7897 (
            .O(N__40425),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_24));
    InMux I__7896 (
            .O(N__40422),
            .I(N__40419));
    LocalMux I__7895 (
            .O(N__40419),
            .I(N__40416));
    Odrv4 I__7894 (
            .O(N__40416),
            .I(\serializer_mod_inst.shift_regZ0Z_82 ));
    InMux I__7893 (
            .O(N__40413),
            .I(N__40410));
    LocalMux I__7892 (
            .O(N__40410),
            .I(N__40407));
    Span4Mux_h I__7891 (
            .O(N__40407),
            .I(N__40404));
    Odrv4 I__7890 (
            .O(N__40404),
            .I(\serializer_mod_inst.shift_regZ0Z_80 ));
    InMux I__7889 (
            .O(N__40401),
            .I(N__40398));
    LocalMux I__7888 (
            .O(N__40398),
            .I(\serializer_mod_inst.shift_regZ0Z_81 ));
    InMux I__7887 (
            .O(N__40395),
            .I(N__40392));
    LocalMux I__7886 (
            .O(N__40392),
            .I(N__40389));
    Span4Mux_v I__7885 (
            .O(N__40389),
            .I(N__40386));
    Span4Mux_h I__7884 (
            .O(N__40386),
            .I(N__40383));
    Span4Mux_h I__7883 (
            .O(N__40383),
            .I(N__40380));
    Span4Mux_v I__7882 (
            .O(N__40380),
            .I(N__40377));
    Odrv4 I__7881 (
            .O(N__40377),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_29));
    CascadeMux I__7880 (
            .O(N__40374),
            .I(N__40371));
    InMux I__7879 (
            .O(N__40371),
            .I(N__40368));
    LocalMux I__7878 (
            .O(N__40368),
            .I(N__40365));
    Span4Mux_v I__7877 (
            .O(N__40365),
            .I(N__40362));
    Span4Mux_h I__7876 (
            .O(N__40362),
            .I(N__40359));
    Span4Mux_h I__7875 (
            .O(N__40359),
            .I(N__40356));
    Odrv4 I__7874 (
            .O(N__40356),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_29));
    CascadeMux I__7873 (
            .O(N__40353),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_29_cascade_ ));
    InMux I__7872 (
            .O(N__40350),
            .I(N__40347));
    LocalMux I__7871 (
            .O(N__40347),
            .I(N__40344));
    Span4Mux_v I__7870 (
            .O(N__40344),
            .I(N__40341));
    Span4Mux_h I__7869 (
            .O(N__40341),
            .I(N__40338));
    Odrv4 I__7868 (
            .O(N__40338),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_29 ));
    InMux I__7867 (
            .O(N__40335),
            .I(N__40332));
    LocalMux I__7866 (
            .O(N__40332),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_29 ));
    CascadeMux I__7865 (
            .O(N__40329),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_29_cascade_ ));
    InMux I__7864 (
            .O(N__40326),
            .I(N__40323));
    LocalMux I__7863 (
            .O(N__40323),
            .I(N__40320));
    Span4Mux_h I__7862 (
            .O(N__40320),
            .I(N__40317));
    Span4Mux_h I__7861 (
            .O(N__40317),
            .I(N__40314));
    Odrv4 I__7860 (
            .O(N__40314),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_632 ));
    InMux I__7859 (
            .O(N__40311),
            .I(N__40308));
    LocalMux I__7858 (
            .O(N__40308),
            .I(N__40305));
    Span4Mux_h I__7857 (
            .O(N__40305),
            .I(N__40302));
    Span4Mux_h I__7856 (
            .O(N__40302),
            .I(N__40299));
    Odrv4 I__7855 (
            .O(N__40299),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_29 ));
    InMux I__7854 (
            .O(N__40296),
            .I(N__40293));
    LocalMux I__7853 (
            .O(N__40293),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_29 ));
    InMux I__7852 (
            .O(N__40290),
            .I(N__40287));
    LocalMux I__7851 (
            .O(N__40287),
            .I(\serializer_mod_inst.shift_regZ0Z_42 ));
    InMux I__7850 (
            .O(N__40284),
            .I(N__40281));
    LocalMux I__7849 (
            .O(N__40281),
            .I(\serializer_mod_inst.shift_regZ0Z_43 ));
    InMux I__7848 (
            .O(N__40278),
            .I(N__40275));
    LocalMux I__7847 (
            .O(N__40275),
            .I(\serializer_mod_inst.shift_regZ0Z_44 ));
    InMux I__7846 (
            .O(N__40272),
            .I(N__40269));
    LocalMux I__7845 (
            .O(N__40269),
            .I(N__40266));
    Odrv4 I__7844 (
            .O(N__40266),
            .I(\serializer_mod_inst.shift_regZ0Z_45 ));
    InMux I__7843 (
            .O(N__40263),
            .I(N__40260));
    LocalMux I__7842 (
            .O(N__40260),
            .I(\serializer_mod_inst.shift_regZ0Z_70 ));
    InMux I__7841 (
            .O(N__40257),
            .I(N__40254));
    LocalMux I__7840 (
            .O(N__40254),
            .I(\serializer_mod_inst.shift_regZ0Z_71 ));
    InMux I__7839 (
            .O(N__40251),
            .I(N__40248));
    LocalMux I__7838 (
            .O(N__40248),
            .I(\serializer_mod_inst.shift_regZ0Z_74 ));
    InMux I__7837 (
            .O(N__40245),
            .I(N__40242));
    LocalMux I__7836 (
            .O(N__40242),
            .I(N__40239));
    Odrv4 I__7835 (
            .O(N__40239),
            .I(\serializer_mod_inst.shift_regZ0Z_75 ));
    InMux I__7834 (
            .O(N__40236),
            .I(N__40233));
    LocalMux I__7833 (
            .O(N__40233),
            .I(N__40230));
    Odrv4 I__7832 (
            .O(N__40230),
            .I(\serializer_mod_inst.shift_regZ0Z_98 ));
    InMux I__7831 (
            .O(N__40227),
            .I(N__40224));
    LocalMux I__7830 (
            .O(N__40224),
            .I(N__40221));
    Odrv4 I__7829 (
            .O(N__40221),
            .I(\serializer_mod_inst.shift_regZ0Z_99 ));
    InMux I__7828 (
            .O(N__40218),
            .I(N__40215));
    LocalMux I__7827 (
            .O(N__40215),
            .I(\serializer_mod_inst.shift_regZ0Z_72 ));
    InMux I__7826 (
            .O(N__40212),
            .I(N__40209));
    LocalMux I__7825 (
            .O(N__40209),
            .I(\serializer_mod_inst.shift_regZ0Z_73 ));
    CascadeMux I__7824 (
            .O(N__40206),
            .I(N__40203));
    InMux I__7823 (
            .O(N__40203),
            .I(N__40200));
    LocalMux I__7822 (
            .O(N__40200),
            .I(\serializer_mod_inst.shift_regZ0Z_83 ));
    InMux I__7821 (
            .O(N__40197),
            .I(N__40194));
    LocalMux I__7820 (
            .O(N__40194),
            .I(N__40191));
    Odrv4 I__7819 (
            .O(N__40191),
            .I(\serializer_mod_inst.shift_regZ0Z_85 ));
    InMux I__7818 (
            .O(N__40188),
            .I(N__40185));
    LocalMux I__7817 (
            .O(N__40185),
            .I(\serializer_mod_inst.shift_regZ0Z_1 ));
    InMux I__7816 (
            .O(N__40182),
            .I(N__40179));
    LocalMux I__7815 (
            .O(N__40179),
            .I(\serializer_mod_inst.shift_regZ0Z_101 ));
    InMux I__7814 (
            .O(N__40176),
            .I(N__40173));
    LocalMux I__7813 (
            .O(N__40173),
            .I(N__40170));
    Span4Mux_h I__7812 (
            .O(N__40170),
            .I(N__40167));
    Odrv4 I__7811 (
            .O(N__40167),
            .I(\serializer_mod_inst.shift_regZ0Z_66 ));
    InMux I__7810 (
            .O(N__40164),
            .I(N__40161));
    LocalMux I__7809 (
            .O(N__40161),
            .I(\serializer_mod_inst.shift_regZ0Z_102 ));
    CascadeMux I__7808 (
            .O(N__40158),
            .I(N__40155));
    InMux I__7807 (
            .O(N__40155),
            .I(N__40152));
    LocalMux I__7806 (
            .O(N__40152),
            .I(N__40149));
    Odrv4 I__7805 (
            .O(N__40149),
            .I(\serializer_mod_inst.shift_regZ0Z_103 ));
    InMux I__7804 (
            .O(N__40146),
            .I(N__40143));
    LocalMux I__7803 (
            .O(N__40143),
            .I(\serializer_mod_inst.shift_regZ0Z_84 ));
    InMux I__7802 (
            .O(N__40140),
            .I(N__40137));
    LocalMux I__7801 (
            .O(N__40137),
            .I(N__40134));
    Odrv12 I__7800 (
            .O(N__40134),
            .I(\serializer_mod_inst.shift_regZ0Z_41 ));
    InMux I__7799 (
            .O(N__40131),
            .I(N__40128));
    LocalMux I__7798 (
            .O(N__40128),
            .I(N__40125));
    Odrv4 I__7797 (
            .O(N__40125),
            .I(\serializer_mod_inst.shift_regZ0Z_100 ));
    InMux I__7796 (
            .O(N__40122),
            .I(N__40119));
    LocalMux I__7795 (
            .O(N__40119),
            .I(N__40116));
    Odrv4 I__7794 (
            .O(N__40116),
            .I(\serializer_mod_inst.shift_regZ0Z_54 ));
    InMux I__7793 (
            .O(N__40113),
            .I(N__40108));
    InMux I__7792 (
            .O(N__40112),
            .I(N__40105));
    InMux I__7791 (
            .O(N__40111),
            .I(N__40102));
    LocalMux I__7790 (
            .O(N__40108),
            .I(N__40099));
    LocalMux I__7789 (
            .O(N__40105),
            .I(N__40093));
    LocalMux I__7788 (
            .O(N__40102),
            .I(N__40090));
    Span4Mux_h I__7787 (
            .O(N__40099),
            .I(N__40087));
    InMux I__7786 (
            .O(N__40098),
            .I(N__40080));
    InMux I__7785 (
            .O(N__40097),
            .I(N__40080));
    InMux I__7784 (
            .O(N__40096),
            .I(N__40080));
    Span4Mux_v I__7783 (
            .O(N__40093),
            .I(N__40077));
    Span4Mux_v I__7782 (
            .O(N__40090),
            .I(N__40074));
    Span4Mux_v I__7781 (
            .O(N__40087),
            .I(N__40069));
    LocalMux I__7780 (
            .O(N__40080),
            .I(N__40069));
    Sp12to4 I__7779 (
            .O(N__40077),
            .I(N__40064));
    Sp12to4 I__7778 (
            .O(N__40074),
            .I(N__40064));
    Span4Mux_h I__7777 (
            .O(N__40069),
            .I(N__40061));
    Span12Mux_h I__7776 (
            .O(N__40064),
            .I(N__40056));
    Span4Mux_h I__7775 (
            .O(N__40061),
            .I(N__40053));
    InMux I__7774 (
            .O(N__40060),
            .I(N__40048));
    InMux I__7773 (
            .O(N__40059),
            .I(N__40048));
    Odrv12 I__7772 (
            .O(N__40056),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_0));
    Odrv4 I__7771 (
            .O(N__40053),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_0));
    LocalMux I__7770 (
            .O(N__40048),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_0));
    InMux I__7769 (
            .O(N__40041),
            .I(N__40038));
    LocalMux I__7768 (
            .O(N__40038),
            .I(N__40034));
    InMux I__7767 (
            .O(N__40037),
            .I(N__40030));
    Span4Mux_h I__7766 (
            .O(N__40034),
            .I(N__40027));
    InMux I__7765 (
            .O(N__40033),
            .I(N__40024));
    LocalMux I__7764 (
            .O(N__40030),
            .I(N__40021));
    Span4Mux_v I__7763 (
            .O(N__40027),
            .I(N__40018));
    LocalMux I__7762 (
            .O(N__40024),
            .I(N__40015));
    Span4Mux_h I__7761 (
            .O(N__40021),
            .I(N__40012));
    Span4Mux_v I__7760 (
            .O(N__40018),
            .I(N__40009));
    Odrv4 I__7759 (
            .O(N__40015),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0 ));
    Odrv4 I__7758 (
            .O(N__40012),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0 ));
    Odrv4 I__7757 (
            .O(N__40009),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0 ));
    InMux I__7756 (
            .O(N__40002),
            .I(N__39997));
    InMux I__7755 (
            .O(N__40001),
            .I(N__39994));
    InMux I__7754 (
            .O(N__40000),
            .I(N__39991));
    LocalMux I__7753 (
            .O(N__39997),
            .I(N__39988));
    LocalMux I__7752 (
            .O(N__39994),
            .I(N__39985));
    LocalMux I__7751 (
            .O(N__39991),
            .I(N__39982));
    Span4Mux_v I__7750 (
            .O(N__39988),
            .I(N__39979));
    Span4Mux_h I__7749 (
            .O(N__39985),
            .I(N__39976));
    Span12Mux_h I__7748 (
            .O(N__39982),
            .I(N__39971));
    Sp12to4 I__7747 (
            .O(N__39979),
            .I(N__39971));
    Odrv4 I__7746 (
            .O(N__39976),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6 ));
    Odrv12 I__7745 (
            .O(N__39971),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6 ));
    CascadeMux I__7744 (
            .O(N__39966),
            .I(N__39963));
    InMux I__7743 (
            .O(N__39963),
            .I(N__39960));
    LocalMux I__7742 (
            .O(N__39960),
            .I(\serializer_mod_inst.shift_regZ0Z_52 ));
    InMux I__7741 (
            .O(N__39957),
            .I(N__39954));
    LocalMux I__7740 (
            .O(N__39954),
            .I(\serializer_mod_inst.shift_regZ0Z_53 ));
    CascadeMux I__7739 (
            .O(N__39951),
            .I(N__39948));
    InMux I__7738 (
            .O(N__39948),
            .I(N__39945));
    LocalMux I__7737 (
            .O(N__39945),
            .I(\serializer_mod_inst.shift_regZ0Z_87 ));
    InMux I__7736 (
            .O(N__39942),
            .I(N__39939));
    LocalMux I__7735 (
            .O(N__39939),
            .I(\serializer_mod_inst.shift_regZ0Z_88 ));
    InMux I__7734 (
            .O(N__39936),
            .I(N__39933));
    LocalMux I__7733 (
            .O(N__39933),
            .I(\serializer_mod_inst.shift_regZ0Z_49 ));
    CascadeMux I__7732 (
            .O(N__39930),
            .I(N__39927));
    InMux I__7731 (
            .O(N__39927),
            .I(N__39924));
    LocalMux I__7730 (
            .O(N__39924),
            .I(\serializer_mod_inst.shift_regZ0Z_50 ));
    InMux I__7729 (
            .O(N__39921),
            .I(N__39918));
    LocalMux I__7728 (
            .O(N__39918),
            .I(\serializer_mod_inst.shift_regZ0Z_89 ));
    InMux I__7727 (
            .O(N__39915),
            .I(N__39912));
    LocalMux I__7726 (
            .O(N__39912),
            .I(\serializer_mod_inst.shift_regZ0Z_90 ));
    InMux I__7725 (
            .O(N__39909),
            .I(N__39905));
    InMux I__7724 (
            .O(N__39908),
            .I(N__39902));
    LocalMux I__7723 (
            .O(N__39905),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_9));
    LocalMux I__7722 (
            .O(N__39902),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_9));
    InMux I__7721 (
            .O(N__39897),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8 ));
    InMux I__7720 (
            .O(N__39894),
            .I(N__39890));
    InMux I__7719 (
            .O(N__39893),
            .I(N__39887));
    LocalMux I__7718 (
            .O(N__39890),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_10));
    LocalMux I__7717 (
            .O(N__39887),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_10));
    InMux I__7716 (
            .O(N__39882),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9 ));
    InMux I__7715 (
            .O(N__39879),
            .I(N__39875));
    InMux I__7714 (
            .O(N__39878),
            .I(N__39872));
    LocalMux I__7713 (
            .O(N__39875),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_11));
    LocalMux I__7712 (
            .O(N__39872),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_11));
    InMux I__7711 (
            .O(N__39867),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10 ));
    InMux I__7710 (
            .O(N__39864),
            .I(N__39860));
    InMux I__7709 (
            .O(N__39863),
            .I(N__39857));
    LocalMux I__7708 (
            .O(N__39860),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_12));
    LocalMux I__7707 (
            .O(N__39857),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_12));
    InMux I__7706 (
            .O(N__39852),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11 ));
    InMux I__7705 (
            .O(N__39849),
            .I(N__39845));
    InMux I__7704 (
            .O(N__39848),
            .I(N__39842));
    LocalMux I__7703 (
            .O(N__39845),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_13));
    LocalMux I__7702 (
            .O(N__39842),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_13));
    InMux I__7701 (
            .O(N__39837),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12 ));
    CascadeMux I__7700 (
            .O(N__39834),
            .I(N__39830));
    InMux I__7699 (
            .O(N__39833),
            .I(N__39827));
    InMux I__7698 (
            .O(N__39830),
            .I(N__39824));
    LocalMux I__7697 (
            .O(N__39827),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_14));
    LocalMux I__7696 (
            .O(N__39824),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_14));
    InMux I__7695 (
            .O(N__39819),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13 ));
    InMux I__7694 (
            .O(N__39816),
            .I(N__39800));
    InMux I__7693 (
            .O(N__39815),
            .I(N__39800));
    InMux I__7692 (
            .O(N__39814),
            .I(N__39800));
    InMux I__7691 (
            .O(N__39813),
            .I(N__39800));
    InMux I__7690 (
            .O(N__39812),
            .I(N__39782));
    InMux I__7689 (
            .O(N__39811),
            .I(N__39782));
    InMux I__7688 (
            .O(N__39810),
            .I(N__39782));
    InMux I__7687 (
            .O(N__39809),
            .I(N__39782));
    LocalMux I__7686 (
            .O(N__39800),
            .I(N__39779));
    InMux I__7685 (
            .O(N__39799),
            .I(N__39770));
    InMux I__7684 (
            .O(N__39798),
            .I(N__39770));
    InMux I__7683 (
            .O(N__39797),
            .I(N__39770));
    InMux I__7682 (
            .O(N__39796),
            .I(N__39770));
    InMux I__7681 (
            .O(N__39795),
            .I(N__39761));
    InMux I__7680 (
            .O(N__39794),
            .I(N__39761));
    InMux I__7679 (
            .O(N__39793),
            .I(N__39761));
    InMux I__7678 (
            .O(N__39792),
            .I(N__39761));
    InMux I__7677 (
            .O(N__39791),
            .I(N__39758));
    LocalMux I__7676 (
            .O(N__39782),
            .I(N__39754));
    Span4Mux_v I__7675 (
            .O(N__39779),
            .I(N__39747));
    LocalMux I__7674 (
            .O(N__39770),
            .I(N__39747));
    LocalMux I__7673 (
            .O(N__39761),
            .I(N__39747));
    LocalMux I__7672 (
            .O(N__39758),
            .I(N__39744));
    InMux I__7671 (
            .O(N__39757),
            .I(N__39739));
    Span4Mux_h I__7670 (
            .O(N__39754),
            .I(N__39736));
    Span4Mux_h I__7669 (
            .O(N__39747),
            .I(N__39733));
    Span12Mux_v I__7668 (
            .O(N__39744),
            .I(N__39730));
    InMux I__7667 (
            .O(N__39743),
            .I(N__39725));
    InMux I__7666 (
            .O(N__39742),
            .I(N__39725));
    LocalMux I__7665 (
            .O(N__39739),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ));
    Odrv4 I__7664 (
            .O(N__39736),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ));
    Odrv4 I__7663 (
            .O(N__39733),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ));
    Odrv12 I__7662 (
            .O(N__39730),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ));
    LocalMux I__7661 (
            .O(N__39725),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ));
    InMux I__7660 (
            .O(N__39714),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_14 ));
    CascadeMux I__7659 (
            .O(N__39711),
            .I(N__39707));
    InMux I__7658 (
            .O(N__39710),
            .I(N__39704));
    InMux I__7657 (
            .O(N__39707),
            .I(N__39701));
    LocalMux I__7656 (
            .O(N__39704),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_15));
    LocalMux I__7655 (
            .O(N__39701),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_15));
    CEMux I__7654 (
            .O(N__39696),
            .I(N__39692));
    CEMux I__7653 (
            .O(N__39695),
            .I(N__39689));
    LocalMux I__7652 (
            .O(N__39692),
            .I(N__39686));
    LocalMux I__7651 (
            .O(N__39689),
            .I(N__39683));
    Span4Mux_h I__7650 (
            .O(N__39686),
            .I(N__39680));
    Span4Mux_h I__7649 (
            .O(N__39683),
            .I(N__39677));
    Span4Mux_h I__7648 (
            .O(N__39680),
            .I(N__39674));
    Span4Mux_h I__7647 (
            .O(N__39677),
            .I(N__39671));
    Odrv4 I__7646 (
            .O(N__39674),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0 ));
    Odrv4 I__7645 (
            .O(N__39671),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0 ));
    InMux I__7644 (
            .O(N__39666),
            .I(N__39663));
    LocalMux I__7643 (
            .O(N__39663),
            .I(\serializer_mod_inst.shift_regZ0Z_86 ));
    CascadeMux I__7642 (
            .O(N__39660),
            .I(N__39657));
    InMux I__7641 (
            .O(N__39657),
            .I(N__39654));
    LocalMux I__7640 (
            .O(N__39654),
            .I(N__39650));
    InMux I__7639 (
            .O(N__39653),
            .I(N__39647));
    Span4Mux_h I__7638 (
            .O(N__39650),
            .I(N__39643));
    LocalMux I__7637 (
            .O(N__39647),
            .I(N__39640));
    InMux I__7636 (
            .O(N__39646),
            .I(N__39637));
    Span4Mux_v I__7635 (
            .O(N__39643),
            .I(N__39634));
    Span12Mux_v I__7634 (
            .O(N__39640),
            .I(N__39631));
    LocalMux I__7633 (
            .O(N__39637),
            .I(\cemf_module_64ch_ctrl_inst1.paddr_fsm_1 ));
    Odrv4 I__7632 (
            .O(N__39634),
            .I(\cemf_module_64ch_ctrl_inst1.paddr_fsm_1 ));
    Odrv12 I__7631 (
            .O(N__39631),
            .I(\cemf_module_64ch_ctrl_inst1.paddr_fsm_1 ));
    InMux I__7630 (
            .O(N__39624),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0 ));
    InMux I__7629 (
            .O(N__39621),
            .I(N__39618));
    LocalMux I__7628 (
            .O(N__39618),
            .I(N__39614));
    CascadeMux I__7627 (
            .O(N__39617),
            .I(N__39608));
    Span4Mux_h I__7626 (
            .O(N__39614),
            .I(N__39605));
    InMux I__7625 (
            .O(N__39613),
            .I(N__39596));
    InMux I__7624 (
            .O(N__39612),
            .I(N__39596));
    InMux I__7623 (
            .O(N__39611),
            .I(N__39596));
    InMux I__7622 (
            .O(N__39608),
            .I(N__39596));
    Span4Mux_h I__7621 (
            .O(N__39605),
            .I(N__39590));
    LocalMux I__7620 (
            .O(N__39596),
            .I(N__39590));
    InMux I__7619 (
            .O(N__39595),
            .I(N__39587));
    Span4Mux_h I__7618 (
            .O(N__39590),
            .I(N__39584));
    LocalMux I__7617 (
            .O(N__39587),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_2));
    Odrv4 I__7616 (
            .O(N__39584),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_2));
    InMux I__7615 (
            .O(N__39579),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1 ));
    InMux I__7614 (
            .O(N__39576),
            .I(N__39573));
    LocalMux I__7613 (
            .O(N__39573),
            .I(N__39570));
    Span4Mux_h I__7612 (
            .O(N__39570),
            .I(N__39567));
    Span4Mux_h I__7611 (
            .O(N__39567),
            .I(N__39561));
    InMux I__7610 (
            .O(N__39566),
            .I(N__39558));
    InMux I__7609 (
            .O(N__39565),
            .I(N__39555));
    InMux I__7608 (
            .O(N__39564),
            .I(N__39552));
    Span4Mux_h I__7607 (
            .O(N__39561),
            .I(N__39547));
    LocalMux I__7606 (
            .O(N__39558),
            .I(N__39547));
    LocalMux I__7605 (
            .O(N__39555),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_3));
    LocalMux I__7604 (
            .O(N__39552),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_3));
    Odrv4 I__7603 (
            .O(N__39547),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_3));
    InMux I__7602 (
            .O(N__39540),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2 ));
    InMux I__7601 (
            .O(N__39537),
            .I(N__39532));
    InMux I__7600 (
            .O(N__39536),
            .I(N__39529));
    InMux I__7599 (
            .O(N__39535),
            .I(N__39526));
    LocalMux I__7598 (
            .O(N__39532),
            .I(N__39521));
    LocalMux I__7597 (
            .O(N__39529),
            .I(N__39521));
    LocalMux I__7596 (
            .O(N__39526),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_4));
    Odrv4 I__7595 (
            .O(N__39521),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_4));
    InMux I__7594 (
            .O(N__39516),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3 ));
    InMux I__7593 (
            .O(N__39513),
            .I(N__39509));
    InMux I__7592 (
            .O(N__39512),
            .I(N__39506));
    LocalMux I__7591 (
            .O(N__39509),
            .I(N__39500));
    LocalMux I__7590 (
            .O(N__39506),
            .I(N__39500));
    InMux I__7589 (
            .O(N__39505),
            .I(N__39497));
    Span4Mux_v I__7588 (
            .O(N__39500),
            .I(N__39494));
    LocalMux I__7587 (
            .O(N__39497),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_5));
    Odrv4 I__7586 (
            .O(N__39494),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_5));
    InMux I__7585 (
            .O(N__39489),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4 ));
    CascadeMux I__7584 (
            .O(N__39486),
            .I(N__39482));
    InMux I__7583 (
            .O(N__39485),
            .I(N__39479));
    InMux I__7582 (
            .O(N__39482),
            .I(N__39476));
    LocalMux I__7581 (
            .O(N__39479),
            .I(N__39470));
    LocalMux I__7580 (
            .O(N__39476),
            .I(N__39470));
    InMux I__7579 (
            .O(N__39475),
            .I(N__39467));
    Span4Mux_h I__7578 (
            .O(N__39470),
            .I(N__39464));
    LocalMux I__7577 (
            .O(N__39467),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_6));
    Odrv4 I__7576 (
            .O(N__39464),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_6));
    InMux I__7575 (
            .O(N__39459),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5 ));
    InMux I__7574 (
            .O(N__39456),
            .I(N__39452));
    InMux I__7573 (
            .O(N__39455),
            .I(N__39449));
    LocalMux I__7572 (
            .O(N__39452),
            .I(N__39445));
    LocalMux I__7571 (
            .O(N__39449),
            .I(N__39442));
    InMux I__7570 (
            .O(N__39448),
            .I(N__39439));
    Span4Mux_h I__7569 (
            .O(N__39445),
            .I(N__39434));
    Span4Mux_h I__7568 (
            .O(N__39442),
            .I(N__39434));
    LocalMux I__7567 (
            .O(N__39439),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7 ));
    Odrv4 I__7566 (
            .O(N__39434),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7 ));
    InMux I__7565 (
            .O(N__39429),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6 ));
    InMux I__7564 (
            .O(N__39426),
            .I(N__39422));
    InMux I__7563 (
            .O(N__39425),
            .I(N__39418));
    LocalMux I__7562 (
            .O(N__39422),
            .I(N__39415));
    InMux I__7561 (
            .O(N__39421),
            .I(N__39412));
    LocalMux I__7560 (
            .O(N__39418),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_8));
    Odrv4 I__7559 (
            .O(N__39415),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_8));
    LocalMux I__7558 (
            .O(N__39412),
            .I(cemf_module_64ch_ctrl_inst1_paddr_fsm_8));
    InMux I__7557 (
            .O(N__39405),
            .I(bfn_18_21_0_));
    SRMux I__7556 (
            .O(N__39402),
            .I(N__39397));
    SRMux I__7555 (
            .O(N__39401),
            .I(N__39393));
    SRMux I__7554 (
            .O(N__39400),
            .I(N__39389));
    LocalMux I__7553 (
            .O(N__39397),
            .I(N__39386));
    SRMux I__7552 (
            .O(N__39396),
            .I(N__39383));
    LocalMux I__7551 (
            .O(N__39393),
            .I(N__39378));
    SRMux I__7550 (
            .O(N__39392),
            .I(N__39375));
    LocalMux I__7549 (
            .O(N__39389),
            .I(N__39366));
    Span4Mux_s0_v I__7548 (
            .O(N__39386),
            .I(N__39366));
    LocalMux I__7547 (
            .O(N__39383),
            .I(N__39366));
    SRMux I__7546 (
            .O(N__39382),
            .I(N__39363));
    SRMux I__7545 (
            .O(N__39381),
            .I(N__39359));
    Span4Mux_v I__7544 (
            .O(N__39378),
            .I(N__39354));
    LocalMux I__7543 (
            .O(N__39375),
            .I(N__39354));
    SRMux I__7542 (
            .O(N__39374),
            .I(N__39351));
    SRMux I__7541 (
            .O(N__39373),
            .I(N__39347));
    Span4Mux_v I__7540 (
            .O(N__39366),
            .I(N__39340));
    LocalMux I__7539 (
            .O(N__39363),
            .I(N__39340));
    SRMux I__7538 (
            .O(N__39362),
            .I(N__39337));
    LocalMux I__7537 (
            .O(N__39359),
            .I(N__39329));
    Span4Mux_h I__7536 (
            .O(N__39354),
            .I(N__39329));
    LocalMux I__7535 (
            .O(N__39351),
            .I(N__39329));
    SRMux I__7534 (
            .O(N__39350),
            .I(N__39326));
    LocalMux I__7533 (
            .O(N__39347),
            .I(N__39322));
    CascadeMux I__7532 (
            .O(N__39346),
            .I(N__39319));
    CascadeMux I__7531 (
            .O(N__39345),
            .I(N__39316));
    Span4Mux_v I__7530 (
            .O(N__39340),
            .I(N__39309));
    LocalMux I__7529 (
            .O(N__39337),
            .I(N__39309));
    SRMux I__7528 (
            .O(N__39336),
            .I(N__39306));
    Span4Mux_v I__7527 (
            .O(N__39329),
            .I(N__39300));
    LocalMux I__7526 (
            .O(N__39326),
            .I(N__39300));
    SRMux I__7525 (
            .O(N__39325),
            .I(N__39297));
    Span4Mux_h I__7524 (
            .O(N__39322),
            .I(N__39293));
    InMux I__7523 (
            .O(N__39319),
            .I(N__39290));
    InMux I__7522 (
            .O(N__39316),
            .I(N__39287));
    CascadeMux I__7521 (
            .O(N__39315),
            .I(N__39283));
    SRMux I__7520 (
            .O(N__39314),
            .I(N__39278));
    Span4Mux_h I__7519 (
            .O(N__39309),
            .I(N__39273));
    LocalMux I__7518 (
            .O(N__39306),
            .I(N__39273));
    SRMux I__7517 (
            .O(N__39305),
            .I(N__39270));
    Span4Mux_v I__7516 (
            .O(N__39300),
            .I(N__39265));
    LocalMux I__7515 (
            .O(N__39297),
            .I(N__39265));
    SRMux I__7514 (
            .O(N__39296),
            .I(N__39262));
    Span4Mux_v I__7513 (
            .O(N__39293),
            .I(N__39259));
    LocalMux I__7512 (
            .O(N__39290),
            .I(N__39254));
    LocalMux I__7511 (
            .O(N__39287),
            .I(N__39254));
    InMux I__7510 (
            .O(N__39286),
            .I(N__39244));
    InMux I__7509 (
            .O(N__39283),
            .I(N__39244));
    InMux I__7508 (
            .O(N__39282),
            .I(N__39244));
    InMux I__7507 (
            .O(N__39281),
            .I(N__39244));
    LocalMux I__7506 (
            .O(N__39278),
            .I(N__39241));
    Span4Mux_v I__7505 (
            .O(N__39273),
            .I(N__39236));
    LocalMux I__7504 (
            .O(N__39270),
            .I(N__39236));
    Span4Mux_h I__7503 (
            .O(N__39265),
            .I(N__39231));
    LocalMux I__7502 (
            .O(N__39262),
            .I(N__39231));
    Span4Mux_v I__7501 (
            .O(N__39259),
            .I(N__39226));
    Span4Mux_h I__7500 (
            .O(N__39254),
            .I(N__39226));
    InMux I__7499 (
            .O(N__39253),
            .I(N__39223));
    LocalMux I__7498 (
            .O(N__39244),
            .I(N__39220));
    Span4Mux_v I__7497 (
            .O(N__39241),
            .I(N__39217));
    Span4Mux_v I__7496 (
            .O(N__39236),
            .I(N__39212));
    Span4Mux_v I__7495 (
            .O(N__39231),
            .I(N__39212));
    Span4Mux_h I__7494 (
            .O(N__39226),
            .I(N__39207));
    LocalMux I__7493 (
            .O(N__39223),
            .I(N__39207));
    Span4Mux_v I__7492 (
            .O(N__39220),
            .I(N__39204));
    Span4Mux_h I__7491 (
            .O(N__39217),
            .I(N__39199));
    Span4Mux_h I__7490 (
            .O(N__39212),
            .I(N__39199));
    Span4Mux_h I__7489 (
            .O(N__39207),
            .I(N__39196));
    Sp12to4 I__7488 (
            .O(N__39204),
            .I(N__39193));
    Odrv4 I__7487 (
            .O(N__39199),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__7486 (
            .O(N__39196),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__7485 (
            .O(N__39193),
            .I(CONSTANT_ONE_NET));
    InMux I__7484 (
            .O(N__39186),
            .I(N__39183));
    LocalMux I__7483 (
            .O(N__39183),
            .I(N__39180));
    Span4Mux_v I__7482 (
            .O(N__39180),
            .I(N__39177));
    Odrv4 I__7481 (
            .O(N__39177),
            .I(\I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rstZ0 ));
    SRMux I__7480 (
            .O(N__39174),
            .I(N__39171));
    LocalMux I__7479 (
            .O(N__39171),
            .I(N__39168));
    Span4Mux_v I__7478 (
            .O(N__39168),
            .I(N__39165));
    Span4Mux_h I__7477 (
            .O(N__39165),
            .I(N__39162));
    Span4Mux_h I__7476 (
            .O(N__39162),
            .I(N__39159));
    Span4Mux_v I__7475 (
            .O(N__39159),
            .I(N__39156));
    Odrv4 I__7474 (
            .O(N__39156),
            .I(\I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNOZ0 ));
    CascadeMux I__7473 (
            .O(N__39153),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa_cascade_ ));
    CascadeMux I__7472 (
            .O(N__39150),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_3_cascade_ ));
    CascadeMux I__7471 (
            .O(N__39147),
            .I(N__39137));
    InMux I__7470 (
            .O(N__39146),
            .I(N__39134));
    InMux I__7469 (
            .O(N__39145),
            .I(N__39125));
    InMux I__7468 (
            .O(N__39144),
            .I(N__39125));
    InMux I__7467 (
            .O(N__39143),
            .I(N__39125));
    InMux I__7466 (
            .O(N__39142),
            .I(N__39120));
    InMux I__7465 (
            .O(N__39141),
            .I(N__39120));
    InMux I__7464 (
            .O(N__39140),
            .I(N__39117));
    InMux I__7463 (
            .O(N__39137),
            .I(N__39110));
    LocalMux I__7462 (
            .O(N__39134),
            .I(N__39102));
    InMux I__7461 (
            .O(N__39133),
            .I(N__39099));
    InMux I__7460 (
            .O(N__39132),
            .I(N__39096));
    LocalMux I__7459 (
            .O(N__39125),
            .I(N__39093));
    LocalMux I__7458 (
            .O(N__39120),
            .I(N__39088));
    LocalMux I__7457 (
            .O(N__39117),
            .I(N__39088));
    InMux I__7456 (
            .O(N__39116),
            .I(N__39079));
    InMux I__7455 (
            .O(N__39115),
            .I(N__39079));
    InMux I__7454 (
            .O(N__39114),
            .I(N__39079));
    InMux I__7453 (
            .O(N__39113),
            .I(N__39079));
    LocalMux I__7452 (
            .O(N__39110),
            .I(N__39076));
    InMux I__7451 (
            .O(N__39109),
            .I(N__39073));
    InMux I__7450 (
            .O(N__39108),
            .I(N__39064));
    InMux I__7449 (
            .O(N__39107),
            .I(N__39064));
    InMux I__7448 (
            .O(N__39106),
            .I(N__39064));
    InMux I__7447 (
            .O(N__39105),
            .I(N__39064));
    Span4Mux_v I__7446 (
            .O(N__39102),
            .I(N__39059));
    LocalMux I__7445 (
            .O(N__39099),
            .I(N__39059));
    LocalMux I__7444 (
            .O(N__39096),
            .I(N_1975));
    Odrv4 I__7443 (
            .O(N__39093),
            .I(N_1975));
    Odrv12 I__7442 (
            .O(N__39088),
            .I(N_1975));
    LocalMux I__7441 (
            .O(N__39079),
            .I(N_1975));
    Odrv12 I__7440 (
            .O(N__39076),
            .I(N_1975));
    LocalMux I__7439 (
            .O(N__39073),
            .I(N_1975));
    LocalMux I__7438 (
            .O(N__39064),
            .I(N_1975));
    Odrv4 I__7437 (
            .O(N__39059),
            .I(N_1975));
    InMux I__7436 (
            .O(N__39042),
            .I(N__39039));
    LocalMux I__7435 (
            .O(N__39039),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNOZ0 ));
    InMux I__7434 (
            .O(N__39036),
            .I(N__39033));
    LocalMux I__7433 (
            .O(N__39033),
            .I(N__39029));
    InMux I__7432 (
            .O(N__39032),
            .I(N__39026));
    Span4Mux_h I__7431 (
            .O(N__39029),
            .I(N__39023));
    LocalMux I__7430 (
            .O(N__39026),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0 ));
    Odrv4 I__7429 (
            .O(N__39023),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0 ));
    InMux I__7428 (
            .O(N__39018),
            .I(bfn_18_20_0_));
    InMux I__7427 (
            .O(N__39015),
            .I(N__39012));
    LocalMux I__7426 (
            .O(N__39012),
            .I(N__39008));
    CascadeMux I__7425 (
            .O(N__39011),
            .I(N__39005));
    Span12Mux_v I__7424 (
            .O(N__39008),
            .I(N__39002));
    InMux I__7423 (
            .O(N__39005),
            .I(N__38999));
    Odrv12 I__7422 (
            .O(N__39002),
            .I(\cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4 ));
    LocalMux I__7421 (
            .O(N__38999),
            .I(\cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4 ));
    InMux I__7420 (
            .O(N__38994),
            .I(N__38991));
    LocalMux I__7419 (
            .O(N__38991),
            .I(N__38988));
    Span4Mux_h I__7418 (
            .O(N__38988),
            .I(N__38985));
    Span4Mux_v I__7417 (
            .O(N__38985),
            .I(N__38982));
    Span4Mux_h I__7416 (
            .O(N__38982),
            .I(N__38979));
    Odrv4 I__7415 (
            .O(N__38979),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_CO ));
    InMux I__7414 (
            .O(N__38976),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0 ));
    InMux I__7413 (
            .O(N__38973),
            .I(N__38970));
    LocalMux I__7412 (
            .O(N__38970),
            .I(N__38967));
    Span4Mux_h I__7411 (
            .O(N__38967),
            .I(N__38964));
    Span4Mux_h I__7410 (
            .O(N__38964),
            .I(N__38961));
    Span4Mux_h I__7409 (
            .O(N__38961),
            .I(N__38957));
    InMux I__7408 (
            .O(N__38960),
            .I(N__38954));
    Odrv4 I__7407 (
            .O(N__38957),
            .I(\cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5 ));
    LocalMux I__7406 (
            .O(N__38954),
            .I(\cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5 ));
    InMux I__7405 (
            .O(N__38949),
            .I(N__38946));
    LocalMux I__7404 (
            .O(N__38946),
            .I(N__38943));
    Span4Mux_h I__7403 (
            .O(N__38943),
            .I(N__38940));
    Span4Mux_h I__7402 (
            .O(N__38940),
            .I(N__38937));
    Span4Mux_h I__7401 (
            .O(N__38937),
            .I(N__38934));
    Odrv4 I__7400 (
            .O(N__38934),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_CO ));
    InMux I__7399 (
            .O(N__38931),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1 ));
    CascadeMux I__7398 (
            .O(N__38928),
            .I(N__38925));
    InMux I__7397 (
            .O(N__38925),
            .I(N__38922));
    LocalMux I__7396 (
            .O(N__38922),
            .I(\cemf_module_64ch_ctrl_inst1.c_addr_RNI3UAS1_6 ));
    InMux I__7395 (
            .O(N__38919),
            .I(N__38916));
    LocalMux I__7394 (
            .O(N__38916),
            .I(N__38913));
    Span4Mux_s1_v I__7393 (
            .O(N__38913),
            .I(N__38909));
    InMux I__7392 (
            .O(N__38912),
            .I(N__38906));
    Span4Mux_v I__7391 (
            .O(N__38909),
            .I(N__38900));
    LocalMux I__7390 (
            .O(N__38906),
            .I(N__38897));
    InMux I__7389 (
            .O(N__38905),
            .I(N__38894));
    InMux I__7388 (
            .O(N__38904),
            .I(N__38886));
    InMux I__7387 (
            .O(N__38903),
            .I(N__38886));
    Span4Mux_v I__7386 (
            .O(N__38900),
            .I(N__38881));
    Span4Mux_h I__7385 (
            .O(N__38897),
            .I(N__38881));
    LocalMux I__7384 (
            .O(N__38894),
            .I(N__38878));
    InMux I__7383 (
            .O(N__38893),
            .I(N__38873));
    InMux I__7382 (
            .O(N__38892),
            .I(N__38873));
    InMux I__7381 (
            .O(N__38891),
            .I(N__38870));
    LocalMux I__7380 (
            .O(N__38886),
            .I(N__38867));
    Span4Mux_v I__7379 (
            .O(N__38881),
            .I(N__38862));
    Span4Mux_h I__7378 (
            .O(N__38878),
            .I(N__38862));
    LocalMux I__7377 (
            .O(N__38873),
            .I(N__38859));
    LocalMux I__7376 (
            .O(N__38870),
            .I(N__38856));
    Span4Mux_v I__7375 (
            .O(N__38867),
            .I(N__38851));
    Span4Mux_h I__7374 (
            .O(N__38862),
            .I(N__38851));
    Span4Mux_h I__7373 (
            .O(N__38859),
            .I(N__38848));
    Span12Mux_h I__7372 (
            .O(N__38856),
            .I(N__38845));
    Span4Mux_h I__7371 (
            .O(N__38851),
            .I(N__38842));
    Odrv4 I__7370 (
            .O(N__38848),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1 ));
    Odrv12 I__7369 (
            .O(N__38845),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1 ));
    Odrv4 I__7368 (
            .O(N__38842),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1 ));
    InMux I__7367 (
            .O(N__38835),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2 ));
    CascadeMux I__7366 (
            .O(N__38832),
            .I(N__38829));
    InMux I__7365 (
            .O(N__38829),
            .I(N__38826));
    LocalMux I__7364 (
            .O(N__38826),
            .I(\cemf_module_64ch_ctrl_inst1.c_addr_RNI50BS1_7 ));
    InMux I__7363 (
            .O(N__38823),
            .I(N__38817));
    InMux I__7362 (
            .O(N__38822),
            .I(N__38814));
    InMux I__7361 (
            .O(N__38821),
            .I(N__38809));
    InMux I__7360 (
            .O(N__38820),
            .I(N__38809));
    LocalMux I__7359 (
            .O(N__38817),
            .I(N__38803));
    LocalMux I__7358 (
            .O(N__38814),
            .I(N__38799));
    LocalMux I__7357 (
            .O(N__38809),
            .I(N__38796));
    InMux I__7356 (
            .O(N__38808),
            .I(N__38791));
    InMux I__7355 (
            .O(N__38807),
            .I(N__38791));
    InMux I__7354 (
            .O(N__38806),
            .I(N__38788));
    Sp12to4 I__7353 (
            .O(N__38803),
            .I(N__38785));
    InMux I__7352 (
            .O(N__38802),
            .I(N__38782));
    Span4Mux_h I__7351 (
            .O(N__38799),
            .I(N__38779));
    Span4Mux_v I__7350 (
            .O(N__38796),
            .I(N__38774));
    LocalMux I__7349 (
            .O(N__38791),
            .I(N__38774));
    LocalMux I__7348 (
            .O(N__38788),
            .I(N__38771));
    Span12Mux_s5_v I__7347 (
            .O(N__38785),
            .I(N__38766));
    LocalMux I__7346 (
            .O(N__38782),
            .I(N__38766));
    Span4Mux_h I__7345 (
            .O(N__38779),
            .I(N__38763));
    Span4Mux_h I__7344 (
            .O(N__38774),
            .I(N__38760));
    Span12Mux_h I__7343 (
            .O(N__38771),
            .I(N__38757));
    Span12Mux_v I__7342 (
            .O(N__38766),
            .I(N__38754));
    Span4Mux_h I__7341 (
            .O(N__38763),
            .I(N__38751));
    Odrv4 I__7340 (
            .O(N__38760),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1 ));
    Odrv12 I__7339 (
            .O(N__38757),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1 ));
    Odrv12 I__7338 (
            .O(N__38754),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1 ));
    Odrv4 I__7337 (
            .O(N__38751),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1 ));
    InMux I__7336 (
            .O(N__38742),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3 ));
    InMux I__7335 (
            .O(N__38739),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4 ));
    InMux I__7334 (
            .O(N__38736),
            .I(N__38733));
    LocalMux I__7333 (
            .O(N__38733),
            .I(N__38730));
    Span4Mux_h I__7332 (
            .O(N__38730),
            .I(N__38727));
    Span4Mux_v I__7331 (
            .O(N__38727),
            .I(N__38723));
    InMux I__7330 (
            .O(N__38726),
            .I(N__38720));
    Span4Mux_v I__7329 (
            .O(N__38723),
            .I(N__38715));
    LocalMux I__7328 (
            .O(N__38720),
            .I(N__38715));
    Span4Mux_h I__7327 (
            .O(N__38715),
            .I(N__38712));
    Odrv4 I__7326 (
            .O(N__38712),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93STZ0Z1 ));
    CascadeMux I__7325 (
            .O(N__38709),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_8_0_m2_ns_1_cascade_ ));
    InMux I__7324 (
            .O(N__38706),
            .I(N__38703));
    LocalMux I__7323 (
            .O(N__38703),
            .I(N__38700));
    Span4Mux_v I__7322 (
            .O(N__38700),
            .I(N__38696));
    InMux I__7321 (
            .O(N__38699),
            .I(N__38693));
    Span4Mux_h I__7320 (
            .O(N__38696),
            .I(N__38690));
    LocalMux I__7319 (
            .O(N__38693),
            .I(N__38687));
    Odrv4 I__7318 (
            .O(N__38690),
            .I(N_1842_0));
    Odrv12 I__7317 (
            .O(N__38687),
            .I(N_1842_0));
    CascadeMux I__7316 (
            .O(N__38682),
            .I(N_1842_0_cascade_));
    InMux I__7315 (
            .O(N__38679),
            .I(N__38676));
    LocalMux I__7314 (
            .O(N__38676),
            .I(N__38670));
    InMux I__7313 (
            .O(N__38675),
            .I(N__38667));
    InMux I__7312 (
            .O(N__38674),
            .I(N__38661));
    InMux I__7311 (
            .O(N__38673),
            .I(N__38658));
    Span12Mux_h I__7310 (
            .O(N__38670),
            .I(N__38653));
    LocalMux I__7309 (
            .O(N__38667),
            .I(N__38650));
    InMux I__7308 (
            .O(N__38666),
            .I(N__38643));
    InMux I__7307 (
            .O(N__38665),
            .I(N__38643));
    InMux I__7306 (
            .O(N__38664),
            .I(N__38643));
    LocalMux I__7305 (
            .O(N__38661),
            .I(N__38638));
    LocalMux I__7304 (
            .O(N__38658),
            .I(N__38638));
    InMux I__7303 (
            .O(N__38657),
            .I(N__38634));
    InMux I__7302 (
            .O(N__38656),
            .I(N__38631));
    Span12Mux_v I__7301 (
            .O(N__38653),
            .I(N__38626));
    Span12Mux_v I__7300 (
            .O(N__38650),
            .I(N__38626));
    LocalMux I__7299 (
            .O(N__38643),
            .I(N__38621));
    Span4Mux_v I__7298 (
            .O(N__38638),
            .I(N__38621));
    InMux I__7297 (
            .O(N__38637),
            .I(N__38618));
    LocalMux I__7296 (
            .O(N__38634),
            .I(N_1841_0));
    LocalMux I__7295 (
            .O(N__38631),
            .I(N_1841_0));
    Odrv12 I__7294 (
            .O(N__38626),
            .I(N_1841_0));
    Odrv4 I__7293 (
            .O(N__38621),
            .I(N_1841_0));
    LocalMux I__7292 (
            .O(N__38618),
            .I(N_1841_0));
    InMux I__7291 (
            .O(N__38607),
            .I(N__38604));
    LocalMux I__7290 (
            .O(N__38604),
            .I(N__38601));
    Span4Mux_v I__7289 (
            .O(N__38601),
            .I(N__38598));
    Span4Mux_h I__7288 (
            .O(N__38598),
            .I(N__38593));
    InMux I__7287 (
            .O(N__38597),
            .I(N__38588));
    InMux I__7286 (
            .O(N__38596),
            .I(N__38588));
    Odrv4 I__7285 (
            .O(N__38593),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_22));
    LocalMux I__7284 (
            .O(N__38588),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_22));
    InMux I__7283 (
            .O(N__38583),
            .I(N__38580));
    LocalMux I__7282 (
            .O(N__38580),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_22 ));
    CascadeMux I__7281 (
            .O(N__38577),
            .I(N__38573));
    InMux I__7280 (
            .O(N__38576),
            .I(N__38570));
    InMux I__7279 (
            .O(N__38573),
            .I(N__38567));
    LocalMux I__7278 (
            .O(N__38570),
            .I(N__38561));
    LocalMux I__7277 (
            .O(N__38567),
            .I(N__38561));
    InMux I__7276 (
            .O(N__38566),
            .I(N__38558));
    Span4Mux_h I__7275 (
            .O(N__38561),
            .I(N__38555));
    LocalMux I__7274 (
            .O(N__38558),
            .I(cemf_module_64ch_ctrl_inst1_data_config_20));
    Odrv4 I__7273 (
            .O(N__38555),
            .I(cemf_module_64ch_ctrl_inst1_data_config_20));
    InMux I__7272 (
            .O(N__38550),
            .I(N__38547));
    LocalMux I__7271 (
            .O(N__38547),
            .I(N__38544));
    Span4Mux_v I__7270 (
            .O(N__38544),
            .I(N__38541));
    Span4Mux_v I__7269 (
            .O(N__38541),
            .I(N__38538));
    Sp12to4 I__7268 (
            .O(N__38538),
            .I(N__38535));
    Odrv12 I__7267 (
            .O(N__38535),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_30));
    InMux I__7266 (
            .O(N__38532),
            .I(N__38529));
    LocalMux I__7265 (
            .O(N__38529),
            .I(N__38526));
    Span4Mux_h I__7264 (
            .O(N__38526),
            .I(N__38523));
    Span4Mux_v I__7263 (
            .O(N__38523),
            .I(N__38520));
    Span4Mux_v I__7262 (
            .O(N__38520),
            .I(N__38515));
    InMux I__7261 (
            .O(N__38519),
            .I(N__38510));
    InMux I__7260 (
            .O(N__38518),
            .I(N__38510));
    Odrv4 I__7259 (
            .O(N__38515),
            .I(cemf_module_64ch_ctrl_inst1_data_config_22));
    LocalMux I__7258 (
            .O(N__38510),
            .I(cemf_module_64ch_ctrl_inst1_data_config_22));
    CascadeMux I__7257 (
            .O(N__38505),
            .I(N__38502));
    InMux I__7256 (
            .O(N__38502),
            .I(N__38499));
    LocalMux I__7255 (
            .O(N__38499),
            .I(N__38496));
    Span4Mux_h I__7254 (
            .O(N__38496),
            .I(N__38493));
    Span4Mux_h I__7253 (
            .O(N__38493),
            .I(N__38490));
    Odrv4 I__7252 (
            .O(N__38490),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_31));
    InMux I__7251 (
            .O(N__38487),
            .I(N__38484));
    LocalMux I__7250 (
            .O(N__38484),
            .I(N__38481));
    Span4Mux_h I__7249 (
            .O(N__38481),
            .I(N__38476));
    CascadeMux I__7248 (
            .O(N__38480),
            .I(N__38473));
    InMux I__7247 (
            .O(N__38479),
            .I(N__38470));
    Span4Mux_h I__7246 (
            .O(N__38476),
            .I(N__38467));
    InMux I__7245 (
            .O(N__38473),
            .I(N__38464));
    LocalMux I__7244 (
            .O(N__38470),
            .I(N__38461));
    Sp12to4 I__7243 (
            .O(N__38467),
            .I(N__38458));
    LocalMux I__7242 (
            .O(N__38464),
            .I(N__38455));
    Span4Mux_h I__7241 (
            .O(N__38461),
            .I(N__38452));
    Odrv12 I__7240 (
            .O(N__38458),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_14));
    Odrv12 I__7239 (
            .O(N__38455),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_14));
    Odrv4 I__7238 (
            .O(N__38452),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_14));
    CascadeMux I__7237 (
            .O(N__38445),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_22_cascade_ ));
    InMux I__7236 (
            .O(N__38442),
            .I(N__38439));
    LocalMux I__7235 (
            .O(N__38439),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_22 ));
    InMux I__7234 (
            .O(N__38436),
            .I(N__38433));
    LocalMux I__7233 (
            .O(N__38433),
            .I(N__38430));
    Span4Mux_v I__7232 (
            .O(N__38430),
            .I(N__38426));
    CascadeMux I__7231 (
            .O(N__38429),
            .I(N__38422));
    Span4Mux_h I__7230 (
            .O(N__38426),
            .I(N__38419));
    InMux I__7229 (
            .O(N__38425),
            .I(N__38416));
    InMux I__7228 (
            .O(N__38422),
            .I(N__38413));
    Odrv4 I__7227 (
            .O(N__38419),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_22));
    LocalMux I__7226 (
            .O(N__38416),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_22));
    LocalMux I__7225 (
            .O(N__38413),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_22));
    CascadeMux I__7224 (
            .O(N__38406),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_22_cascade_ ));
    InMux I__7223 (
            .O(N__38403),
            .I(N__38400));
    LocalMux I__7222 (
            .O(N__38400),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDDZ0Z7 ));
    CascadeMux I__7221 (
            .O(N__38397),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_21_cascade_ ));
    InMux I__7220 (
            .O(N__38394),
            .I(N__38391));
    LocalMux I__7219 (
            .O(N__38391),
            .I(N__38388));
    Span12Mux_h I__7218 (
            .O(N__38388),
            .I(N__38385));
    Odrv12 I__7217 (
            .O(N__38385),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_21));
    InMux I__7216 (
            .O(N__38382),
            .I(N__38379));
    LocalMux I__7215 (
            .O(N__38379),
            .I(N__38376));
    Span4Mux_v I__7214 (
            .O(N__38376),
            .I(N__38369));
    InMux I__7213 (
            .O(N__38375),
            .I(N__38366));
    InMux I__7212 (
            .O(N__38374),
            .I(N__38363));
    InMux I__7211 (
            .O(N__38373),
            .I(N__38360));
    InMux I__7210 (
            .O(N__38372),
            .I(N__38357));
    Span4Mux_h I__7209 (
            .O(N__38369),
            .I(N__38352));
    LocalMux I__7208 (
            .O(N__38366),
            .I(N__38352));
    LocalMux I__7207 (
            .O(N__38363),
            .I(N__38347));
    LocalMux I__7206 (
            .O(N__38360),
            .I(N__38347));
    LocalMux I__7205 (
            .O(N__38357),
            .I(N__38344));
    Span4Mux_h I__7204 (
            .O(N__38352),
            .I(N__38339));
    Span4Mux_v I__7203 (
            .O(N__38347),
            .I(N__38339));
    Span12Mux_v I__7202 (
            .O(N__38344),
            .I(N__38336));
    Span4Mux_v I__7201 (
            .O(N__38339),
            .I(N__38333));
    Odrv12 I__7200 (
            .O(N__38336),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1320 ));
    Odrv4 I__7199 (
            .O(N__38333),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1320 ));
    InMux I__7198 (
            .O(N__38328),
            .I(N__38325));
    LocalMux I__7197 (
            .O(N__38325),
            .I(N__38322));
    Odrv12 I__7196 (
            .O(N__38322),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1896 ));
    CascadeMux I__7195 (
            .O(N__38319),
            .I(N__38312));
    CascadeMux I__7194 (
            .O(N__38318),
            .I(N__38308));
    CascadeMux I__7193 (
            .O(N__38317),
            .I(N__38305));
    InMux I__7192 (
            .O(N__38316),
            .I(N__38298));
    InMux I__7191 (
            .O(N__38315),
            .I(N__38295));
    InMux I__7190 (
            .O(N__38312),
            .I(N__38292));
    InMux I__7189 (
            .O(N__38311),
            .I(N__38285));
    InMux I__7188 (
            .O(N__38308),
            .I(N__38285));
    InMux I__7187 (
            .O(N__38305),
            .I(N__38285));
    CascadeMux I__7186 (
            .O(N__38304),
            .I(N__38282));
    InMux I__7185 (
            .O(N__38303),
            .I(N__38279));
    InMux I__7184 (
            .O(N__38302),
            .I(N__38273));
    InMux I__7183 (
            .O(N__38301),
            .I(N__38270));
    LocalMux I__7182 (
            .O(N__38298),
            .I(N__38263));
    LocalMux I__7181 (
            .O(N__38295),
            .I(N__38263));
    LocalMux I__7180 (
            .O(N__38292),
            .I(N__38260));
    LocalMux I__7179 (
            .O(N__38285),
            .I(N__38257));
    InMux I__7178 (
            .O(N__38282),
            .I(N__38254));
    LocalMux I__7177 (
            .O(N__38279),
            .I(N__38251));
    InMux I__7176 (
            .O(N__38278),
            .I(N__38248));
    InMux I__7175 (
            .O(N__38277),
            .I(N__38243));
    InMux I__7174 (
            .O(N__38276),
            .I(N__38243));
    LocalMux I__7173 (
            .O(N__38273),
            .I(N__38240));
    LocalMux I__7172 (
            .O(N__38270),
            .I(N__38234));
    InMux I__7171 (
            .O(N__38269),
            .I(N__38231));
    InMux I__7170 (
            .O(N__38268),
            .I(N__38228));
    Span4Mux_v I__7169 (
            .O(N__38263),
            .I(N__38223));
    Span4Mux_v I__7168 (
            .O(N__38260),
            .I(N__38223));
    Span4Mux_v I__7167 (
            .O(N__38257),
            .I(N__38208));
    LocalMux I__7166 (
            .O(N__38254),
            .I(N__38203));
    Span4Mux_v I__7165 (
            .O(N__38251),
            .I(N__38203));
    LocalMux I__7164 (
            .O(N__38248),
            .I(N__38196));
    LocalMux I__7163 (
            .O(N__38243),
            .I(N__38196));
    Span4Mux_v I__7162 (
            .O(N__38240),
            .I(N__38196));
    InMux I__7161 (
            .O(N__38239),
            .I(N__38189));
    InMux I__7160 (
            .O(N__38238),
            .I(N__38189));
    InMux I__7159 (
            .O(N__38237),
            .I(N__38189));
    Span4Mux_h I__7158 (
            .O(N__38234),
            .I(N__38184));
    LocalMux I__7157 (
            .O(N__38231),
            .I(N__38184));
    LocalMux I__7156 (
            .O(N__38228),
            .I(N__38179));
    Span4Mux_h I__7155 (
            .O(N__38223),
            .I(N__38179));
    InMux I__7154 (
            .O(N__38222),
            .I(N__38176));
    InMux I__7153 (
            .O(N__38221),
            .I(N__38161));
    InMux I__7152 (
            .O(N__38220),
            .I(N__38161));
    InMux I__7151 (
            .O(N__38219),
            .I(N__38161));
    InMux I__7150 (
            .O(N__38218),
            .I(N__38161));
    InMux I__7149 (
            .O(N__38217),
            .I(N__38161));
    InMux I__7148 (
            .O(N__38216),
            .I(N__38161));
    InMux I__7147 (
            .O(N__38215),
            .I(N__38161));
    InMux I__7146 (
            .O(N__38214),
            .I(N__38152));
    InMux I__7145 (
            .O(N__38213),
            .I(N__38152));
    InMux I__7144 (
            .O(N__38212),
            .I(N__38152));
    InMux I__7143 (
            .O(N__38211),
            .I(N__38152));
    Span4Mux_v I__7142 (
            .O(N__38208),
            .I(N__38147));
    Span4Mux_h I__7141 (
            .O(N__38203),
            .I(N__38147));
    Span4Mux_h I__7140 (
            .O(N__38196),
            .I(N__38138));
    LocalMux I__7139 (
            .O(N__38189),
            .I(N__38138));
    Span4Mux_v I__7138 (
            .O(N__38184),
            .I(N__38138));
    Span4Mux_h I__7137 (
            .O(N__38179),
            .I(N__38138));
    LocalMux I__7136 (
            .O(N__38176),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ));
    LocalMux I__7135 (
            .O(N__38161),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ));
    LocalMux I__7134 (
            .O(N__38152),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ));
    Odrv4 I__7133 (
            .O(N__38147),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ));
    Odrv4 I__7132 (
            .O(N__38138),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ));
    CascadeMux I__7131 (
            .O(N__38127),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_21_cascade_ ));
    InMux I__7130 (
            .O(N__38124),
            .I(N__38121));
    LocalMux I__7129 (
            .O(N__38121),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_21 ));
    InMux I__7128 (
            .O(N__38118),
            .I(N__38115));
    LocalMux I__7127 (
            .O(N__38115),
            .I(N__38112));
    Span4Mux_h I__7126 (
            .O(N__38112),
            .I(N__38109));
    Odrv4 I__7125 (
            .O(N__38109),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_21 ));
    CascadeMux I__7124 (
            .O(N__38106),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_21_cascade_ ));
    InMux I__7123 (
            .O(N__38103),
            .I(N__38100));
    LocalMux I__7122 (
            .O(N__38100),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_21 ));
    CascadeMux I__7121 (
            .O(N__38097),
            .I(N__38094));
    InMux I__7120 (
            .O(N__38094),
            .I(N__38091));
    LocalMux I__7119 (
            .O(N__38091),
            .I(N__38088));
    Sp12to4 I__7118 (
            .O(N__38088),
            .I(N__38085));
    Span12Mux_v I__7117 (
            .O(N__38085),
            .I(N__38082));
    Odrv12 I__7116 (
            .O(N__38082),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_30));
    InMux I__7115 (
            .O(N__38079),
            .I(N__38074));
    CascadeMux I__7114 (
            .O(N__38078),
            .I(N__38071));
    CascadeMux I__7113 (
            .O(N__38077),
            .I(N__38068));
    LocalMux I__7112 (
            .O(N__38074),
            .I(N__38065));
    InMux I__7111 (
            .O(N__38071),
            .I(N__38062));
    InMux I__7110 (
            .O(N__38068),
            .I(N__38059));
    Span4Mux_v I__7109 (
            .O(N__38065),
            .I(N__38056));
    LocalMux I__7108 (
            .O(N__38062),
            .I(N__38053));
    LocalMux I__7107 (
            .O(N__38059),
            .I(N__38050));
    Span4Mux_h I__7106 (
            .O(N__38056),
            .I(N__38047));
    Span4Mux_v I__7105 (
            .O(N__38053),
            .I(N__38044));
    Span12Mux_h I__7104 (
            .O(N__38050),
            .I(N__38041));
    Odrv4 I__7103 (
            .O(N__38047),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_13));
    Odrv4 I__7102 (
            .O(N__38044),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_13));
    Odrv12 I__7101 (
            .O(N__38041),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_13));
    InMux I__7100 (
            .O(N__38034),
            .I(N__38031));
    LocalMux I__7099 (
            .O(N__38031),
            .I(N__38028));
    Odrv12 I__7098 (
            .O(N__38028),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_20 ));
    InMux I__7097 (
            .O(N__38025),
            .I(N__38022));
    LocalMux I__7096 (
            .O(N__38022),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21 ));
    CascadeMux I__7095 (
            .O(N__38019),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21_cascade_ ));
    CascadeMux I__7094 (
            .O(N__38016),
            .I(N__38013));
    InMux I__7093 (
            .O(N__38013),
            .I(N__38010));
    LocalMux I__7092 (
            .O(N__38010),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_20 ));
    InMux I__7091 (
            .O(N__38007),
            .I(N__38004));
    LocalMux I__7090 (
            .O(N__38004),
            .I(N__38001));
    Odrv4 I__7089 (
            .O(N__38001),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_20 ));
    CascadeMux I__7088 (
            .O(N__37998),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LHZ0Z5_cascade_ ));
    InMux I__7087 (
            .O(N__37995),
            .I(N__37992));
    LocalMux I__7086 (
            .O(N__37992),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20 ));
    CascadeMux I__7085 (
            .O(N__37989),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20_cascade_ ));
    InMux I__7084 (
            .O(N__37986),
            .I(N__37983));
    LocalMux I__7083 (
            .O(N__37983),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_20 ));
    InMux I__7082 (
            .O(N__37980),
            .I(N__37977));
    LocalMux I__7081 (
            .O(N__37977),
            .I(N__37974));
    Span4Mux_h I__7080 (
            .O(N__37974),
            .I(N__37971));
    Span4Mux_h I__7079 (
            .O(N__37971),
            .I(N__37968));
    Span4Mux_v I__7078 (
            .O(N__37968),
            .I(N__37965));
    Span4Mux_v I__7077 (
            .O(N__37965),
            .I(N__37962));
    Odrv4 I__7076 (
            .O(N__37962),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_21));
    CascadeMux I__7075 (
            .O(N__37959),
            .I(N__37956));
    InMux I__7074 (
            .O(N__37956),
            .I(N__37953));
    LocalMux I__7073 (
            .O(N__37953),
            .I(N__37950));
    Span4Mux_v I__7072 (
            .O(N__37950),
            .I(N__37947));
    Span4Mux_h I__7071 (
            .O(N__37947),
            .I(N__37944));
    Span4Mux_h I__7070 (
            .O(N__37944),
            .I(N__37941));
    Odrv4 I__7069 (
            .O(N__37941),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_21));
    CascadeMux I__7068 (
            .O(N__37938),
            .I(N__37935));
    InMux I__7067 (
            .O(N__37935),
            .I(N__37931));
    CascadeMux I__7066 (
            .O(N__37934),
            .I(N__37928));
    LocalMux I__7065 (
            .O(N__37931),
            .I(N__37925));
    InMux I__7064 (
            .O(N__37928),
            .I(N__37922));
    Span12Mux_v I__7063 (
            .O(N__37925),
            .I(N__37919));
    LocalMux I__7062 (
            .O(N__37922),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_23));
    Odrv12 I__7061 (
            .O(N__37919),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_23));
    InMux I__7060 (
            .O(N__37914),
            .I(N__37911));
    LocalMux I__7059 (
            .O(N__37911),
            .I(N__37908));
    Span4Mux_v I__7058 (
            .O(N__37908),
            .I(N__37905));
    Sp12to4 I__7057 (
            .O(N__37905),
            .I(N__37901));
    InMux I__7056 (
            .O(N__37904),
            .I(N__37898));
    Span12Mux_h I__7055 (
            .O(N__37901),
            .I(N__37895));
    LocalMux I__7054 (
            .O(N__37898),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_10));
    Odrv12 I__7053 (
            .O(N__37895),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_10));
    InMux I__7052 (
            .O(N__37890),
            .I(N__37887));
    LocalMux I__7051 (
            .O(N__37887),
            .I(N__37884));
    Odrv12 I__7050 (
            .O(N__37884),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_10 ));
    InMux I__7049 (
            .O(N__37881),
            .I(N__37870));
    InMux I__7048 (
            .O(N__37880),
            .I(N__37848));
    InMux I__7047 (
            .O(N__37879),
            .I(N__37848));
    InMux I__7046 (
            .O(N__37878),
            .I(N__37848));
    InMux I__7045 (
            .O(N__37877),
            .I(N__37848));
    InMux I__7044 (
            .O(N__37876),
            .I(N__37848));
    InMux I__7043 (
            .O(N__37875),
            .I(N__37848));
    InMux I__7042 (
            .O(N__37874),
            .I(N__37848));
    InMux I__7041 (
            .O(N__37873),
            .I(N__37845));
    LocalMux I__7040 (
            .O(N__37870),
            .I(N__37840));
    InMux I__7039 (
            .O(N__37869),
            .I(N__37825));
    InMux I__7038 (
            .O(N__37868),
            .I(N__37825));
    InMux I__7037 (
            .O(N__37867),
            .I(N__37825));
    InMux I__7036 (
            .O(N__37866),
            .I(N__37825));
    InMux I__7035 (
            .O(N__37865),
            .I(N__37825));
    InMux I__7034 (
            .O(N__37864),
            .I(N__37825));
    InMux I__7033 (
            .O(N__37863),
            .I(N__37825));
    LocalMux I__7032 (
            .O(N__37848),
            .I(N__37820));
    LocalMux I__7031 (
            .O(N__37845),
            .I(N__37817));
    InMux I__7030 (
            .O(N__37844),
            .I(N__37814));
    InMux I__7029 (
            .O(N__37843),
            .I(N__37811));
    Span4Mux_v I__7028 (
            .O(N__37840),
            .I(N__37798));
    LocalMux I__7027 (
            .O(N__37825),
            .I(N__37798));
    CascadeMux I__7026 (
            .O(N__37824),
            .I(N__37795));
    CascadeMux I__7025 (
            .O(N__37823),
            .I(N__37792));
    Span4Mux_h I__7024 (
            .O(N__37820),
            .I(N__37789));
    Span4Mux_v I__7023 (
            .O(N__37817),
            .I(N__37784));
    LocalMux I__7022 (
            .O(N__37814),
            .I(N__37784));
    LocalMux I__7021 (
            .O(N__37811),
            .I(N__37781));
    InMux I__7020 (
            .O(N__37810),
            .I(N__37768));
    InMux I__7019 (
            .O(N__37809),
            .I(N__37768));
    InMux I__7018 (
            .O(N__37808),
            .I(N__37768));
    InMux I__7017 (
            .O(N__37807),
            .I(N__37768));
    InMux I__7016 (
            .O(N__37806),
            .I(N__37768));
    InMux I__7015 (
            .O(N__37805),
            .I(N__37768));
    InMux I__7014 (
            .O(N__37804),
            .I(N__37765));
    InMux I__7013 (
            .O(N__37803),
            .I(N__37762));
    Span4Mux_v I__7012 (
            .O(N__37798),
            .I(N__37759));
    InMux I__7011 (
            .O(N__37795),
            .I(N__37754));
    InMux I__7010 (
            .O(N__37792),
            .I(N__37754));
    Span4Mux_v I__7009 (
            .O(N__37789),
            .I(N__37749));
    Span4Mux_h I__7008 (
            .O(N__37784),
            .I(N__37749));
    Span12Mux_v I__7007 (
            .O(N__37781),
            .I(N__37742));
    LocalMux I__7006 (
            .O(N__37768),
            .I(N__37742));
    LocalMux I__7005 (
            .O(N__37765),
            .I(N__37742));
    LocalMux I__7004 (
            .O(N__37762),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable));
    Odrv4 I__7003 (
            .O(N__37759),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable));
    LocalMux I__7002 (
            .O(N__37754),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable));
    Odrv4 I__7001 (
            .O(N__37749),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable));
    Odrv12 I__7000 (
            .O(N__37742),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable));
    CascadeMux I__6999 (
            .O(N__37731),
            .I(N__37728));
    InMux I__6998 (
            .O(N__37728),
            .I(N__37725));
    LocalMux I__6997 (
            .O(N__37725),
            .I(N__37722));
    Span4Mux_v I__6996 (
            .O(N__37722),
            .I(N__37719));
    Sp12to4 I__6995 (
            .O(N__37719),
            .I(N__37716));
    Odrv12 I__6994 (
            .O(N__37716),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_24));
    InMux I__6993 (
            .O(N__37713),
            .I(N__37710));
    LocalMux I__6992 (
            .O(N__37710),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_676 ));
    InMux I__6991 (
            .O(N__37707),
            .I(N__37702));
    InMux I__6990 (
            .O(N__37706),
            .I(N__37695));
    InMux I__6989 (
            .O(N__37705),
            .I(N__37691));
    LocalMux I__6988 (
            .O(N__37702),
            .I(N__37685));
    InMux I__6987 (
            .O(N__37701),
            .I(N__37682));
    InMux I__6986 (
            .O(N__37700),
            .I(N__37675));
    InMux I__6985 (
            .O(N__37699),
            .I(N__37675));
    InMux I__6984 (
            .O(N__37698),
            .I(N__37675));
    LocalMux I__6983 (
            .O(N__37695),
            .I(N__37672));
    InMux I__6982 (
            .O(N__37694),
            .I(N__37669));
    LocalMux I__6981 (
            .O(N__37691),
            .I(N__37666));
    InMux I__6980 (
            .O(N__37690),
            .I(N__37659));
    InMux I__6979 (
            .O(N__37689),
            .I(N__37659));
    InMux I__6978 (
            .O(N__37688),
            .I(N__37659));
    Span4Mux_h I__6977 (
            .O(N__37685),
            .I(N__37635));
    LocalMux I__6976 (
            .O(N__37682),
            .I(N__37635));
    LocalMux I__6975 (
            .O(N__37675),
            .I(N__37632));
    Span4Mux_h I__6974 (
            .O(N__37672),
            .I(N__37627));
    LocalMux I__6973 (
            .O(N__37669),
            .I(N__37627));
    Span4Mux_v I__6972 (
            .O(N__37666),
            .I(N__37622));
    LocalMux I__6971 (
            .O(N__37659),
            .I(N__37622));
    InMux I__6970 (
            .O(N__37658),
            .I(N__37613));
    InMux I__6969 (
            .O(N__37657),
            .I(N__37613));
    InMux I__6968 (
            .O(N__37656),
            .I(N__37613));
    InMux I__6967 (
            .O(N__37655),
            .I(N__37613));
    InMux I__6966 (
            .O(N__37654),
            .I(N__37604));
    InMux I__6965 (
            .O(N__37653),
            .I(N__37604));
    InMux I__6964 (
            .O(N__37652),
            .I(N__37604));
    InMux I__6963 (
            .O(N__37651),
            .I(N__37604));
    InMux I__6962 (
            .O(N__37650),
            .I(N__37589));
    InMux I__6961 (
            .O(N__37649),
            .I(N__37589));
    InMux I__6960 (
            .O(N__37648),
            .I(N__37589));
    InMux I__6959 (
            .O(N__37647),
            .I(N__37589));
    InMux I__6958 (
            .O(N__37646),
            .I(N__37589));
    InMux I__6957 (
            .O(N__37645),
            .I(N__37589));
    InMux I__6956 (
            .O(N__37644),
            .I(N__37589));
    InMux I__6955 (
            .O(N__37643),
            .I(N__37580));
    InMux I__6954 (
            .O(N__37642),
            .I(N__37580));
    InMux I__6953 (
            .O(N__37641),
            .I(N__37580));
    InMux I__6952 (
            .O(N__37640),
            .I(N__37580));
    Span4Mux_v I__6951 (
            .O(N__37635),
            .I(N__37575));
    Span4Mux_v I__6950 (
            .O(N__37632),
            .I(N__37575));
    Span4Mux_v I__6949 (
            .O(N__37627),
            .I(N__37570));
    Span4Mux_h I__6948 (
            .O(N__37622),
            .I(N__37570));
    LocalMux I__6947 (
            .O(N__37613),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ));
    LocalMux I__6946 (
            .O(N__37604),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ));
    LocalMux I__6945 (
            .O(N__37589),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ));
    LocalMux I__6944 (
            .O(N__37580),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ));
    Odrv4 I__6943 (
            .O(N__37575),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ));
    Odrv4 I__6942 (
            .O(N__37570),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ));
    InMux I__6941 (
            .O(N__37557),
            .I(N__37554));
    LocalMux I__6940 (
            .O(N__37554),
            .I(N__37551));
    Odrv12 I__6939 (
            .O(N__37551),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_23 ));
    CascadeMux I__6938 (
            .O(N__37548),
            .I(N__37545));
    InMux I__6937 (
            .O(N__37545),
            .I(N__37542));
    LocalMux I__6936 (
            .O(N__37542),
            .I(N__37539));
    Span4Mux_v I__6935 (
            .O(N__37539),
            .I(N__37536));
    Odrv4 I__6934 (
            .O(N__37536),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_687 ));
    InMux I__6933 (
            .O(N__37533),
            .I(N__37530));
    LocalMux I__6932 (
            .O(N__37530),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_23 ));
    CascadeMux I__6931 (
            .O(N__37527),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_23_cascade_ ));
    InMux I__6930 (
            .O(N__37524),
            .I(N__37521));
    LocalMux I__6929 (
            .O(N__37521),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_23 ));
    InMux I__6928 (
            .O(N__37518),
            .I(N__37515));
    LocalMux I__6927 (
            .O(N__37515),
            .I(N__37512));
    Span4Mux_h I__6926 (
            .O(N__37512),
            .I(N__37509));
    Span4Mux_h I__6925 (
            .O(N__37509),
            .I(N__37506));
    Span4Mux_h I__6924 (
            .O(N__37506),
            .I(N__37503));
    Span4Mux_v I__6923 (
            .O(N__37503),
            .I(N__37500));
    Odrv4 I__6922 (
            .O(N__37500),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_23));
    CascadeMux I__6921 (
            .O(N__37497),
            .I(N__37494));
    InMux I__6920 (
            .O(N__37494),
            .I(N__37491));
    LocalMux I__6919 (
            .O(N__37491),
            .I(N__37488));
    Span4Mux_v I__6918 (
            .O(N__37488),
            .I(N__37485));
    Span4Mux_h I__6917 (
            .O(N__37485),
            .I(N__37482));
    Span4Mux_h I__6916 (
            .O(N__37482),
            .I(N__37479));
    Odrv4 I__6915 (
            .O(N__37479),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_23));
    CascadeMux I__6914 (
            .O(N__37476),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_23_cascade_ ));
    InMux I__6913 (
            .O(N__37473),
            .I(N__37470));
    LocalMux I__6912 (
            .O(N__37470),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_23 ));
    InMux I__6911 (
            .O(N__37467),
            .I(N__37464));
    LocalMux I__6910 (
            .O(N__37464),
            .I(\serializer_mod_inst.shift_regZ0Z_95 ));
    InMux I__6909 (
            .O(N__37461),
            .I(N__37458));
    LocalMux I__6908 (
            .O(N__37458),
            .I(\serializer_mod_inst.shift_regZ0Z_96 ));
    InMux I__6907 (
            .O(N__37455),
            .I(N__37452));
    LocalMux I__6906 (
            .O(N__37452),
            .I(\serializer_mod_inst.shift_regZ0Z_97 ));
    IoInMux I__6905 (
            .O(N__37449),
            .I(N__37446));
    LocalMux I__6904 (
            .O(N__37446),
            .I(N__37443));
    Span12Mux_s3_v I__6903 (
            .O(N__37443),
            .I(N__37440));
    Odrv12 I__6902 (
            .O(N__37440),
            .I(enable_config_c));
    IoInMux I__6901 (
            .O(N__37437),
            .I(N__37434));
    LocalMux I__6900 (
            .O(N__37434),
            .I(N__37431));
    Span12Mux_s9_v I__6899 (
            .O(N__37431),
            .I(N__37428));
    Span12Mux_h I__6898 (
            .O(N__37428),
            .I(N__37425));
    Odrv12 I__6897 (
            .O(N__37425),
            .I(elec_config_out_c));
    InMux I__6896 (
            .O(N__37422),
            .I(N__37419));
    LocalMux I__6895 (
            .O(N__37419),
            .I(N__37416));
    Span4Mux_v I__6894 (
            .O(N__37416),
            .I(N__37413));
    Odrv4 I__6893 (
            .O(N__37413),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_24 ));
    CascadeMux I__6892 (
            .O(N__37410),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_24_cascade_ ));
    InMux I__6891 (
            .O(N__37407),
            .I(N__37404));
    LocalMux I__6890 (
            .O(N__37404),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_24 ));
    InMux I__6889 (
            .O(N__37401),
            .I(N__37398));
    LocalMux I__6888 (
            .O(N__37398),
            .I(N__37395));
    Span4Mux_h I__6887 (
            .O(N__37395),
            .I(N__37392));
    Sp12to4 I__6886 (
            .O(N__37392),
            .I(N__37389));
    Span12Mux_v I__6885 (
            .O(N__37389),
            .I(N__37386));
    Odrv12 I__6884 (
            .O(N__37386),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_24));
    CascadeMux I__6883 (
            .O(N__37383),
            .I(N__37380));
    InMux I__6882 (
            .O(N__37380),
            .I(N__37377));
    LocalMux I__6881 (
            .O(N__37377),
            .I(N__37374));
    Span4Mux_h I__6880 (
            .O(N__37374),
            .I(N__37371));
    Span4Mux_h I__6879 (
            .O(N__37371),
            .I(N__37368));
    Span4Mux_h I__6878 (
            .O(N__37368),
            .I(N__37365));
    Odrv4 I__6877 (
            .O(N__37365),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_24));
    CascadeMux I__6876 (
            .O(N__37362),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_24_cascade_ ));
    InMux I__6875 (
            .O(N__37359),
            .I(N__37356));
    LocalMux I__6874 (
            .O(N__37356),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_24 ));
    InMux I__6873 (
            .O(N__37353),
            .I(N__37350));
    LocalMux I__6872 (
            .O(N__37350),
            .I(\serializer_mod_inst.shift_regZ0Z_106 ));
    InMux I__6871 (
            .O(N__37347),
            .I(N__37344));
    LocalMux I__6870 (
            .O(N__37344),
            .I(N__37341));
    Span4Mux_h I__6869 (
            .O(N__37341),
            .I(N__37338));
    Odrv4 I__6868 (
            .O(N__37338),
            .I(\serializer_mod_inst.shift_regZ0Z_47 ));
    InMux I__6867 (
            .O(N__37335),
            .I(N__37332));
    LocalMux I__6866 (
            .O(N__37332),
            .I(\serializer_mod_inst.shift_regZ0Z_94 ));
    InMux I__6865 (
            .O(N__37329),
            .I(N__37326));
    LocalMux I__6864 (
            .O(N__37326),
            .I(\serializer_mod_inst.shift_regZ0Z_104 ));
    CascadeMux I__6863 (
            .O(N__37323),
            .I(N__37320));
    InMux I__6862 (
            .O(N__37320),
            .I(N__37317));
    LocalMux I__6861 (
            .O(N__37317),
            .I(\serializer_mod_inst.shift_regZ0Z_105 ));
    InMux I__6860 (
            .O(N__37314),
            .I(N__37311));
    LocalMux I__6859 (
            .O(N__37311),
            .I(\serializer_mod_inst.shift_regZ0Z_46 ));
    InMux I__6858 (
            .O(N__37308),
            .I(N__37305));
    LocalMux I__6857 (
            .O(N__37305),
            .I(N__37302));
    Odrv12 I__6856 (
            .O(N__37302),
            .I(\serializer_mod_inst.shift_regZ0Z_91 ));
    InMux I__6855 (
            .O(N__37299),
            .I(N__37296));
    LocalMux I__6854 (
            .O(N__37296),
            .I(\serializer_mod_inst.shift_regZ0Z_92 ));
    InMux I__6853 (
            .O(N__37293),
            .I(N__37290));
    LocalMux I__6852 (
            .O(N__37290),
            .I(\serializer_mod_inst.shift_regZ0Z_93 ));
    InMux I__6851 (
            .O(N__37287),
            .I(N__37284));
    LocalMux I__6850 (
            .O(N__37284),
            .I(\serializer_mod_inst.shift_regZ0Z_15 ));
    InMux I__6849 (
            .O(N__37281),
            .I(N__37278));
    LocalMux I__6848 (
            .O(N__37278),
            .I(\serializer_mod_inst.shift_regZ0Z_79 ));
    InMux I__6847 (
            .O(N__37275),
            .I(N__37272));
    LocalMux I__6846 (
            .O(N__37272),
            .I(\serializer_mod_inst.shift_regZ0Z_16 ));
    InMux I__6845 (
            .O(N__37269),
            .I(N__37266));
    LocalMux I__6844 (
            .O(N__37266),
            .I(\serializer_mod_inst.shift_regZ0Z_17 ));
    InMux I__6843 (
            .O(N__37263),
            .I(N__37260));
    LocalMux I__6842 (
            .O(N__37260),
            .I(\serializer_mod_inst.shift_regZ0Z_18 ));
    InMux I__6841 (
            .O(N__37257),
            .I(N__37254));
    LocalMux I__6840 (
            .O(N__37254),
            .I(\serializer_mod_inst.shift_regZ0Z_107 ));
    InMux I__6839 (
            .O(N__37251),
            .I(N__37248));
    LocalMux I__6838 (
            .O(N__37248),
            .I(\serializer_mod_inst.shift_regZ0Z_69 ));
    InMux I__6837 (
            .O(N__37245),
            .I(N__37242));
    LocalMux I__6836 (
            .O(N__37242),
            .I(\serializer_mod_inst.shift_regZ0Z_51 ));
    InMux I__6835 (
            .O(N__37239),
            .I(N__37236));
    LocalMux I__6834 (
            .O(N__37236),
            .I(\serializer_mod_inst.shift_regZ0Z_10 ));
    InMux I__6833 (
            .O(N__37233),
            .I(N__37230));
    LocalMux I__6832 (
            .O(N__37230),
            .I(N__37227));
    Span4Mux_h I__6831 (
            .O(N__37227),
            .I(N__37224));
    Odrv4 I__6830 (
            .O(N__37224),
            .I(\serializer_mod_inst.shift_regZ0Z_55 ));
    InMux I__6829 (
            .O(N__37221),
            .I(N__37218));
    LocalMux I__6828 (
            .O(N__37218),
            .I(N__37215));
    Odrv4 I__6827 (
            .O(N__37215),
            .I(\serializer_mod_inst.shift_regZ0Z_121 ));
    InMux I__6826 (
            .O(N__37212),
            .I(N__37209));
    LocalMux I__6825 (
            .O(N__37209),
            .I(\serializer_mod_inst.shift_regZ0Z_14 ));
    InMux I__6824 (
            .O(N__37206),
            .I(N__37203));
    LocalMux I__6823 (
            .O(N__37203),
            .I(\serializer_mod_inst.shift_regZ0Z_12 ));
    InMux I__6822 (
            .O(N__37200),
            .I(N__37197));
    LocalMux I__6821 (
            .O(N__37197),
            .I(\serializer_mod_inst.shift_regZ0Z_13 ));
    InMux I__6820 (
            .O(N__37194),
            .I(N__37191));
    LocalMux I__6819 (
            .O(N__37191),
            .I(\serializer_mod_inst.shift_regZ0Z_8 ));
    InMux I__6818 (
            .O(N__37188),
            .I(N__37185));
    LocalMux I__6817 (
            .O(N__37185),
            .I(\serializer_mod_inst.shift_regZ0Z_9 ));
    InMux I__6816 (
            .O(N__37182),
            .I(N__37179));
    LocalMux I__6815 (
            .O(N__37179),
            .I(N__37176));
    Odrv12 I__6814 (
            .O(N__37176),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8Z0Z_26 ));
    InMux I__6813 (
            .O(N__37173),
            .I(N__37170));
    LocalMux I__6812 (
            .O(N__37170),
            .I(N__37165));
    InMux I__6811 (
            .O(N__37169),
            .I(N__37162));
    InMux I__6810 (
            .O(N__37168),
            .I(N__37156));
    Span4Mux_v I__6809 (
            .O(N__37165),
            .I(N__37153));
    LocalMux I__6808 (
            .O(N__37162),
            .I(N__37150));
    InMux I__6807 (
            .O(N__37161),
            .I(N__37145));
    InMux I__6806 (
            .O(N__37160),
            .I(N__37140));
    InMux I__6805 (
            .O(N__37159),
            .I(N__37140));
    LocalMux I__6804 (
            .O(N__37156),
            .I(N__37137));
    Sp12to4 I__6803 (
            .O(N__37153),
            .I(N__37132));
    Span12Mux_v I__6802 (
            .O(N__37150),
            .I(N__37132));
    InMux I__6801 (
            .O(N__37149),
            .I(N__37127));
    InMux I__6800 (
            .O(N__37148),
            .I(N__37127));
    LocalMux I__6799 (
            .O(N__37145),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ));
    LocalMux I__6798 (
            .O(N__37140),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ));
    Odrv4 I__6797 (
            .O(N__37137),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ));
    Odrv12 I__6796 (
            .O(N__37132),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ));
    LocalMux I__6795 (
            .O(N__37127),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ));
    InMux I__6794 (
            .O(N__37116),
            .I(N__37113));
    LocalMux I__6793 (
            .O(N__37113),
            .I(N__37110));
    Span4Mux_h I__6792 (
            .O(N__37110),
            .I(N__37103));
    InMux I__6791 (
            .O(N__37109),
            .I(N__37100));
    InMux I__6790 (
            .O(N__37108),
            .I(N__37097));
    InMux I__6789 (
            .O(N__37107),
            .I(N__37092));
    InMux I__6788 (
            .O(N__37106),
            .I(N__37092));
    Odrv4 I__6787 (
            .O(N__37103),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_12 ));
    LocalMux I__6786 (
            .O(N__37100),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_12 ));
    LocalMux I__6785 (
            .O(N__37097),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_12 ));
    LocalMux I__6784 (
            .O(N__37092),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_12 ));
    InMux I__6783 (
            .O(N__37083),
            .I(N__37077));
    InMux I__6782 (
            .O(N__37082),
            .I(N__37077));
    LocalMux I__6781 (
            .O(N__37077),
            .I(N__37074));
    Span4Mux_v I__6780 (
            .O(N__37074),
            .I(N__37071));
    Odrv4 I__6779 (
            .O(N__37071),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1862 ));
    InMux I__6778 (
            .O(N__37068),
            .I(N__37065));
    LocalMux I__6777 (
            .O(N__37065),
            .I(N__37061));
    InMux I__6776 (
            .O(N__37064),
            .I(N__37058));
    Span4Mux_h I__6775 (
            .O(N__37061),
            .I(N__37053));
    LocalMux I__6774 (
            .O(N__37058),
            .I(N__37053));
    Odrv4 I__6773 (
            .O(N__37053),
            .I(\cemf_module_64ch_ctrl_inst1.N_1816_0 ));
    CascadeMux I__6772 (
            .O(N__37050),
            .I(N__37045));
    InMux I__6771 (
            .O(N__37049),
            .I(N__37042));
    InMux I__6770 (
            .O(N__37048),
            .I(N__37037));
    InMux I__6769 (
            .O(N__37045),
            .I(N__37037));
    LocalMux I__6768 (
            .O(N__37042),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_8 ));
    LocalMux I__6767 (
            .O(N__37037),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_8 ));
    InMux I__6766 (
            .O(N__37032),
            .I(N__37028));
    InMux I__6765 (
            .O(N__37031),
            .I(N__37025));
    LocalMux I__6764 (
            .O(N__37028),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9 ));
    LocalMux I__6763 (
            .O(N__37025),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9 ));
    InMux I__6762 (
            .O(N__37020),
            .I(N__37016));
    InMux I__6761 (
            .O(N__37019),
            .I(N__37013));
    LocalMux I__6760 (
            .O(N__37016),
            .I(N__37008));
    LocalMux I__6759 (
            .O(N__37013),
            .I(N__37008));
    Odrv12 I__6758 (
            .O(N__37008),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_reti_0 ));
    InMux I__6757 (
            .O(N__37005),
            .I(N__37002));
    LocalMux I__6756 (
            .O(N__37002),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_6 ));
    InMux I__6755 (
            .O(N__36999),
            .I(N__36996));
    LocalMux I__6754 (
            .O(N__36996),
            .I(\serializer_mod_inst.shift_regZ0Z_11 ));
    InMux I__6753 (
            .O(N__36993),
            .I(N__36990));
    LocalMux I__6752 (
            .O(N__36990),
            .I(\serializer_mod_inst.shift_regZ0Z_48 ));
    InMux I__6751 (
            .O(N__36987),
            .I(N__36984));
    LocalMux I__6750 (
            .O(N__36984),
            .I(\I2C_top_level_inst1.s_sda_o_qZ0Z_1 ));
    InMux I__6749 (
            .O(N__36981),
            .I(N__36978));
    LocalMux I__6748 (
            .O(N__36978),
            .I(\I2C_top_level_inst1.s_sda_o_txZ0 ));
    InMux I__6747 (
            .O(N__36975),
            .I(N__36972));
    LocalMux I__6746 (
            .O(N__36972),
            .I(\I2C_top_level_inst1.s_sda_o_qZ0Z_0 ));
    InMux I__6745 (
            .O(N__36969),
            .I(N__36964));
    CascadeMux I__6744 (
            .O(N__36968),
            .I(N__36961));
    InMux I__6743 (
            .O(N__36967),
            .I(N__36951));
    LocalMux I__6742 (
            .O(N__36964),
            .I(N__36948));
    InMux I__6741 (
            .O(N__36961),
            .I(N__36939));
    InMux I__6740 (
            .O(N__36960),
            .I(N__36939));
    InMux I__6739 (
            .O(N__36959),
            .I(N__36939));
    InMux I__6738 (
            .O(N__36958),
            .I(N__36939));
    InMux I__6737 (
            .O(N__36957),
            .I(N__36934));
    InMux I__6736 (
            .O(N__36956),
            .I(N__36934));
    InMux I__6735 (
            .O(N__36955),
            .I(N__36929));
    InMux I__6734 (
            .O(N__36954),
            .I(N__36929));
    LocalMux I__6733 (
            .O(N__36951),
            .I(N__36926));
    Span4Mux_v I__6732 (
            .O(N__36948),
            .I(N__36923));
    LocalMux I__6731 (
            .O(N__36939),
            .I(N__36918));
    LocalMux I__6730 (
            .O(N__36934),
            .I(N__36918));
    LocalMux I__6729 (
            .O(N__36929),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_a ));
    Odrv12 I__6728 (
            .O(N__36926),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_a ));
    Odrv4 I__6727 (
            .O(N__36923),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_a ));
    Odrv4 I__6726 (
            .O(N__36918),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_a ));
    CascadeMux I__6725 (
            .O(N__36909),
            .I(N__36905));
    InMux I__6724 (
            .O(N__36908),
            .I(N__36901));
    InMux I__6723 (
            .O(N__36905),
            .I(N__36897));
    InMux I__6722 (
            .O(N__36904),
            .I(N__36894));
    LocalMux I__6721 (
            .O(N__36901),
            .I(N__36891));
    InMux I__6720 (
            .O(N__36900),
            .I(N__36888));
    LocalMux I__6719 (
            .O(N__36897),
            .I(N__36883));
    LocalMux I__6718 (
            .O(N__36894),
            .I(N__36883));
    Span4Mux_h I__6717 (
            .O(N__36891),
            .I(N__36880));
    LocalMux I__6716 (
            .O(N__36888),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0 ));
    Odrv4 I__6715 (
            .O(N__36883),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0 ));
    Odrv4 I__6714 (
            .O(N__36880),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0 ));
    InMux I__6713 (
            .O(N__36873),
            .I(N__36870));
    LocalMux I__6712 (
            .O(N__36870),
            .I(N__36865));
    InMux I__6711 (
            .O(N__36869),
            .I(N__36862));
    InMux I__6710 (
            .O(N__36868),
            .I(N__36859));
    Span4Mux_h I__6709 (
            .O(N__36865),
            .I(N__36856));
    LocalMux I__6708 (
            .O(N__36862),
            .I(N__36851));
    LocalMux I__6707 (
            .O(N__36859),
            .I(N__36851));
    Odrv4 I__6706 (
            .O(N__36856),
            .I(\cemf_module_64ch_ctrl_inst1.N_1855_0 ));
    Odrv12 I__6705 (
            .O(N__36851),
            .I(\cemf_module_64ch_ctrl_inst1.N_1855_0 ));
    CascadeMux I__6704 (
            .O(N__36846),
            .I(\cemf_module_64ch_ctrl_inst1.N_1855_0_cascade_ ));
    CascadeMux I__6703 (
            .O(N__36843),
            .I(N__36840));
    InMux I__6702 (
            .O(N__36840),
            .I(N__36831));
    InMux I__6701 (
            .O(N__36839),
            .I(N__36831));
    InMux I__6700 (
            .O(N__36838),
            .I(N__36828));
    InMux I__6699 (
            .O(N__36837),
            .I(N__36825));
    InMux I__6698 (
            .O(N__36836),
            .I(N__36822));
    LocalMux I__6697 (
            .O(N__36831),
            .I(N__36819));
    LocalMux I__6696 (
            .O(N__36828),
            .I(N__36816));
    LocalMux I__6695 (
            .O(N__36825),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0 ));
    LocalMux I__6694 (
            .O(N__36822),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0 ));
    Odrv4 I__6693 (
            .O(N__36819),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0 ));
    Odrv4 I__6692 (
            .O(N__36816),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0 ));
    InMux I__6691 (
            .O(N__36807),
            .I(N__36804));
    LocalMux I__6690 (
            .O(N__36804),
            .I(N__36801));
    Span4Mux_h I__6689 (
            .O(N__36801),
            .I(N__36798));
    Span4Mux_v I__6688 (
            .O(N__36798),
            .I(N__36795));
    Odrv4 I__6687 (
            .O(N__36795),
            .I(\cemf_module_64ch_ctrl_inst1.N_1857_0 ));
    CascadeMux I__6686 (
            .O(N__36792),
            .I(\cemf_module_64ch_ctrl_inst1.N_1857_0_cascade_ ));
    CascadeMux I__6685 (
            .O(N__36789),
            .I(N__36786));
    InMux I__6684 (
            .O(N__36786),
            .I(N__36780));
    InMux I__6683 (
            .O(N__36785),
            .I(N__36780));
    LocalMux I__6682 (
            .O(N__36780),
            .I(N__36777));
    Span4Mux_v I__6681 (
            .O(N__36777),
            .I(N__36774));
    Odrv4 I__6680 (
            .O(N__36774),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_384 ));
    InMux I__6679 (
            .O(N__36771),
            .I(N__36767));
    InMux I__6678 (
            .O(N__36770),
            .I(N__36764));
    LocalMux I__6677 (
            .O(N__36767),
            .I(N__36759));
    LocalMux I__6676 (
            .O(N__36764),
            .I(N__36759));
    Span12Mux_v I__6675 (
            .O(N__36759),
            .I(N__36756));
    Odrv12 I__6674 (
            .O(N__36756),
            .I(\cemf_module_64ch_ctrl_inst1.N_1854_0 ));
    InMux I__6673 (
            .O(N__36753),
            .I(N__36750));
    LocalMux I__6672 (
            .O(N__36750),
            .I(N__36747));
    Span4Mux_h I__6671 (
            .O(N__36747),
            .I(N__36744));
    Span4Mux_v I__6670 (
            .O(N__36744),
            .I(N__36741));
    Odrv4 I__6669 (
            .O(N__36741),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1840_0 ));
    InMux I__6668 (
            .O(N__36738),
            .I(N__36731));
    InMux I__6667 (
            .O(N__36737),
            .I(N__36722));
    InMux I__6666 (
            .O(N__36736),
            .I(N__36722));
    InMux I__6665 (
            .O(N__36735),
            .I(N__36722));
    InMux I__6664 (
            .O(N__36734),
            .I(N__36722));
    LocalMux I__6663 (
            .O(N__36731),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i ));
    LocalMux I__6662 (
            .O(N__36722),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i ));
    InMux I__6661 (
            .O(N__36717),
            .I(N__36711));
    InMux I__6660 (
            .O(N__36716),
            .I(N__36708));
    InMux I__6659 (
            .O(N__36715),
            .I(N__36703));
    InMux I__6658 (
            .O(N__36714),
            .I(N__36703));
    LocalMux I__6657 (
            .O(N__36711),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0 ));
    LocalMux I__6656 (
            .O(N__36708),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0 ));
    LocalMux I__6655 (
            .O(N__36703),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0 ));
    InMux I__6654 (
            .O(N__36696),
            .I(N__36690));
    InMux I__6653 (
            .O(N__36695),
            .I(N__36690));
    LocalMux I__6652 (
            .O(N__36690),
            .I(N__36686));
    InMux I__6651 (
            .O(N__36689),
            .I(N__36683));
    Odrv4 I__6650 (
            .O(N__36686),
            .I(\cemf_module_64ch_ctrl_inst1.N_383 ));
    LocalMux I__6649 (
            .O(N__36683),
            .I(\cemf_module_64ch_ctrl_inst1.N_383 ));
    InMux I__6648 (
            .O(N__36678),
            .I(N__36672));
    InMux I__6647 (
            .O(N__36677),
            .I(N__36665));
    InMux I__6646 (
            .O(N__36676),
            .I(N__36665));
    InMux I__6645 (
            .O(N__36675),
            .I(N__36665));
    LocalMux I__6644 (
            .O(N__36672),
            .I(N__36662));
    LocalMux I__6643 (
            .O(N__36665),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0 ));
    Odrv4 I__6642 (
            .O(N__36662),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0 ));
    InMux I__6641 (
            .O(N__36657),
            .I(N__36654));
    LocalMux I__6640 (
            .O(N__36654),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_6 ));
    InMux I__6639 (
            .O(N__36651),
            .I(N__36648));
    LocalMux I__6638 (
            .O(N__36648),
            .I(N__36644));
    CascadeMux I__6637 (
            .O(N__36647),
            .I(N__36635));
    Span4Mux_h I__6636 (
            .O(N__36644),
            .I(N__36631));
    InMux I__6635 (
            .O(N__36643),
            .I(N__36626));
    InMux I__6634 (
            .O(N__36642),
            .I(N__36626));
    InMux I__6633 (
            .O(N__36641),
            .I(N__36623));
    InMux I__6632 (
            .O(N__36640),
            .I(N__36616));
    InMux I__6631 (
            .O(N__36639),
            .I(N__36616));
    InMux I__6630 (
            .O(N__36638),
            .I(N__36616));
    InMux I__6629 (
            .O(N__36635),
            .I(N__36611));
    InMux I__6628 (
            .O(N__36634),
            .I(N__36611));
    Odrv4 I__6627 (
            .O(N__36631),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ));
    LocalMux I__6626 (
            .O(N__36626),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ));
    LocalMux I__6625 (
            .O(N__36623),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ));
    LocalMux I__6624 (
            .O(N__36616),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ));
    LocalMux I__6623 (
            .O(N__36611),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ));
    InMux I__6622 (
            .O(N__36600),
            .I(N__36596));
    InMux I__6621 (
            .O(N__36599),
            .I(N__36592));
    LocalMux I__6620 (
            .O(N__36596),
            .I(N__36589));
    InMux I__6619 (
            .O(N__36595),
            .I(N__36586));
    LocalMux I__6618 (
            .O(N__36592),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4 ));
    Odrv4 I__6617 (
            .O(N__36589),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4 ));
    LocalMux I__6616 (
            .O(N__36586),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4 ));
    InMux I__6615 (
            .O(N__36579),
            .I(N__36576));
    LocalMux I__6614 (
            .O(N__36576),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_3_1 ));
    InMux I__6613 (
            .O(N__36573),
            .I(N__36570));
    LocalMux I__6612 (
            .O(N__36570),
            .I(N__36567));
    Span4Mux_v I__6611 (
            .O(N__36567),
            .I(N__36564));
    Odrv4 I__6610 (
            .O(N__36564),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_5_1 ));
    InMux I__6609 (
            .O(N__36561),
            .I(N__36558));
    LocalMux I__6608 (
            .O(N__36558),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_2_1 ));
    CascadeMux I__6607 (
            .O(N__36555),
            .I(\I2C_top_level_inst1.N_4_0_cascade_ ));
    InMux I__6606 (
            .O(N__36552),
            .I(N__36549));
    LocalMux I__6605 (
            .O(N__36549),
            .I(N__36546));
    Span12Mux_h I__6604 (
            .O(N__36546),
            .I(N__36543));
    Odrv12 I__6603 (
            .O(N__36543),
            .I(\I2C_top_level_inst1.N_259 ));
    InMux I__6602 (
            .O(N__36540),
            .I(N__36537));
    LocalMux I__6601 (
            .O(N__36537),
            .I(N__36534));
    Span4Mux_h I__6600 (
            .O(N__36534),
            .I(N__36531));
    Span4Mux_v I__6599 (
            .O(N__36531),
            .I(N__36527));
    InMux I__6598 (
            .O(N__36530),
            .I(N__36524));
    Odrv4 I__6597 (
            .O(N__36527),
            .I(\cemf_module_64ch_ctrl_inst1.N_1848_0 ));
    LocalMux I__6596 (
            .O(N__36524),
            .I(\cemf_module_64ch_ctrl_inst1.N_1848_0 ));
    InMux I__6595 (
            .O(N__36519),
            .I(N__36516));
    LocalMux I__6594 (
            .O(N__36516),
            .I(N__36513));
    Odrv4 I__6593 (
            .O(N__36513),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7Z0Z_26 ));
    CEMux I__6592 (
            .O(N__36510),
            .I(N__36507));
    LocalMux I__6591 (
            .O(N__36507),
            .I(N__36504));
    Span4Mux_v I__6590 (
            .O(N__36504),
            .I(N__36500));
    CEMux I__6589 (
            .O(N__36503),
            .I(N__36497));
    Span4Mux_h I__6588 (
            .O(N__36500),
            .I(N__36494));
    LocalMux I__6587 (
            .O(N__36497),
            .I(N__36491));
    Odrv4 I__6586 (
            .O(N__36494),
            .I(\I2C_top_level_inst1.N_327_i ));
    Odrv12 I__6585 (
            .O(N__36491),
            .I(\I2C_top_level_inst1.N_327_i ));
    InMux I__6584 (
            .O(N__36486),
            .I(N__36483));
    LocalMux I__6583 (
            .O(N__36483),
            .I(N__36480));
    Odrv4 I__6582 (
            .O(N__36480),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1367_0 ));
    InMux I__6581 (
            .O(N__36477),
            .I(N__36474));
    LocalMux I__6580 (
            .O(N__36474),
            .I(N__36469));
    InMux I__6579 (
            .O(N__36473),
            .I(N__36466));
    InMux I__6578 (
            .O(N__36472),
            .I(N__36463));
    Span4Mux_v I__6577 (
            .O(N__36469),
            .I(N__36460));
    LocalMux I__6576 (
            .O(N__36466),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0 ));
    LocalMux I__6575 (
            .O(N__36463),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0 ));
    Odrv4 I__6574 (
            .O(N__36460),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0 ));
    CascadeMux I__6573 (
            .O(N__36453),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1367_0_cascade_ ));
    InMux I__6572 (
            .O(N__36450),
            .I(N__36444));
    InMux I__6571 (
            .O(N__36449),
            .I(N__36444));
    LocalMux I__6570 (
            .O(N__36444),
            .I(N__36441));
    Span4Mux_h I__6569 (
            .O(N__36441),
            .I(N__36438));
    Odrv4 I__6568 (
            .O(N__36438),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_113_0 ));
    InMux I__6567 (
            .O(N__36435),
            .I(N__36432));
    LocalMux I__6566 (
            .O(N__36432),
            .I(N__36428));
    InMux I__6565 (
            .O(N__36431),
            .I(N__36425));
    Span4Mux_h I__6564 (
            .O(N__36428),
            .I(N__36422));
    LocalMux I__6563 (
            .O(N__36425),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1 ));
    Odrv4 I__6562 (
            .O(N__36422),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1 ));
    CascadeMux I__6561 (
            .O(N__36417),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0_cascade_ ));
    InMux I__6560 (
            .O(N__36414),
            .I(N__36411));
    LocalMux I__6559 (
            .O(N__36411),
            .I(\I2C_top_level_inst1.s_command_4 ));
    InMux I__6558 (
            .O(N__36408),
            .I(N__36405));
    LocalMux I__6557 (
            .O(N__36405),
            .I(\I2C_top_level_inst1.s_command_5 ));
    InMux I__6556 (
            .O(N__36402),
            .I(N__36399));
    LocalMux I__6555 (
            .O(N__36399),
            .I(\I2C_top_level_inst1.s_command_6 ));
    InMux I__6554 (
            .O(N__36396),
            .I(N__36393));
    LocalMux I__6553 (
            .O(N__36393),
            .I(N__36390));
    Odrv4 I__6552 (
            .O(N__36390),
            .I(N_1803));
    CascadeMux I__6551 (
            .O(N__36387),
            .I(N_1803_cascade_));
    CascadeMux I__6550 (
            .O(N__36384),
            .I(N__36381));
    InMux I__6549 (
            .O(N__36381),
            .I(N__36378));
    LocalMux I__6548 (
            .O(N__36378),
            .I(\I2C_top_level_inst1.s_command_7 ));
    InMux I__6547 (
            .O(N__36375),
            .I(N__36372));
    LocalMux I__6546 (
            .O(N__36372),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6Z0Z_26 ));
    CascadeMux I__6545 (
            .O(N__36369),
            .I(N_1613_cascade_));
    InMux I__6544 (
            .O(N__36366),
            .I(N__36363));
    LocalMux I__6543 (
            .O(N__36363),
            .I(N__36359));
    InMux I__6542 (
            .O(N__36362),
            .I(N__36356));
    Sp12to4 I__6541 (
            .O(N__36359),
            .I(N__36351));
    LocalMux I__6540 (
            .O(N__36356),
            .I(N__36348));
    InMux I__6539 (
            .O(N__36355),
            .I(N__36345));
    InMux I__6538 (
            .O(N__36354),
            .I(N__36342));
    Span12Mux_s7_v I__6537 (
            .O(N__36351),
            .I(N__36339));
    Span4Mux_v I__6536 (
            .O(N__36348),
            .I(N__36336));
    LocalMux I__6535 (
            .O(N__36345),
            .I(N__36333));
    LocalMux I__6534 (
            .O(N__36342),
            .I(N_1860_0));
    Odrv12 I__6533 (
            .O(N__36339),
            .I(N_1860_0));
    Odrv4 I__6532 (
            .O(N__36336),
            .I(N_1860_0));
    Odrv12 I__6531 (
            .O(N__36333),
            .I(N_1860_0));
    InMux I__6530 (
            .O(N__36324),
            .I(N__36321));
    LocalMux I__6529 (
            .O(N__36321),
            .I(N__36318));
    Span4Mux_h I__6528 (
            .O(N__36318),
            .I(N__36314));
    InMux I__6527 (
            .O(N__36317),
            .I(N__36311));
    Odrv4 I__6526 (
            .O(N__36314),
            .I(N_202_0));
    LocalMux I__6525 (
            .O(N__36311),
            .I(N_202_0));
    InMux I__6524 (
            .O(N__36306),
            .I(N__36302));
    InMux I__6523 (
            .O(N__36305),
            .I(N__36299));
    LocalMux I__6522 (
            .O(N__36302),
            .I(N__36296));
    LocalMux I__6521 (
            .O(N__36299),
            .I(N__36291));
    Span4Mux_h I__6520 (
            .O(N__36296),
            .I(N__36288));
    InMux I__6519 (
            .O(N__36295),
            .I(N__36283));
    InMux I__6518 (
            .O(N__36294),
            .I(N__36283));
    Span4Mux_v I__6517 (
            .O(N__36291),
            .I(N__36280));
    Odrv4 I__6516 (
            .O(N__36288),
            .I(N_1859_0));
    LocalMux I__6515 (
            .O(N__36283),
            .I(N_1859_0));
    Odrv4 I__6514 (
            .O(N__36280),
            .I(N_1859_0));
    CascadeMux I__6513 (
            .O(N__36273),
            .I(N__36269));
    InMux I__6512 (
            .O(N__36272),
            .I(N__36265));
    InMux I__6511 (
            .O(N__36269),
            .I(N__36260));
    InMux I__6510 (
            .O(N__36268),
            .I(N__36260));
    LocalMux I__6509 (
            .O(N__36265),
            .I(N__36256));
    LocalMux I__6508 (
            .O(N__36260),
            .I(N__36253));
    InMux I__6507 (
            .O(N__36259),
            .I(N__36250));
    Span4Mux_h I__6506 (
            .O(N__36256),
            .I(N__36247));
    Span4Mux_v I__6505 (
            .O(N__36253),
            .I(N__36244));
    LocalMux I__6504 (
            .O(N__36250),
            .I(N_1861_0));
    Odrv4 I__6503 (
            .O(N__36247),
            .I(N_1861_0));
    Odrv4 I__6502 (
            .O(N__36244),
            .I(N_1861_0));
    InMux I__6501 (
            .O(N__36237),
            .I(N__36228));
    InMux I__6500 (
            .O(N__36236),
            .I(N__36228));
    InMux I__6499 (
            .O(N__36235),
            .I(N__36228));
    LocalMux I__6498 (
            .O(N__36228),
            .I(N__36225));
    Span4Mux_h I__6497 (
            .O(N__36225),
            .I(N__36222));
    Span4Mux_h I__6496 (
            .O(N__36222),
            .I(N__36215));
    InMux I__6495 (
            .O(N__36221),
            .I(N__36206));
    InMux I__6494 (
            .O(N__36220),
            .I(N__36206));
    InMux I__6493 (
            .O(N__36219),
            .I(N__36206));
    InMux I__6492 (
            .O(N__36218),
            .I(N__36206));
    Odrv4 I__6491 (
            .O(N__36215),
            .I(N_1613));
    LocalMux I__6490 (
            .O(N__36206),
            .I(N_1613));
    InMux I__6489 (
            .O(N__36201),
            .I(N__36198));
    LocalMux I__6488 (
            .O(N__36198),
            .I(N__36195));
    Odrv12 I__6487 (
            .O(N__36195),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_604 ));
    CascadeMux I__6486 (
            .O(N__36192),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20_cascade_ ));
    InMux I__6485 (
            .O(N__36189),
            .I(N__36186));
    LocalMux I__6484 (
            .O(N__36186),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_20 ));
    InMux I__6483 (
            .O(N__36183),
            .I(N__36179));
    InMux I__6482 (
            .O(N__36182),
            .I(N__36176));
    LocalMux I__6481 (
            .O(N__36179),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21 ));
    LocalMux I__6480 (
            .O(N__36176),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21 ));
    InMux I__6479 (
            .O(N__36171),
            .I(N__36168));
    LocalMux I__6478 (
            .O(N__36168),
            .I(N__36165));
    Sp12to4 I__6477 (
            .O(N__36165),
            .I(N__36162));
    Odrv12 I__6476 (
            .O(N__36162),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_21 ));
    InMux I__6475 (
            .O(N__36159),
            .I(N__36155));
    InMux I__6474 (
            .O(N__36158),
            .I(N__36152));
    LocalMux I__6473 (
            .O(N__36155),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22 ));
    LocalMux I__6472 (
            .O(N__36152),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22 ));
    InMux I__6471 (
            .O(N__36147),
            .I(N__36144));
    LocalMux I__6470 (
            .O(N__36144),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_22 ));
    InMux I__6469 (
            .O(N__36141),
            .I(N__36137));
    InMux I__6468 (
            .O(N__36140),
            .I(N__36134));
    LocalMux I__6467 (
            .O(N__36137),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23 ));
    LocalMux I__6466 (
            .O(N__36134),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23 ));
    InMux I__6465 (
            .O(N__36129),
            .I(N__36126));
    LocalMux I__6464 (
            .O(N__36126),
            .I(N__36123));
    Span4Mux_v I__6463 (
            .O(N__36123),
            .I(N__36120));
    Sp12to4 I__6462 (
            .O(N__36120),
            .I(N__36117));
    Odrv12 I__6461 (
            .O(N__36117),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_conf ));
    CascadeMux I__6460 (
            .O(N__36114),
            .I(N__36110));
    CascadeMux I__6459 (
            .O(N__36113),
            .I(N__36107));
    CascadeBuf I__6458 (
            .O(N__36110),
            .I(N__36104));
    CascadeBuf I__6457 (
            .O(N__36107),
            .I(N__36101));
    CascadeMux I__6456 (
            .O(N__36104),
            .I(N__36098));
    CascadeMux I__6455 (
            .O(N__36101),
            .I(N__36095));
    CascadeBuf I__6454 (
            .O(N__36098),
            .I(N__36092));
    CascadeBuf I__6453 (
            .O(N__36095),
            .I(N__36089));
    CascadeMux I__6452 (
            .O(N__36092),
            .I(N__36086));
    CascadeMux I__6451 (
            .O(N__36089),
            .I(N__36083));
    CascadeBuf I__6450 (
            .O(N__36086),
            .I(N__36080));
    CascadeBuf I__6449 (
            .O(N__36083),
            .I(N__36077));
    CascadeMux I__6448 (
            .O(N__36080),
            .I(N__36074));
    CascadeMux I__6447 (
            .O(N__36077),
            .I(N__36071));
    CascadeBuf I__6446 (
            .O(N__36074),
            .I(N__36068));
    CascadeBuf I__6445 (
            .O(N__36071),
            .I(N__36065));
    CascadeMux I__6444 (
            .O(N__36068),
            .I(N__36062));
    CascadeMux I__6443 (
            .O(N__36065),
            .I(N__36059));
    CascadeBuf I__6442 (
            .O(N__36062),
            .I(N__36056));
    CascadeBuf I__6441 (
            .O(N__36059),
            .I(N__36053));
    CascadeMux I__6440 (
            .O(N__36056),
            .I(N__36050));
    CascadeMux I__6439 (
            .O(N__36053),
            .I(N__36047));
    CascadeBuf I__6438 (
            .O(N__36050),
            .I(N__36044));
    CascadeBuf I__6437 (
            .O(N__36047),
            .I(N__36041));
    CascadeMux I__6436 (
            .O(N__36044),
            .I(N__36038));
    CascadeMux I__6435 (
            .O(N__36041),
            .I(N__36035));
    CascadeBuf I__6434 (
            .O(N__36038),
            .I(N__36032));
    CascadeBuf I__6433 (
            .O(N__36035),
            .I(N__36029));
    CascadeMux I__6432 (
            .O(N__36032),
            .I(N__36026));
    CascadeMux I__6431 (
            .O(N__36029),
            .I(N__36023));
    InMux I__6430 (
            .O(N__36026),
            .I(N__36020));
    InMux I__6429 (
            .O(N__36023),
            .I(N__36017));
    LocalMux I__6428 (
            .O(N__36020),
            .I(N__36014));
    LocalMux I__6427 (
            .O(N__36017),
            .I(N__36011));
    Span4Mux_v I__6426 (
            .O(N__36014),
            .I(N__36006));
    Span4Mux_h I__6425 (
            .O(N__36011),
            .I(N__36006));
    Span4Mux_h I__6424 (
            .O(N__36006),
            .I(N__36003));
    Span4Mux_h I__6423 (
            .O(N__36003),
            .I(N__36000));
    Odrv4 I__6422 (
            .O(N__36000),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1831_0 ));
    CascadeMux I__6421 (
            .O(N__35997),
            .I(N__35993));
    InMux I__6420 (
            .O(N__35996),
            .I(N__35983));
    InMux I__6419 (
            .O(N__35993),
            .I(N__35974));
    InMux I__6418 (
            .O(N__35992),
            .I(N__35974));
    InMux I__6417 (
            .O(N__35991),
            .I(N__35974));
    InMux I__6416 (
            .O(N__35990),
            .I(N__35974));
    InMux I__6415 (
            .O(N__35989),
            .I(N__35968));
    InMux I__6414 (
            .O(N__35988),
            .I(N__35968));
    InMux I__6413 (
            .O(N__35987),
            .I(N__35963));
    InMux I__6412 (
            .O(N__35986),
            .I(N__35963));
    LocalMux I__6411 (
            .O(N__35983),
            .I(N__35960));
    LocalMux I__6410 (
            .O(N__35974),
            .I(N__35957));
    InMux I__6409 (
            .O(N__35973),
            .I(N__35954));
    LocalMux I__6408 (
            .O(N__35968),
            .I(N__35949));
    LocalMux I__6407 (
            .O(N__35963),
            .I(N__35949));
    Span4Mux_v I__6406 (
            .O(N__35960),
            .I(N__35944));
    Span4Mux_v I__6405 (
            .O(N__35957),
            .I(N__35944));
    LocalMux I__6404 (
            .O(N__35954),
            .I(N__35941));
    Span4Mux_v I__6403 (
            .O(N__35949),
            .I(N__35938));
    Span4Mux_h I__6402 (
            .O(N__35944),
            .I(N__35935));
    Span4Mux_h I__6401 (
            .O(N__35941),
            .I(N__35930));
    Span4Mux_v I__6400 (
            .O(N__35938),
            .I(N__35930));
    Odrv4 I__6399 (
            .O(N__35935),
            .I(N_1614));
    Odrv4 I__6398 (
            .O(N__35930),
            .I(N_1614));
    CascadeMux I__6397 (
            .O(N__35925),
            .I(N_1841_0_cascade_));
    InMux I__6396 (
            .O(N__35922),
            .I(N__35919));
    LocalMux I__6395 (
            .O(N__35919),
            .I(N__35916));
    Span4Mux_h I__6394 (
            .O(N__35916),
            .I(N__35912));
    InMux I__6393 (
            .O(N__35915),
            .I(N__35909));
    Span4Mux_v I__6392 (
            .O(N__35912),
            .I(N__35906));
    LocalMux I__6391 (
            .O(N__35909),
            .I(N__35903));
    Span4Mux_v I__6390 (
            .O(N__35906),
            .I(N__35900));
    Sp12to4 I__6389 (
            .O(N__35903),
            .I(N__35897));
    Odrv4 I__6388 (
            .O(N__35900),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0 ));
    Odrv12 I__6387 (
            .O(N__35897),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0 ));
    InMux I__6386 (
            .O(N__35892),
            .I(N__35889));
    LocalMux I__6385 (
            .O(N__35889),
            .I(N__35885));
    InMux I__6384 (
            .O(N__35888),
            .I(N__35882));
    Span4Mux_h I__6383 (
            .O(N__35885),
            .I(N__35878));
    LocalMux I__6382 (
            .O(N__35882),
            .I(N__35875));
    InMux I__6381 (
            .O(N__35881),
            .I(N__35872));
    Span4Mux_v I__6380 (
            .O(N__35878),
            .I(N__35869));
    Odrv4 I__6379 (
            .O(N__35875),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4 ));
    LocalMux I__6378 (
            .O(N__35872),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4 ));
    Odrv4 I__6377 (
            .O(N__35869),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4 ));
    InMux I__6376 (
            .O(N__35862),
            .I(N__35857));
    InMux I__6375 (
            .O(N__35861),
            .I(N__35848));
    InMux I__6374 (
            .O(N__35860),
            .I(N__35848));
    LocalMux I__6373 (
            .O(N__35857),
            .I(N__35845));
    InMux I__6372 (
            .O(N__35856),
            .I(N__35838));
    InMux I__6371 (
            .O(N__35855),
            .I(N__35838));
    InMux I__6370 (
            .O(N__35854),
            .I(N__35838));
    InMux I__6369 (
            .O(N__35853),
            .I(N__35835));
    LocalMux I__6368 (
            .O(N__35848),
            .I(N__35832));
    Span4Mux_h I__6367 (
            .O(N__35845),
            .I(N__35829));
    LocalMux I__6366 (
            .O(N__35838),
            .I(N__35826));
    LocalMux I__6365 (
            .O(N__35835),
            .I(N__35823));
    Span4Mux_v I__6364 (
            .O(N__35832),
            .I(N__35820));
    Span4Mux_v I__6363 (
            .O(N__35829),
            .I(N__35813));
    Span4Mux_h I__6362 (
            .O(N__35826),
            .I(N__35813));
    Span4Mux_v I__6361 (
            .O(N__35823),
            .I(N__35808));
    Span4Mux_h I__6360 (
            .O(N__35820),
            .I(N__35808));
    InMux I__6359 (
            .O(N__35819),
            .I(N__35803));
    InMux I__6358 (
            .O(N__35818),
            .I(N__35803));
    Odrv4 I__6357 (
            .O(N__35813),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_b ));
    Odrv4 I__6356 (
            .O(N__35808),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_b ));
    LocalMux I__6355 (
            .O(N__35803),
            .I(\cemf_module_64ch_ctrl_inst1.start_conf_b ));
    InMux I__6354 (
            .O(N__35796),
            .I(N__35792));
    InMux I__6353 (
            .O(N__35795),
            .I(N__35789));
    LocalMux I__6352 (
            .O(N__35792),
            .I(N__35786));
    LocalMux I__6351 (
            .O(N__35789),
            .I(N__35783));
    Span4Mux_v I__6350 (
            .O(N__35786),
            .I(N__35780));
    Sp12to4 I__6349 (
            .O(N__35783),
            .I(N__35777));
    Span4Mux_v I__6348 (
            .O(N__35780),
            .I(N__35774));
    Span12Mux_v I__6347 (
            .O(N__35777),
            .I(N__35771));
    Sp12to4 I__6346 (
            .O(N__35774),
            .I(N__35768));
    Odrv12 I__6345 (
            .O(N__35771),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0 ));
    Odrv12 I__6344 (
            .O(N__35768),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0 ));
    CascadeMux I__6343 (
            .O(N__35763),
            .I(N__35758));
    InMux I__6342 (
            .O(N__35762),
            .I(N__35752));
    InMux I__6341 (
            .O(N__35761),
            .I(N__35749));
    InMux I__6340 (
            .O(N__35758),
            .I(N__35743));
    InMux I__6339 (
            .O(N__35757),
            .I(N__35743));
    InMux I__6338 (
            .O(N__35756),
            .I(N__35738));
    InMux I__6337 (
            .O(N__35755),
            .I(N__35738));
    LocalMux I__6336 (
            .O(N__35752),
            .I(N__35735));
    LocalMux I__6335 (
            .O(N__35749),
            .I(N__35732));
    InMux I__6334 (
            .O(N__35748),
            .I(N__35729));
    LocalMux I__6333 (
            .O(N__35743),
            .I(N__35726));
    LocalMux I__6332 (
            .O(N__35738),
            .I(N__35719));
    Span4Mux_v I__6331 (
            .O(N__35735),
            .I(N__35719));
    Sp12to4 I__6330 (
            .O(N__35732),
            .I(N__35716));
    LocalMux I__6329 (
            .O(N__35729),
            .I(N__35711));
    Span4Mux_h I__6328 (
            .O(N__35726),
            .I(N__35711));
    InMux I__6327 (
            .O(N__35725),
            .I(N__35708));
    InMux I__6326 (
            .O(N__35724),
            .I(N__35705));
    Sp12to4 I__6325 (
            .O(N__35719),
            .I(N__35700));
    Span12Mux_v I__6324 (
            .O(N__35716),
            .I(N__35700));
    Odrv4 I__6323 (
            .O(N__35711),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15 ));
    LocalMux I__6322 (
            .O(N__35708),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15 ));
    LocalMux I__6321 (
            .O(N__35705),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15 ));
    Odrv12 I__6320 (
            .O(N__35700),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15 ));
    InMux I__6319 (
            .O(N__35691),
            .I(N__35688));
    LocalMux I__6318 (
            .O(N__35688),
            .I(N__35685));
    Span4Mux_v I__6317 (
            .O(N__35685),
            .I(N__35682));
    Sp12to4 I__6316 (
            .O(N__35682),
            .I(N__35677));
    InMux I__6315 (
            .O(N__35681),
            .I(N__35672));
    InMux I__6314 (
            .O(N__35680),
            .I(N__35672));
    Odrv12 I__6313 (
            .O(N__35677),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_20));
    LocalMux I__6312 (
            .O(N__35672),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_20));
    CascadeMux I__6311 (
            .O(N__35667),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_20_cascade_ ));
    CascadeMux I__6310 (
            .O(N__35664),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DDZ0Z7_cascade_ ));
    InMux I__6309 (
            .O(N__35661),
            .I(N__35658));
    LocalMux I__6308 (
            .O(N__35658),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20 ));
    InMux I__6307 (
            .O(N__35655),
            .I(N__35652));
    LocalMux I__6306 (
            .O(N__35652),
            .I(N__35648));
    InMux I__6305 (
            .O(N__35651),
            .I(N__35645));
    Span4Mux_v I__6304 (
            .O(N__35648),
            .I(N__35642));
    LocalMux I__6303 (
            .O(N__35645),
            .I(N__35639));
    Span4Mux_h I__6302 (
            .O(N__35642),
            .I(N__35636));
    Odrv4 I__6301 (
            .O(N__35639),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_28));
    Odrv4 I__6300 (
            .O(N__35636),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_28));
    InMux I__6299 (
            .O(N__35631),
            .I(N__35628));
    LocalMux I__6298 (
            .O(N__35628),
            .I(N__35625));
    Span4Mux_h I__6297 (
            .O(N__35625),
            .I(N__35622));
    Odrv4 I__6296 (
            .O(N__35622),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_28 ));
    CascadeMux I__6295 (
            .O(N__35619),
            .I(N__35616));
    InMux I__6294 (
            .O(N__35616),
            .I(N__35613));
    LocalMux I__6293 (
            .O(N__35613),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_28));
    InMux I__6292 (
            .O(N__35610),
            .I(N__35607));
    LocalMux I__6291 (
            .O(N__35607),
            .I(N__35604));
    Span4Mux_v I__6290 (
            .O(N__35604),
            .I(N__35600));
    InMux I__6289 (
            .O(N__35603),
            .I(N__35597));
    Span4Mux_h I__6288 (
            .O(N__35600),
            .I(N__35594));
    LocalMux I__6287 (
            .O(N__35597),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_29));
    Odrv4 I__6286 (
            .O(N__35594),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_29));
    CascadeMux I__6285 (
            .O(N__35589),
            .I(N__35586));
    InMux I__6284 (
            .O(N__35586),
            .I(N__35583));
    LocalMux I__6283 (
            .O(N__35583),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_29));
    InMux I__6282 (
            .O(N__35580),
            .I(N__35577));
    LocalMux I__6281 (
            .O(N__35577),
            .I(N__35574));
    Span4Mux_v I__6280 (
            .O(N__35574),
            .I(N__35570));
    CascadeMux I__6279 (
            .O(N__35573),
            .I(N__35567));
    Span4Mux_h I__6278 (
            .O(N__35570),
            .I(N__35564));
    InMux I__6277 (
            .O(N__35567),
            .I(N__35561));
    Sp12to4 I__6276 (
            .O(N__35564),
            .I(N__35558));
    LocalMux I__6275 (
            .O(N__35561),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_3));
    Odrv12 I__6274 (
            .O(N__35558),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_3));
    InMux I__6273 (
            .O(N__35553),
            .I(N__35550));
    LocalMux I__6272 (
            .O(N__35550),
            .I(N__35547));
    Span4Mux_h I__6271 (
            .O(N__35547),
            .I(N__35544));
    Span4Mux_h I__6270 (
            .O(N__35544),
            .I(N__35541));
    Odrv4 I__6269 (
            .O(N__35541),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_3 ));
    CascadeMux I__6268 (
            .O(N__35538),
            .I(N__35534));
    InMux I__6267 (
            .O(N__35537),
            .I(N__35530));
    InMux I__6266 (
            .O(N__35534),
            .I(N__35527));
    CascadeMux I__6265 (
            .O(N__35533),
            .I(N__35524));
    LocalMux I__6264 (
            .O(N__35530),
            .I(N__35519));
    LocalMux I__6263 (
            .O(N__35527),
            .I(N__35519));
    InMux I__6262 (
            .O(N__35524),
            .I(N__35516));
    Span4Mux_h I__6261 (
            .O(N__35519),
            .I(N__35513));
    LocalMux I__6260 (
            .O(N__35516),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_3));
    Odrv4 I__6259 (
            .O(N__35513),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_3));
    IoInMux I__6258 (
            .O(N__35508),
            .I(N__35505));
    LocalMux I__6257 (
            .O(N__35505),
            .I(N__35502));
    IoSpan4Mux I__6256 (
            .O(N__35502),
            .I(N__35499));
    Span4Mux_s2_h I__6255 (
            .O(N__35499),
            .I(N__35496));
    Sp12to4 I__6254 (
            .O(N__35496),
            .I(N__35493));
    Span12Mux_h I__6253 (
            .O(N__35493),
            .I(N__35490));
    Odrv12 I__6252 (
            .O(N__35490),
            .I(serial_out_testing_c));
    CascadeMux I__6251 (
            .O(N__35487),
            .I(N__35484));
    InMux I__6250 (
            .O(N__35484),
            .I(N__35474));
    InMux I__6249 (
            .O(N__35483),
            .I(N__35474));
    InMux I__6248 (
            .O(N__35482),
            .I(N__35474));
    CEMux I__6247 (
            .O(N__35481),
            .I(N__35471));
    LocalMux I__6246 (
            .O(N__35474),
            .I(N__35468));
    LocalMux I__6245 (
            .O(N__35471),
            .I(N__35465));
    Span4Mux_h I__6244 (
            .O(N__35468),
            .I(N__35461));
    Span4Mux_h I__6243 (
            .O(N__35465),
            .I(N__35458));
    InMux I__6242 (
            .O(N__35464),
            .I(N__35454));
    Span4Mux_h I__6241 (
            .O(N__35461),
            .I(N__35451));
    Span4Mux_h I__6240 (
            .O(N__35458),
            .I(N__35448));
    InMux I__6239 (
            .O(N__35457),
            .I(N__35445));
    LocalMux I__6238 (
            .O(N__35454),
            .I(N__35442));
    Sp12to4 I__6237 (
            .O(N__35451),
            .I(N__35439));
    Span4Mux_h I__6236 (
            .O(N__35448),
            .I(N__35436));
    LocalMux I__6235 (
            .O(N__35445),
            .I(N__35433));
    Span4Mux_h I__6234 (
            .O(N__35442),
            .I(N__35430));
    Span12Mux_v I__6233 (
            .O(N__35439),
            .I(N__35427));
    Sp12to4 I__6232 (
            .O(N__35436),
            .I(N__35424));
    Span12Mux_h I__6231 (
            .O(N__35433),
            .I(N__35421));
    Span4Mux_h I__6230 (
            .O(N__35430),
            .I(N__35418));
    Span12Mux_h I__6229 (
            .O(N__35427),
            .I(N__35415));
    Span12Mux_v I__6228 (
            .O(N__35424),
            .I(N__35410));
    Span12Mux_h I__6227 (
            .O(N__35421),
            .I(N__35410));
    Span4Mux_h I__6226 (
            .O(N__35418),
            .I(N__35407));
    Odrv12 I__6225 (
            .O(N__35415),
            .I(rst_n_c));
    Odrv12 I__6224 (
            .O(N__35410),
            .I(rst_n_c));
    Odrv4 I__6223 (
            .O(N__35407),
            .I(rst_n_c));
    InMux I__6222 (
            .O(N__35400),
            .I(N__35397));
    LocalMux I__6221 (
            .O(N__35397),
            .I(N__35391));
    InMux I__6220 (
            .O(N__35396),
            .I(N__35388));
    InMux I__6219 (
            .O(N__35395),
            .I(N__35383));
    InMux I__6218 (
            .O(N__35394),
            .I(N__35383));
    Span4Mux_h I__6217 (
            .O(N__35391),
            .I(N__35380));
    LocalMux I__6216 (
            .O(N__35388),
            .I(N__35375));
    LocalMux I__6215 (
            .O(N__35383),
            .I(N__35375));
    Sp12to4 I__6214 (
            .O(N__35380),
            .I(N__35370));
    Span12Mux_h I__6213 (
            .O(N__35375),
            .I(N__35370));
    Odrv12 I__6212 (
            .O(N__35370),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1965 ));
    InMux I__6211 (
            .O(N__35367),
            .I(N__35364));
    LocalMux I__6210 (
            .O(N__35364),
            .I(N__35361));
    Span4Mux_v I__6209 (
            .O(N__35361),
            .I(N__35357));
    InMux I__6208 (
            .O(N__35360),
            .I(N__35354));
    Sp12to4 I__6207 (
            .O(N__35357),
            .I(N__35351));
    LocalMux I__6206 (
            .O(N__35354),
            .I(N__35348));
    Span12Mux_h I__6205 (
            .O(N__35351),
            .I(N__35343));
    Sp12to4 I__6204 (
            .O(N__35348),
            .I(N__35343));
    Odrv12 I__6203 (
            .O(N__35343),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_522_0 ));
    CascadeMux I__6202 (
            .O(N__35340),
            .I(N__35337));
    InMux I__6201 (
            .O(N__35337),
            .I(N__35334));
    LocalMux I__6200 (
            .O(N__35334),
            .I(N__35331));
    Span4Mux_h I__6199 (
            .O(N__35331),
            .I(N__35327));
    InMux I__6198 (
            .O(N__35330),
            .I(N__35324));
    Span4Mux_h I__6197 (
            .O(N__35327),
            .I(N__35321));
    LocalMux I__6196 (
            .O(N__35324),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_17));
    Odrv4 I__6195 (
            .O(N__35321),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_17));
    InMux I__6194 (
            .O(N__35316),
            .I(N__35313));
    LocalMux I__6193 (
            .O(N__35313),
            .I(N__35310));
    Span4Mux_h I__6192 (
            .O(N__35310),
            .I(N__35307));
    Odrv4 I__6191 (
            .O(N__35307),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_17 ));
    InMux I__6190 (
            .O(N__35304),
            .I(N__35300));
    CascadeMux I__6189 (
            .O(N__35303),
            .I(N__35297));
    LocalMux I__6188 (
            .O(N__35300),
            .I(N__35294));
    InMux I__6187 (
            .O(N__35297),
            .I(N__35291));
    Span4Mux_v I__6186 (
            .O(N__35294),
            .I(N__35288));
    LocalMux I__6185 (
            .O(N__35291),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_2));
    Odrv4 I__6184 (
            .O(N__35288),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_2));
    CascadeMux I__6183 (
            .O(N__35283),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0_cascade_ ));
    InMux I__6182 (
            .O(N__35280),
            .I(N__35277));
    LocalMux I__6181 (
            .O(N__35277),
            .I(N__35274));
    Span4Mux_h I__6180 (
            .O(N__35274),
            .I(N__35271));
    Odrv4 I__6179 (
            .O(N__35271),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_2 ));
    InMux I__6178 (
            .O(N__35268),
            .I(N__35265));
    LocalMux I__6177 (
            .O(N__35265),
            .I(N__35261));
    InMux I__6176 (
            .O(N__35264),
            .I(N__35258));
    Span4Mux_h I__6175 (
            .O(N__35261),
            .I(N__35255));
    LocalMux I__6174 (
            .O(N__35258),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_24));
    Odrv4 I__6173 (
            .O(N__35255),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_24));
    CascadeMux I__6172 (
            .O(N__35250),
            .I(N__35247));
    InMux I__6171 (
            .O(N__35247),
            .I(N__35244));
    LocalMux I__6170 (
            .O(N__35244),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_24));
    CascadeMux I__6169 (
            .O(N__35241),
            .I(N__35238));
    InMux I__6168 (
            .O(N__35238),
            .I(N__35235));
    LocalMux I__6167 (
            .O(N__35235),
            .I(N__35231));
    InMux I__6166 (
            .O(N__35234),
            .I(N__35228));
    Sp12to4 I__6165 (
            .O(N__35231),
            .I(N__35225));
    LocalMux I__6164 (
            .O(N__35228),
            .I(N__35220));
    Span12Mux_v I__6163 (
            .O(N__35225),
            .I(N__35220));
    Odrv12 I__6162 (
            .O(N__35220),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_19));
    InMux I__6161 (
            .O(N__35217),
            .I(N__35214));
    LocalMux I__6160 (
            .O(N__35214),
            .I(N__35211));
    Span4Mux_v I__6159 (
            .O(N__35211),
            .I(N__35208));
    Odrv4 I__6158 (
            .O(N__35208),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_19 ));
    InMux I__6157 (
            .O(N__35205),
            .I(N__35202));
    LocalMux I__6156 (
            .O(N__35202),
            .I(N__35199));
    Span4Mux_v I__6155 (
            .O(N__35199),
            .I(N__35195));
    InMux I__6154 (
            .O(N__35198),
            .I(N__35192));
    Span4Mux_h I__6153 (
            .O(N__35195),
            .I(N__35189));
    LocalMux I__6152 (
            .O(N__35192),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_25));
    Odrv4 I__6151 (
            .O(N__35189),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_25));
    InMux I__6150 (
            .O(N__35184),
            .I(N__35181));
    LocalMux I__6149 (
            .O(N__35181),
            .I(N__35178));
    Span4Mux_h I__6148 (
            .O(N__35178),
            .I(N__35174));
    InMux I__6147 (
            .O(N__35177),
            .I(N__35171));
    Span4Mux_h I__6146 (
            .O(N__35174),
            .I(N__35168));
    LocalMux I__6145 (
            .O(N__35171),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_27));
    Odrv4 I__6144 (
            .O(N__35168),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_27));
    CascadeMux I__6143 (
            .O(N__35163),
            .I(N__35160));
    InMux I__6142 (
            .O(N__35160),
            .I(N__35157));
    LocalMux I__6141 (
            .O(N__35157),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_27));
    InMux I__6140 (
            .O(N__35154),
            .I(N__35151));
    LocalMux I__6139 (
            .O(N__35151),
            .I(N__35148));
    Span4Mux_h I__6138 (
            .O(N__35148),
            .I(N__35145));
    Span4Mux_h I__6137 (
            .O(N__35145),
            .I(N__35142));
    Span4Mux_h I__6136 (
            .O(N__35142),
            .I(N__35139));
    Odrv4 I__6135 (
            .O(N__35139),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_12));
    InMux I__6134 (
            .O(N__35136),
            .I(N__35133));
    LocalMux I__6133 (
            .O(N__35133),
            .I(N__35130));
    Span12Mux_v I__6132 (
            .O(N__35130),
            .I(N__35127));
    Odrv12 I__6131 (
            .O(N__35127),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_808 ));
    CascadeMux I__6130 (
            .O(N__35124),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_12_cascade_ ));
    InMux I__6129 (
            .O(N__35121),
            .I(N__35118));
    LocalMux I__6128 (
            .O(N__35118),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_12 ));
    CascadeMux I__6127 (
            .O(N__35115),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_12_cascade_ ));
    InMux I__6126 (
            .O(N__35112),
            .I(N__35109));
    LocalMux I__6125 (
            .O(N__35109),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_12 ));
    CascadeMux I__6124 (
            .O(N__35106),
            .I(N__35103));
    InMux I__6123 (
            .O(N__35103),
            .I(N__35100));
    LocalMux I__6122 (
            .O(N__35100),
            .I(N__35096));
    CascadeMux I__6121 (
            .O(N__35099),
            .I(N__35093));
    Span4Mux_v I__6120 (
            .O(N__35096),
            .I(N__35090));
    InMux I__6119 (
            .O(N__35093),
            .I(N__35087));
    Span4Mux_v I__6118 (
            .O(N__35090),
            .I(N__35084));
    LocalMux I__6117 (
            .O(N__35087),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_11));
    Odrv4 I__6116 (
            .O(N__35084),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_11));
    InMux I__6115 (
            .O(N__35079),
            .I(N__35076));
    LocalMux I__6114 (
            .O(N__35076),
            .I(N__35073));
    Odrv4 I__6113 (
            .O(N__35073),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_11 ));
    CascadeMux I__6112 (
            .O(N__35070),
            .I(N__35067));
    InMux I__6111 (
            .O(N__35067),
            .I(N__35064));
    LocalMux I__6110 (
            .O(N__35064),
            .I(N__35061));
    Span4Mux_h I__6109 (
            .O(N__35061),
            .I(N__35057));
    CascadeMux I__6108 (
            .O(N__35060),
            .I(N__35054));
    Span4Mux_v I__6107 (
            .O(N__35057),
            .I(N__35051));
    InMux I__6106 (
            .O(N__35054),
            .I(N__35048));
    Sp12to4 I__6105 (
            .O(N__35051),
            .I(N__35045));
    LocalMux I__6104 (
            .O(N__35048),
            .I(N__35040));
    Span12Mux_v I__6103 (
            .O(N__35045),
            .I(N__35040));
    Odrv12 I__6102 (
            .O(N__35040),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_12));
    InMux I__6101 (
            .O(N__35037),
            .I(N__35034));
    LocalMux I__6100 (
            .O(N__35034),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_12 ));
    CascadeMux I__6099 (
            .O(N__35031),
            .I(N__35028));
    InMux I__6098 (
            .O(N__35028),
            .I(N__35025));
    LocalMux I__6097 (
            .O(N__35025),
            .I(N__35022));
    Span4Mux_v I__6096 (
            .O(N__35022),
            .I(N__35019));
    Span4Mux_v I__6095 (
            .O(N__35019),
            .I(N__35015));
    InMux I__6094 (
            .O(N__35018),
            .I(N__35012));
    Sp12to4 I__6093 (
            .O(N__35015),
            .I(N__35009));
    LocalMux I__6092 (
            .O(N__35012),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_13));
    Odrv12 I__6091 (
            .O(N__35009),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_13));
    InMux I__6090 (
            .O(N__35004),
            .I(N__35001));
    LocalMux I__6089 (
            .O(N__35001),
            .I(N__34998));
    Span4Mux_h I__6088 (
            .O(N__34998),
            .I(N__34995));
    Odrv4 I__6087 (
            .O(N__34995),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_13 ));
    CascadeMux I__6086 (
            .O(N__34992),
            .I(N__34989));
    InMux I__6085 (
            .O(N__34989),
            .I(N__34985));
    CascadeMux I__6084 (
            .O(N__34988),
            .I(N__34982));
    LocalMux I__6083 (
            .O(N__34985),
            .I(N__34979));
    InMux I__6082 (
            .O(N__34982),
            .I(N__34976));
    Span12Mux_v I__6081 (
            .O(N__34979),
            .I(N__34973));
    LocalMux I__6080 (
            .O(N__34976),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_14));
    Odrv12 I__6079 (
            .O(N__34973),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_14));
    InMux I__6078 (
            .O(N__34968),
            .I(N__34965));
    LocalMux I__6077 (
            .O(N__34965),
            .I(N__34962));
    Span4Mux_h I__6076 (
            .O(N__34962),
            .I(N__34959));
    Span4Mux_h I__6075 (
            .O(N__34959),
            .I(N__34956));
    Odrv4 I__6074 (
            .O(N__34956),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_14 ));
    CascadeMux I__6073 (
            .O(N__34953),
            .I(N__34950));
    InMux I__6072 (
            .O(N__34950),
            .I(N__34947));
    LocalMux I__6071 (
            .O(N__34947),
            .I(N__34944));
    Span4Mux_h I__6070 (
            .O(N__34944),
            .I(N__34940));
    CascadeMux I__6069 (
            .O(N__34943),
            .I(N__34937));
    Span4Mux_v I__6068 (
            .O(N__34940),
            .I(N__34934));
    InMux I__6067 (
            .O(N__34937),
            .I(N__34931));
    Span4Mux_v I__6066 (
            .O(N__34934),
            .I(N__34928));
    LocalMux I__6065 (
            .O(N__34931),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_15));
    Odrv4 I__6064 (
            .O(N__34928),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_15));
    InMux I__6063 (
            .O(N__34923),
            .I(N__34920));
    LocalMux I__6062 (
            .O(N__34920),
            .I(N__34917));
    Odrv12 I__6061 (
            .O(N__34917),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_15 ));
    CascadeMux I__6060 (
            .O(N__34914),
            .I(N__34911));
    InMux I__6059 (
            .O(N__34911),
            .I(N__34907));
    CascadeMux I__6058 (
            .O(N__34910),
            .I(N__34904));
    LocalMux I__6057 (
            .O(N__34907),
            .I(N__34901));
    InMux I__6056 (
            .O(N__34904),
            .I(N__34898));
    Span4Mux_v I__6055 (
            .O(N__34901),
            .I(N__34895));
    LocalMux I__6054 (
            .O(N__34898),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_16));
    Odrv4 I__6053 (
            .O(N__34895),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_16));
    InMux I__6052 (
            .O(N__34890),
            .I(N__34887));
    LocalMux I__6051 (
            .O(N__34887),
            .I(\serializer_mod_inst.shift_regZ0Z_67 ));
    InMux I__6050 (
            .O(N__34884),
            .I(N__34881));
    LocalMux I__6049 (
            .O(N__34881),
            .I(\serializer_mod_inst.shift_regZ0Z_68 ));
    InMux I__6048 (
            .O(N__34878),
            .I(N__34875));
    LocalMux I__6047 (
            .O(N__34875),
            .I(N__34872));
    Odrv4 I__6046 (
            .O(N__34872),
            .I(\serializer_mod_inst.shift_regZ0Z_115 ));
    InMux I__6045 (
            .O(N__34869),
            .I(N__34866));
    LocalMux I__6044 (
            .O(N__34866),
            .I(\serializer_mod_inst.shift_regZ0Z_116 ));
    InMux I__6043 (
            .O(N__34863),
            .I(N__34860));
    LocalMux I__6042 (
            .O(N__34860),
            .I(\serializer_mod_inst.shift_regZ0Z_117 ));
    InMux I__6041 (
            .O(N__34857),
            .I(N__34853));
    InMux I__6040 (
            .O(N__34856),
            .I(N__34848));
    LocalMux I__6039 (
            .O(N__34853),
            .I(N__34845));
    InMux I__6038 (
            .O(N__34852),
            .I(N__34840));
    InMux I__6037 (
            .O(N__34851),
            .I(N__34837));
    LocalMux I__6036 (
            .O(N__34848),
            .I(N__34832));
    Span12Mux_s6_v I__6035 (
            .O(N__34845),
            .I(N__34832));
    InMux I__6034 (
            .O(N__34844),
            .I(N__34827));
    InMux I__6033 (
            .O(N__34843),
            .I(N__34827));
    LocalMux I__6032 (
            .O(N__34840),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0 ));
    LocalMux I__6031 (
            .O(N__34837),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0 ));
    Odrv12 I__6030 (
            .O(N__34832),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0 ));
    LocalMux I__6029 (
            .O(N__34827),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0 ));
    IoInMux I__6028 (
            .O(N__34818),
            .I(N__34815));
    LocalMux I__6027 (
            .O(N__34815),
            .I(N__34812));
    Span4Mux_s2_v I__6026 (
            .O(N__34812),
            .I(N__34809));
    Odrv4 I__6025 (
            .O(N__34809),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa ));
    IoInMux I__6024 (
            .O(N__34806),
            .I(N__34803));
    LocalMux I__6023 (
            .O(N__34803),
            .I(rst_n_c_i));
    InMux I__6022 (
            .O(N__34800),
            .I(N__34797));
    LocalMux I__6021 (
            .O(N__34797),
            .I(N__34794));
    Span4Mux_h I__6020 (
            .O(N__34794),
            .I(N__34791));
    Span4Mux_h I__6019 (
            .O(N__34791),
            .I(N__34788));
    Span4Mux_v I__6018 (
            .O(N__34788),
            .I(N__34785));
    Span4Mux_v I__6017 (
            .O(N__34785),
            .I(N__34782));
    Odrv4 I__6016 (
            .O(N__34782),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_12));
    CascadeMux I__6015 (
            .O(N__34779),
            .I(N__34776));
    InMux I__6014 (
            .O(N__34776),
            .I(N__34773));
    LocalMux I__6013 (
            .O(N__34773),
            .I(N__34770));
    Span4Mux_h I__6012 (
            .O(N__34770),
            .I(N__34767));
    Span4Mux_v I__6011 (
            .O(N__34767),
            .I(N__34764));
    Span4Mux_h I__6010 (
            .O(N__34764),
            .I(N__34761));
    Odrv4 I__6009 (
            .O(N__34761),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_12));
    CascadeMux I__6008 (
            .O(N__34758),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_12_cascade_ ));
    InMux I__6007 (
            .O(N__34755),
            .I(N__34752));
    LocalMux I__6006 (
            .O(N__34752),
            .I(N__34749));
    Odrv4 I__6005 (
            .O(N__34749),
            .I(\serializer_mod_inst.shift_regZ0Z_113 ));
    InMux I__6004 (
            .O(N__34746),
            .I(N__34743));
    LocalMux I__6003 (
            .O(N__34743),
            .I(\serializer_mod_inst.shift_regZ0Z_114 ));
    InMux I__6002 (
            .O(N__34740),
            .I(N__34737));
    LocalMux I__6001 (
            .O(N__34737),
            .I(\serializer_mod_inst.shift_regZ0Z_110 ));
    InMux I__6000 (
            .O(N__34734),
            .I(N__34731));
    LocalMux I__5999 (
            .O(N__34731),
            .I(\serializer_mod_inst.shift_regZ0Z_39 ));
    InMux I__5998 (
            .O(N__34728),
            .I(N__34725));
    LocalMux I__5997 (
            .O(N__34725),
            .I(\serializer_mod_inst.shift_regZ0Z_77 ));
    InMux I__5996 (
            .O(N__34722),
            .I(N__34719));
    LocalMux I__5995 (
            .O(N__34719),
            .I(\serializer_mod_inst.shift_regZ0Z_78 ));
    InMux I__5994 (
            .O(N__34716),
            .I(N__34713));
    LocalMux I__5993 (
            .O(N__34713),
            .I(\serializer_mod_inst.shift_regZ0Z_40 ));
    CascadeMux I__5992 (
            .O(N__34710),
            .I(N__34707));
    InMux I__5991 (
            .O(N__34707),
            .I(N__34704));
    LocalMux I__5990 (
            .O(N__34704),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0 ));
    InMux I__5989 (
            .O(N__34701),
            .I(N__34698));
    LocalMux I__5988 (
            .O(N__34698),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_2 ));
    InMux I__5987 (
            .O(N__34695),
            .I(N__34692));
    LocalMux I__5986 (
            .O(N__34692),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_12 ));
    InMux I__5985 (
            .O(N__34689),
            .I(N__34686));
    LocalMux I__5984 (
            .O(N__34686),
            .I(N__34683));
    Odrv4 I__5983 (
            .O(N__34683),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_li_0_1 ));
    InMux I__5982 (
            .O(N__34680),
            .I(N__34677));
    LocalMux I__5981 (
            .O(N__34677),
            .I(c_state_ret_12_RNIDMPS1_0));
    CascadeMux I__5980 (
            .O(N__34674),
            .I(c_state_ret_12_RNIDMPS1_0_cascade_));
    CascadeMux I__5979 (
            .O(N__34671),
            .I(N__34667));
    InMux I__5978 (
            .O(N__34670),
            .I(N__34662));
    InMux I__5977 (
            .O(N__34667),
            .I(N__34662));
    LocalMux I__5976 (
            .O(N__34662),
            .I(N__34659));
    Span4Mux_v I__5975 (
            .O(N__34659),
            .I(N__34656));
    Span4Mux_v I__5974 (
            .O(N__34656),
            .I(N__34651));
    InMux I__5973 (
            .O(N__34655),
            .I(N__34646));
    InMux I__5972 (
            .O(N__34654),
            .I(N__34646));
    Odrv4 I__5971 (
            .O(N__34651),
            .I(\cemf_module_64ch_ctrl_inst1.clr_sys_reg ));
    LocalMux I__5970 (
            .O(N__34646),
            .I(\cemf_module_64ch_ctrl_inst1.clr_sys_reg ));
    CascadeMux I__5969 (
            .O(N__34641),
            .I(N__34636));
    CascadeMux I__5968 (
            .O(N__34640),
            .I(N__34633));
    CascadeMux I__5967 (
            .O(N__34639),
            .I(N__34630));
    InMux I__5966 (
            .O(N__34636),
            .I(N__34626));
    InMux I__5965 (
            .O(N__34633),
            .I(N__34621));
    InMux I__5964 (
            .O(N__34630),
            .I(N__34621));
    InMux I__5963 (
            .O(N__34629),
            .I(N__34618));
    LocalMux I__5962 (
            .O(N__34626),
            .I(N__34615));
    LocalMux I__5961 (
            .O(N__34621),
            .I(N__34612));
    LocalMux I__5960 (
            .O(N__34618),
            .I(N__34609));
    Span4Mux_v I__5959 (
            .O(N__34615),
            .I(N__34604));
    Span4Mux_v I__5958 (
            .O(N__34612),
            .I(N__34604));
    Odrv12 I__5957 (
            .O(N__34609),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_1));
    Odrv4 I__5956 (
            .O(N__34604),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_1));
    InMux I__5955 (
            .O(N__34599),
            .I(N__34594));
    InMux I__5954 (
            .O(N__34598),
            .I(N__34589));
    InMux I__5953 (
            .O(N__34597),
            .I(N__34589));
    LocalMux I__5952 (
            .O(N__34594),
            .I(N__34584));
    LocalMux I__5951 (
            .O(N__34589),
            .I(N__34584));
    Span4Mux_v I__5950 (
            .O(N__34584),
            .I(N__34581));
    Span4Mux_v I__5949 (
            .O(N__34581),
            .I(N__34578));
    Odrv4 I__5948 (
            .O(N__34578),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_349 ));
    InMux I__5947 (
            .O(N__34575),
            .I(N__34572));
    LocalMux I__5946 (
            .O(N__34572),
            .I(\serializer_mod_inst.shift_regZ0Z_7 ));
    InMux I__5945 (
            .O(N__34569),
            .I(N__34566));
    LocalMux I__5944 (
            .O(N__34566),
            .I(\serializer_mod_inst.shift_regZ0Z_31 ));
    InMux I__5943 (
            .O(N__34563),
            .I(N__34560));
    LocalMux I__5942 (
            .O(N__34560),
            .I(\serializer_mod_inst.shift_regZ0Z_32 ));
    CascadeMux I__5941 (
            .O(N__34557),
            .I(N__34552));
    InMux I__5940 (
            .O(N__34556),
            .I(N__34544));
    InMux I__5939 (
            .O(N__34555),
            .I(N__34544));
    InMux I__5938 (
            .O(N__34552),
            .I(N__34544));
    CascadeMux I__5937 (
            .O(N__34551),
            .I(N__34540));
    LocalMux I__5936 (
            .O(N__34544),
            .I(N__34537));
    InMux I__5935 (
            .O(N__34543),
            .I(N__34532));
    InMux I__5934 (
            .O(N__34540),
            .I(N__34532));
    Span4Mux_h I__5933 (
            .O(N__34537),
            .I(N__34529));
    LocalMux I__5932 (
            .O(N__34532),
            .I(N__34526));
    Odrv4 I__5931 (
            .O(N__34529),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13 ));
    Odrv4 I__5930 (
            .O(N__34526),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13 ));
    InMux I__5929 (
            .O(N__34521),
            .I(N__34518));
    LocalMux I__5928 (
            .O(N__34518),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1880 ));
    CascadeMux I__5927 (
            .O(N__34515),
            .I(\cemf_module_64ch_ctrl_inst1.N_1848_0_cascade_ ));
    InMux I__5926 (
            .O(N__34512),
            .I(N__34508));
    InMux I__5925 (
            .O(N__34511),
            .I(N__34505));
    LocalMux I__5924 (
            .O(N__34508),
            .I(N__34502));
    LocalMux I__5923 (
            .O(N__34505),
            .I(N__34497));
    Span4Mux_v I__5922 (
            .O(N__34502),
            .I(N__34497));
    Odrv4 I__5921 (
            .O(N__34497),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1884_0 ));
    InMux I__5920 (
            .O(N__34494),
            .I(N__34491));
    LocalMux I__5919 (
            .O(N__34491),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0 ));
    CascadeMux I__5918 (
            .O(N__34488),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0_cascade_ ));
    InMux I__5917 (
            .O(N__34485),
            .I(N__34482));
    LocalMux I__5916 (
            .O(N__34482),
            .I(N__34479));
    Odrv4 I__5915 (
            .O(N__34479),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392_reti ));
    CascadeMux I__5914 (
            .O(N__34476),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0_a2_6_1_cascade_ ));
    CascadeMux I__5913 (
            .O(N__34473),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1399_cascade_ ));
    CascadeMux I__5912 (
            .O(N__34470),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1373_0_cascade_ ));
    CascadeMux I__5911 (
            .O(N__34467),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1395_cascade_ ));
    InMux I__5910 (
            .O(N__34464),
            .I(N__34461));
    LocalMux I__5909 (
            .O(N__34461),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_0_10 ));
    CascadeMux I__5908 (
            .O(N__34458),
            .I(N__34450));
    InMux I__5907 (
            .O(N__34457),
            .I(N__34442));
    InMux I__5906 (
            .O(N__34456),
            .I(N__34442));
    InMux I__5905 (
            .O(N__34455),
            .I(N__34442));
    InMux I__5904 (
            .O(N__34454),
            .I(N__34433));
    InMux I__5903 (
            .O(N__34453),
            .I(N__34433));
    InMux I__5902 (
            .O(N__34450),
            .I(N__34433));
    InMux I__5901 (
            .O(N__34449),
            .I(N__34433));
    LocalMux I__5900 (
            .O(N__34442),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10 ));
    LocalMux I__5899 (
            .O(N__34433),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10 ));
    InMux I__5898 (
            .O(N__34428),
            .I(N__34425));
    LocalMux I__5897 (
            .O(N__34425),
            .I(N__34422));
    Span4Mux_v I__5896 (
            .O(N__34422),
            .I(N__34417));
    InMux I__5895 (
            .O(N__34421),
            .I(N__34414));
    InMux I__5894 (
            .O(N__34420),
            .I(N__34411));
    Odrv4 I__5893 (
            .O(N__34417),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8 ));
    LocalMux I__5892 (
            .O(N__34414),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8 ));
    LocalMux I__5891 (
            .O(N__34411),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8 ));
    InMux I__5890 (
            .O(N__34404),
            .I(N__34400));
    InMux I__5889 (
            .O(N__34403),
            .I(N__34397));
    LocalMux I__5888 (
            .O(N__34400),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1373_0 ));
    LocalMux I__5887 (
            .O(N__34397),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1373_0 ));
    InMux I__5886 (
            .O(N__34392),
            .I(N__34389));
    LocalMux I__5885 (
            .O(N__34389),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_14 ));
    CascadeMux I__5884 (
            .O(N__34386),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1409_cascade_ ));
    InMux I__5883 (
            .O(N__34383),
            .I(N__34376));
    InMux I__5882 (
            .O(N__34382),
            .I(N__34376));
    InMux I__5881 (
            .O(N__34381),
            .I(N__34372));
    LocalMux I__5880 (
            .O(N__34376),
            .I(N__34369));
    InMux I__5879 (
            .O(N__34375),
            .I(N__34366));
    LocalMux I__5878 (
            .O(N__34372),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1372_0 ));
    Odrv4 I__5877 (
            .O(N__34369),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1372_0 ));
    LocalMux I__5876 (
            .O(N__34366),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1372_0 ));
    InMux I__5875 (
            .O(N__34359),
            .I(N__34355));
    CascadeMux I__5874 (
            .O(N__34358),
            .I(N__34351));
    LocalMux I__5873 (
            .O(N__34355),
            .I(N__34348));
    InMux I__5872 (
            .O(N__34354),
            .I(N__34343));
    InMux I__5871 (
            .O(N__34351),
            .I(N__34343));
    Span4Mux_h I__5870 (
            .O(N__34348),
            .I(N__34340));
    LocalMux I__5869 (
            .O(N__34343),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14 ));
    Odrv4 I__5868 (
            .O(N__34340),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14 ));
    InMux I__5867 (
            .O(N__34335),
            .I(N__34317));
    InMux I__5866 (
            .O(N__34334),
            .I(N__34317));
    InMux I__5865 (
            .O(N__34333),
            .I(N__34317));
    InMux I__5864 (
            .O(N__34332),
            .I(N__34317));
    InMux I__5863 (
            .O(N__34331),
            .I(N__34317));
    InMux I__5862 (
            .O(N__34330),
            .I(N__34317));
    LocalMux I__5861 (
            .O(N__34317),
            .I(N__34314));
    Span4Mux_v I__5860 (
            .O(N__34314),
            .I(N__34310));
    InMux I__5859 (
            .O(N__34313),
            .I(N__34307));
    Odrv4 I__5858 (
            .O(N__34310),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1379_0 ));
    LocalMux I__5857 (
            .O(N__34307),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1379_0 ));
    CascadeMux I__5856 (
            .O(N__34302),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1400_cascade_ ));
    InMux I__5855 (
            .O(N__34299),
            .I(N__34296));
    LocalMux I__5854 (
            .O(N__34296),
            .I(N__34292));
    InMux I__5853 (
            .O(N__34295),
            .I(N__34289));
    Span4Mux_v I__5852 (
            .O(N__34292),
            .I(N__34286));
    LocalMux I__5851 (
            .O(N__34289),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1374_0 ));
    Odrv4 I__5850 (
            .O(N__34286),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1374_0 ));
    InMux I__5849 (
            .O(N__34281),
            .I(N__34277));
    InMux I__5848 (
            .O(N__34280),
            .I(N__34273));
    LocalMux I__5847 (
            .O(N__34277),
            .I(N__34269));
    InMux I__5846 (
            .O(N__34276),
            .I(N__34266));
    LocalMux I__5845 (
            .O(N__34273),
            .I(N__34263));
    InMux I__5844 (
            .O(N__34272),
            .I(N__34260));
    Span4Mux_h I__5843 (
            .O(N__34269),
            .I(N__34257));
    LocalMux I__5842 (
            .O(N__34266),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0 ));
    Odrv12 I__5841 (
            .O(N__34263),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0 ));
    LocalMux I__5840 (
            .O(N__34260),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0 ));
    Odrv4 I__5839 (
            .O(N__34257),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0 ));
    InMux I__5838 (
            .O(N__34248),
            .I(N__34245));
    LocalMux I__5837 (
            .O(N__34245),
            .I(N__34241));
    InMux I__5836 (
            .O(N__34244),
            .I(N__34237));
    Span4Mux_h I__5835 (
            .O(N__34241),
            .I(N__34234));
    InMux I__5834 (
            .O(N__34240),
            .I(N__34231));
    LocalMux I__5833 (
            .O(N__34237),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2 ));
    Odrv4 I__5832 (
            .O(N__34234),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2 ));
    LocalMux I__5831 (
            .O(N__34231),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2 ));
    CascadeMux I__5830 (
            .O(N__34224),
            .I(N__34221));
    InMux I__5829 (
            .O(N__34221),
            .I(N__34218));
    LocalMux I__5828 (
            .O(N__34218),
            .I(N__34213));
    InMux I__5827 (
            .O(N__34217),
            .I(N__34210));
    InMux I__5826 (
            .O(N__34216),
            .I(N__34207));
    Span4Mux_h I__5825 (
            .O(N__34213),
            .I(N__34204));
    LocalMux I__5824 (
            .O(N__34210),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3 ));
    LocalMux I__5823 (
            .O(N__34207),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3 ));
    Odrv4 I__5822 (
            .O(N__34204),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3 ));
    InMux I__5821 (
            .O(N__34197),
            .I(N__34194));
    LocalMux I__5820 (
            .O(N__34194),
            .I(N__34191));
    Span4Mux_h I__5819 (
            .O(N__34191),
            .I(N__34186));
    InMux I__5818 (
            .O(N__34190),
            .I(N__34183));
    InMux I__5817 (
            .O(N__34189),
            .I(N__34180));
    Odrv4 I__5816 (
            .O(N__34186),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1 ));
    LocalMux I__5815 (
            .O(N__34183),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1 ));
    LocalMux I__5814 (
            .O(N__34180),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1 ));
    CascadeMux I__5813 (
            .O(N__34173),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0_cascade_ ));
    InMux I__5812 (
            .O(N__34170),
            .I(N__34163));
    InMux I__5811 (
            .O(N__34169),
            .I(N__34154));
    InMux I__5810 (
            .O(N__34168),
            .I(N__34154));
    InMux I__5809 (
            .O(N__34167),
            .I(N__34154));
    InMux I__5808 (
            .O(N__34166),
            .I(N__34154));
    LocalMux I__5807 (
            .O(N__34163),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6 ));
    LocalMux I__5806 (
            .O(N__34154),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6 ));
    CascadeMux I__5805 (
            .O(N__34149),
            .I(N__34143));
    InMux I__5804 (
            .O(N__34148),
            .I(N__34140));
    InMux I__5803 (
            .O(N__34147),
            .I(N__34137));
    InMux I__5802 (
            .O(N__34146),
            .I(N__34132));
    InMux I__5801 (
            .O(N__34143),
            .I(N__34132));
    LocalMux I__5800 (
            .O(N__34140),
            .I(N__34129));
    LocalMux I__5799 (
            .O(N__34137),
            .I(N__34126));
    LocalMux I__5798 (
            .O(N__34132),
            .I(N__34122));
    Span4Mux_v I__5797 (
            .O(N__34129),
            .I(N__34117));
    Span4Mux_h I__5796 (
            .O(N__34126),
            .I(N__34117));
    CascadeMux I__5795 (
            .O(N__34125),
            .I(N__34113));
    Span4Mux_v I__5794 (
            .O(N__34122),
            .I(N__34110));
    Span4Mux_v I__5793 (
            .O(N__34117),
            .I(N__34107));
    InMux I__5792 (
            .O(N__34116),
            .I(N__34102));
    InMux I__5791 (
            .O(N__34113),
            .I(N__34102));
    Span4Mux_v I__5790 (
            .O(N__34110),
            .I(N__34099));
    Odrv4 I__5789 (
            .O(N__34107),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1 ));
    LocalMux I__5788 (
            .O(N__34102),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1 ));
    Odrv4 I__5787 (
            .O(N__34099),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1 ));
    InMux I__5786 (
            .O(N__34092),
            .I(N__34086));
    InMux I__5785 (
            .O(N__34091),
            .I(N__34086));
    LocalMux I__5784 (
            .O(N__34086),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_1786_2 ));
    InMux I__5783 (
            .O(N__34083),
            .I(N__34080));
    LocalMux I__5782 (
            .O(N__34080),
            .I(N__34077));
    Odrv4 I__5781 (
            .O(N__34077),
            .I(N_979));
    InMux I__5780 (
            .O(N__34074),
            .I(N__34071));
    LocalMux I__5779 (
            .O(N__34071),
            .I(N__34068));
    Span4Mux_h I__5778 (
            .O(N__34068),
            .I(N__34065));
    Odrv4 I__5777 (
            .O(N__34065),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_id_prdata_1_4_u_i_0));
    InMux I__5776 (
            .O(N__34062),
            .I(N__34059));
    LocalMux I__5775 (
            .O(N__34059),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2));
    CascadeMux I__5774 (
            .O(N__34056),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2_cascade_));
    CascadeMux I__5773 (
            .O(N__34053),
            .I(N_1838_0_cascade_));
    InMux I__5772 (
            .O(N__34050),
            .I(N__34046));
    InMux I__5771 (
            .O(N__34049),
            .I(N__34043));
    LocalMux I__5770 (
            .O(N__34046),
            .I(N__34040));
    LocalMux I__5769 (
            .O(N__34043),
            .I(N__34037));
    Span4Mux_h I__5768 (
            .O(N__34040),
            .I(N__34034));
    Span4Mux_h I__5767 (
            .O(N__34037),
            .I(N__34031));
    Odrv4 I__5766 (
            .O(N__34034),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable));
    Odrv4 I__5765 (
            .O(N__34031),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable));
    InMux I__5764 (
            .O(N__34026),
            .I(N__34023));
    LocalMux I__5763 (
            .O(N__34023),
            .I(N__34020));
    Span4Mux_v I__5762 (
            .O(N__34020),
            .I(N__34017));
    Span4Mux_h I__5761 (
            .O(N__34017),
            .I(N__34014));
    Odrv4 I__5760 (
            .O(N__34014),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_30));
    CascadeMux I__5759 (
            .O(N__34011),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1654_cascade_ ));
    CascadeMux I__5758 (
            .O(N__34008),
            .I(N_12_0_cascade_));
    InMux I__5757 (
            .O(N__34005),
            .I(N__34002));
    LocalMux I__5756 (
            .O(N__34002),
            .I(N__33998));
    InMux I__5755 (
            .O(N__34001),
            .I(N__33995));
    Span4Mux_h I__5754 (
            .O(N__33998),
            .I(N__33991));
    LocalMux I__5753 (
            .O(N__33995),
            .I(N__33988));
    InMux I__5752 (
            .O(N__33994),
            .I(N__33985));
    Span4Mux_v I__5751 (
            .O(N__33991),
            .I(N__33980));
    Span4Mux_h I__5750 (
            .O(N__33988),
            .I(N__33980));
    LocalMux I__5749 (
            .O(N__33985),
            .I(N__33977));
    Span4Mux_v I__5748 (
            .O(N__33980),
            .I(N__33971));
    Span4Mux_h I__5747 (
            .O(N__33977),
            .I(N__33971));
    InMux I__5746 (
            .O(N__33976),
            .I(N__33968));
    Span4Mux_v I__5745 (
            .O(N__33971),
            .I(N__33965));
    LocalMux I__5744 (
            .O(N__33968),
            .I(N__33962));
    Span4Mux_h I__5743 (
            .O(N__33965),
            .I(N__33959));
    Span12Mux_h I__5742 (
            .O(N__33962),
            .I(N__33956));
    Odrv4 I__5741 (
            .O(N__33959),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7 ));
    Odrv12 I__5740 (
            .O(N__33956),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7 ));
    InMux I__5739 (
            .O(N__33951),
            .I(N__33926));
    CascadeMux I__5738 (
            .O(N__33950),
            .I(N__33923));
    InMux I__5737 (
            .O(N__33949),
            .I(N__33901));
    InMux I__5736 (
            .O(N__33948),
            .I(N__33901));
    InMux I__5735 (
            .O(N__33947),
            .I(N__33901));
    InMux I__5734 (
            .O(N__33946),
            .I(N__33901));
    InMux I__5733 (
            .O(N__33945),
            .I(N__33901));
    InMux I__5732 (
            .O(N__33944),
            .I(N__33901));
    InMux I__5731 (
            .O(N__33943),
            .I(N__33901));
    InMux I__5730 (
            .O(N__33942),
            .I(N__33886));
    InMux I__5729 (
            .O(N__33941),
            .I(N__33886));
    InMux I__5728 (
            .O(N__33940),
            .I(N__33886));
    InMux I__5727 (
            .O(N__33939),
            .I(N__33886));
    InMux I__5726 (
            .O(N__33938),
            .I(N__33886));
    InMux I__5725 (
            .O(N__33937),
            .I(N__33886));
    InMux I__5724 (
            .O(N__33936),
            .I(N__33886));
    InMux I__5723 (
            .O(N__33935),
            .I(N__33871));
    InMux I__5722 (
            .O(N__33934),
            .I(N__33871));
    InMux I__5721 (
            .O(N__33933),
            .I(N__33871));
    InMux I__5720 (
            .O(N__33932),
            .I(N__33871));
    InMux I__5719 (
            .O(N__33931),
            .I(N__33871));
    InMux I__5718 (
            .O(N__33930),
            .I(N__33871));
    InMux I__5717 (
            .O(N__33929),
            .I(N__33871));
    LocalMux I__5716 (
            .O(N__33926),
            .I(N__33868));
    InMux I__5715 (
            .O(N__33923),
            .I(N__33865));
    InMux I__5714 (
            .O(N__33922),
            .I(N__33862));
    InMux I__5713 (
            .O(N__33921),
            .I(N__33849));
    InMux I__5712 (
            .O(N__33920),
            .I(N__33849));
    InMux I__5711 (
            .O(N__33919),
            .I(N__33849));
    InMux I__5710 (
            .O(N__33918),
            .I(N__33849));
    InMux I__5709 (
            .O(N__33917),
            .I(N__33849));
    InMux I__5708 (
            .O(N__33916),
            .I(N__33849));
    LocalMux I__5707 (
            .O(N__33901),
            .I(N__33846));
    LocalMux I__5706 (
            .O(N__33886),
            .I(N__33841));
    LocalMux I__5705 (
            .O(N__33871),
            .I(N__33841));
    Span12Mux_h I__5704 (
            .O(N__33868),
            .I(N__33838));
    LocalMux I__5703 (
            .O(N__33865),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ));
    LocalMux I__5702 (
            .O(N__33862),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ));
    LocalMux I__5701 (
            .O(N__33849),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ));
    Odrv4 I__5700 (
            .O(N__33846),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ));
    Odrv12 I__5699 (
            .O(N__33841),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ));
    Odrv12 I__5698 (
            .O(N__33838),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ));
    InMux I__5697 (
            .O(N__33825),
            .I(N__33822));
    LocalMux I__5696 (
            .O(N__33822),
            .I(N__33818));
    InMux I__5695 (
            .O(N__33821),
            .I(N__33815));
    Span4Mux_v I__5694 (
            .O(N__33818),
            .I(N__33812));
    LocalMux I__5693 (
            .O(N__33815),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_7));
    Odrv4 I__5692 (
            .O(N__33812),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_7));
    CascadeMux I__5691 (
            .O(N__33807),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0_cascade_ ));
    InMux I__5690 (
            .O(N__33804),
            .I(N__33801));
    LocalMux I__5689 (
            .O(N__33801),
            .I(N_12_0));
    InMux I__5688 (
            .O(N__33798),
            .I(N__33795));
    LocalMux I__5687 (
            .O(N__33795),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_0_7 ));
    CascadeMux I__5686 (
            .O(N__33792),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_23_cascade_ ));
    CascadeMux I__5685 (
            .O(N__33789),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDDZ0Z7_cascade_ ));
    CascadeMux I__5684 (
            .O(N__33786),
            .I(N__33783));
    InMux I__5683 (
            .O(N__33783),
            .I(N__33780));
    LocalMux I__5682 (
            .O(N__33780),
            .I(N__33776));
    InMux I__5681 (
            .O(N__33779),
            .I(N__33772));
    Span4Mux_h I__5680 (
            .O(N__33776),
            .I(N__33769));
    InMux I__5679 (
            .O(N__33775),
            .I(N__33766));
    LocalMux I__5678 (
            .O(N__33772),
            .I(N__33761));
    Span4Mux_h I__5677 (
            .O(N__33769),
            .I(N__33761));
    LocalMux I__5676 (
            .O(N__33766),
            .I(N__33758));
    Span4Mux_v I__5675 (
            .O(N__33761),
            .I(N__33755));
    Span12Mux_h I__5674 (
            .O(N__33758),
            .I(N__33752));
    Odrv4 I__5673 (
            .O(N__33755),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_6));
    Odrv12 I__5672 (
            .O(N__33752),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_6));
    InMux I__5671 (
            .O(N__33747),
            .I(N__33744));
    LocalMux I__5670 (
            .O(N__33744),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_6 ));
    InMux I__5669 (
            .O(N__33741),
            .I(N__33738));
    LocalMux I__5668 (
            .O(N__33738),
            .I(N__33734));
    CascadeMux I__5667 (
            .O(N__33737),
            .I(N__33731));
    Span4Mux_h I__5666 (
            .O(N__33734),
            .I(N__33727));
    InMux I__5665 (
            .O(N__33731),
            .I(N__33722));
    InMux I__5664 (
            .O(N__33730),
            .I(N__33722));
    Span4Mux_v I__5663 (
            .O(N__33727),
            .I(N__33717));
    LocalMux I__5662 (
            .O(N__33722),
            .I(N__33717));
    Odrv4 I__5661 (
            .O(N__33717),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_3));
    CascadeMux I__5660 (
            .O(N__33714),
            .I(N__33711));
    InMux I__5659 (
            .O(N__33711),
            .I(N__33707));
    InMux I__5658 (
            .O(N__33710),
            .I(N__33704));
    LocalMux I__5657 (
            .O(N__33707),
            .I(N__33700));
    LocalMux I__5656 (
            .O(N__33704),
            .I(N__33697));
    InMux I__5655 (
            .O(N__33703),
            .I(N__33694));
    Span4Mux_v I__5654 (
            .O(N__33700),
            .I(N__33691));
    Span4Mux_h I__5653 (
            .O(N__33697),
            .I(N__33688));
    LocalMux I__5652 (
            .O(N__33694),
            .I(N__33683));
    Sp12to4 I__5651 (
            .O(N__33691),
            .I(N__33683));
    Odrv4 I__5650 (
            .O(N__33688),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_4));
    Odrv12 I__5649 (
            .O(N__33683),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_4));
    InMux I__5648 (
            .O(N__33678),
            .I(N__33675));
    LocalMux I__5647 (
            .O(N__33675),
            .I(N__33670));
    InMux I__5646 (
            .O(N__33674),
            .I(N__33665));
    InMux I__5645 (
            .O(N__33673),
            .I(N__33665));
    Span4Mux_h I__5644 (
            .O(N__33670),
            .I(N__33662));
    LocalMux I__5643 (
            .O(N__33665),
            .I(N__33659));
    Odrv4 I__5642 (
            .O(N__33662),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_6));
    Odrv4 I__5641 (
            .O(N__33659),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_6));
    InMux I__5640 (
            .O(N__33654),
            .I(N__33651));
    LocalMux I__5639 (
            .O(N__33651),
            .I(N__33648));
    Span4Mux_h I__5638 (
            .O(N__33648),
            .I(N__33645));
    Span4Mux_h I__5637 (
            .O(N__33645),
            .I(N__33642));
    Odrv4 I__5636 (
            .O(N__33642),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_0Z0Z_26 ));
    CascadeMux I__5635 (
            .O(N__33639),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGHZ0Z5_cascade_ ));
    InMux I__5634 (
            .O(N__33636),
            .I(N__33630));
    InMux I__5633 (
            .O(N__33635),
            .I(N__33630));
    LocalMux I__5632 (
            .O(N__33630),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_15 ));
    InMux I__5631 (
            .O(N__33627),
            .I(N__33624));
    LocalMux I__5630 (
            .O(N__33624),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14 ));
    InMux I__5629 (
            .O(N__33621),
            .I(N__33618));
    LocalMux I__5628 (
            .O(N__33618),
            .I(N__33615));
    Span4Mux_h I__5627 (
            .O(N__33615),
            .I(N__33612));
    Sp12to4 I__5626 (
            .O(N__33612),
            .I(N__33609));
    Span12Mux_h I__5625 (
            .O(N__33609),
            .I(N__33606));
    Odrv12 I__5624 (
            .O(N__33606),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_13 ));
    CascadeMux I__5623 (
            .O(N__33603),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14_cascade_ ));
    CascadeMux I__5622 (
            .O(N__33600),
            .I(N__33597));
    InMux I__5621 (
            .O(N__33597),
            .I(N__33594));
    LocalMux I__5620 (
            .O(N__33594),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_14 ));
    CascadeMux I__5619 (
            .O(N__33591),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_14_cascade_ ));
    InMux I__5618 (
            .O(N__33588),
            .I(N__33585));
    LocalMux I__5617 (
            .O(N__33585),
            .I(N__33582));
    Odrv4 I__5616 (
            .O(N__33582),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_14 ));
    InMux I__5615 (
            .O(N__33579),
            .I(N__33576));
    LocalMux I__5614 (
            .O(N__33576),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGHZ0Z5 ));
    CascadeMux I__5613 (
            .O(N__33573),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_14_cascade_ ));
    InMux I__5612 (
            .O(N__33570),
            .I(N__33567));
    LocalMux I__5611 (
            .O(N__33567),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_14 ));
    InMux I__5610 (
            .O(N__33564),
            .I(N__33561));
    LocalMux I__5609 (
            .O(N__33561),
            .I(N__33558));
    Span4Mux_v I__5608 (
            .O(N__33558),
            .I(N__33553));
    InMux I__5607 (
            .O(N__33557),
            .I(N__33550));
    InMux I__5606 (
            .O(N__33556),
            .I(N__33547));
    Odrv4 I__5605 (
            .O(N__33553),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_14));
    LocalMux I__5604 (
            .O(N__33550),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_14));
    LocalMux I__5603 (
            .O(N__33547),
            .I(cemf_module_64ch_ctrl_inst1_data_coarseovf_14));
    InMux I__5602 (
            .O(N__33540),
            .I(N__33537));
    LocalMux I__5601 (
            .O(N__33537),
            .I(N__33534));
    Span4Mux_v I__5600 (
            .O(N__33534),
            .I(N__33531));
    Span4Mux_h I__5599 (
            .O(N__33531),
            .I(N__33528));
    Odrv4 I__5598 (
            .O(N__33528),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_1 ));
    InMux I__5597 (
            .O(N__33525),
            .I(N__33522));
    LocalMux I__5596 (
            .O(N__33522),
            .I(N__33518));
    CascadeMux I__5595 (
            .O(N__33521),
            .I(N__33515));
    Span4Mux_v I__5594 (
            .O(N__33518),
            .I(N__33512));
    InMux I__5593 (
            .O(N__33515),
            .I(N__33509));
    Span4Mux_h I__5592 (
            .O(N__33512),
            .I(N__33506));
    LocalMux I__5591 (
            .O(N__33509),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_18));
    Odrv4 I__5590 (
            .O(N__33506),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_18));
    CascadeMux I__5589 (
            .O(N__33501),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0_cascade_ ));
    InMux I__5588 (
            .O(N__33498),
            .I(N__33495));
    LocalMux I__5587 (
            .O(N__33495),
            .I(N__33492));
    Span4Mux_h I__5586 (
            .O(N__33492),
            .I(N__33489));
    Odrv4 I__5585 (
            .O(N__33489),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_18 ));
    CascadeMux I__5584 (
            .O(N__33486),
            .I(N__33483));
    InMux I__5583 (
            .O(N__33483),
            .I(N__33480));
    LocalMux I__5582 (
            .O(N__33480),
            .I(N__33476));
    InMux I__5581 (
            .O(N__33479),
            .I(N__33473));
    Span4Mux_v I__5580 (
            .O(N__33476),
            .I(N__33470));
    LocalMux I__5579 (
            .O(N__33473),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_20));
    Odrv4 I__5578 (
            .O(N__33470),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_20));
    InMux I__5577 (
            .O(N__33465),
            .I(N__33462));
    LocalMux I__5576 (
            .O(N__33462),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_20 ));
    CascadeMux I__5575 (
            .O(N__33459),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0_cascade_ ));
    InMux I__5574 (
            .O(N__33456),
            .I(N__33453));
    LocalMux I__5573 (
            .O(N__33453),
            .I(N__33450));
    Span4Mux_v I__5572 (
            .O(N__33450),
            .I(N__33447));
    Sp12to4 I__5571 (
            .O(N__33447),
            .I(N__33444));
    Odrv12 I__5570 (
            .O(N__33444),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_7 ));
    CascadeMux I__5569 (
            .O(N__33441),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_15_cascade_ ));
    InMux I__5568 (
            .O(N__33438),
            .I(N__33435));
    LocalMux I__5567 (
            .O(N__33435),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_19 ));
    InMux I__5566 (
            .O(N__33432),
            .I(N__33428));
    InMux I__5565 (
            .O(N__33431),
            .I(N__33425));
    LocalMux I__5564 (
            .O(N__33428),
            .I(N__33422));
    LocalMux I__5563 (
            .O(N__33425),
            .I(N__33419));
    Span12Mux_v I__5562 (
            .O(N__33422),
            .I(N__33416));
    Span12Mux_v I__5561 (
            .O(N__33419),
            .I(N__33413));
    Odrv12 I__5560 (
            .O(N__33416),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable));
    Odrv12 I__5559 (
            .O(N__33413),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable));
    InMux I__5558 (
            .O(N__33408),
            .I(N__33405));
    LocalMux I__5557 (
            .O(N__33405),
            .I(N__33402));
    Span4Mux_v I__5556 (
            .O(N__33402),
            .I(N__33399));
    Sp12to4 I__5555 (
            .O(N__33399),
            .I(N__33396));
    Odrv12 I__5554 (
            .O(N__33396),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_0));
    InMux I__5553 (
            .O(N__33393),
            .I(N__33390));
    LocalMux I__5552 (
            .O(N__33390),
            .I(N__33387));
    Span4Mux_v I__5551 (
            .O(N__33387),
            .I(N__33384));
    Span4Mux_v I__5550 (
            .O(N__33384),
            .I(N__33381));
    Sp12to4 I__5549 (
            .O(N__33381),
            .I(N__33378));
    Odrv12 I__5548 (
            .O(N__33378),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_0));
    CascadeMux I__5547 (
            .O(N__33375),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319_cascade_ ));
    CascadeMux I__5546 (
            .O(N__33372),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_0_cascade_ ));
    CascadeMux I__5545 (
            .O(N__33369),
            .I(N__33366));
    InMux I__5544 (
            .O(N__33366),
            .I(N__33362));
    CascadeMux I__5543 (
            .O(N__33365),
            .I(N__33359));
    LocalMux I__5542 (
            .O(N__33362),
            .I(N__33356));
    InMux I__5541 (
            .O(N__33359),
            .I(N__33353));
    Span4Mux_h I__5540 (
            .O(N__33356),
            .I(N__33350));
    LocalMux I__5539 (
            .O(N__33353),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_21));
    Odrv4 I__5538 (
            .O(N__33350),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_21));
    CascadeMux I__5537 (
            .O(N__33345),
            .I(N__33342));
    InMux I__5536 (
            .O(N__33342),
            .I(N__33339));
    LocalMux I__5535 (
            .O(N__33339),
            .I(N__33336));
    Span4Mux_h I__5534 (
            .O(N__33336),
            .I(N__33333));
    Span4Mux_v I__5533 (
            .O(N__33333),
            .I(N__33330));
    Span4Mux_h I__5532 (
            .O(N__33330),
            .I(N__33327));
    Odrv4 I__5531 (
            .O(N__33327),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_22));
    CascadeMux I__5530 (
            .O(N__33324),
            .I(N__33321));
    InMux I__5529 (
            .O(N__33321),
            .I(N__33318));
    LocalMux I__5528 (
            .O(N__33318),
            .I(N__33315));
    Odrv4 I__5527 (
            .O(N__33315),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_698 ));
    InMux I__5526 (
            .O(N__33312),
            .I(N__33309));
    LocalMux I__5525 (
            .O(N__33309),
            .I(N__33306));
    Sp12to4 I__5524 (
            .O(N__33306),
            .I(N__33303));
    Span12Mux_s11_v I__5523 (
            .O(N__33303),
            .I(N__33300));
    Odrv12 I__5522 (
            .O(N__33300),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_23));
    InMux I__5521 (
            .O(N__33297),
            .I(N__33294));
    LocalMux I__5520 (
            .O(N__33294),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_2 ));
    InMux I__5519 (
            .O(N__33291),
            .I(N__33288));
    LocalMux I__5518 (
            .O(N__33288),
            .I(N__33285));
    Span4Mux_h I__5517 (
            .O(N__33285),
            .I(N__33282));
    Span4Mux_h I__5516 (
            .O(N__33282),
            .I(N__33279));
    Span4Mux_h I__5515 (
            .O(N__33279),
            .I(N__33276));
    Odrv4 I__5514 (
            .O(N__33276),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_25));
    CascadeMux I__5513 (
            .O(N__33273),
            .I(N__33270));
    InMux I__5512 (
            .O(N__33270),
            .I(N__33267));
    LocalMux I__5511 (
            .O(N__33267),
            .I(N__33264));
    Span4Mux_v I__5510 (
            .O(N__33264),
            .I(N__33261));
    Span4Mux_h I__5509 (
            .O(N__33261),
            .I(N__33258));
    Odrv4 I__5508 (
            .O(N__33258),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_27));
    InMux I__5507 (
            .O(N__33255),
            .I(N__33252));
    LocalMux I__5506 (
            .O(N__33252),
            .I(N__33249));
    Span4Mux_v I__5505 (
            .O(N__33249),
            .I(N__33246));
    Span4Mux_h I__5504 (
            .O(N__33246),
            .I(N__33243));
    Span4Mux_h I__5503 (
            .O(N__33243),
            .I(N__33240));
    Odrv4 I__5502 (
            .O(N__33240),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_19));
    CascadeMux I__5501 (
            .O(N__33237),
            .I(N__33234));
    InMux I__5500 (
            .O(N__33234),
            .I(N__33231));
    LocalMux I__5499 (
            .O(N__33231),
            .I(N__33228));
    Span4Mux_v I__5498 (
            .O(N__33228),
            .I(N__33225));
    Span4Mux_h I__5497 (
            .O(N__33225),
            .I(N__33222));
    Span4Mux_h I__5496 (
            .O(N__33222),
            .I(N__33219));
    Odrv4 I__5495 (
            .O(N__33219),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_19));
    InMux I__5494 (
            .O(N__33216),
            .I(N__33213));
    LocalMux I__5493 (
            .O(N__33213),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_731 ));
    InMux I__5492 (
            .O(N__33210),
            .I(N__33207));
    LocalMux I__5491 (
            .O(N__33207),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_19 ));
    CascadeMux I__5490 (
            .O(N__33204),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_19_cascade_ ));
    InMux I__5489 (
            .O(N__33201),
            .I(N__33198));
    LocalMux I__5488 (
            .O(N__33198),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_19 ));
    InMux I__5487 (
            .O(N__33195),
            .I(N__33192));
    LocalMux I__5486 (
            .O(N__33192),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_19 ));
    InMux I__5485 (
            .O(N__33189),
            .I(N__33186));
    LocalMux I__5484 (
            .O(N__33186),
            .I(\serializer_mod_inst.shift_regZ0Z_37 ));
    InMux I__5483 (
            .O(N__33183),
            .I(N__33180));
    LocalMux I__5482 (
            .O(N__33180),
            .I(\serializer_mod_inst.shift_regZ0Z_38 ));
    InMux I__5481 (
            .O(N__33177),
            .I(N__33174));
    LocalMux I__5480 (
            .O(N__33174),
            .I(\serializer_mod_inst.shift_regZ0Z_33 ));
    InMux I__5479 (
            .O(N__33171),
            .I(N__33168));
    LocalMux I__5478 (
            .O(N__33168),
            .I(\serializer_mod_inst.shift_regZ0Z_34 ));
    InMux I__5477 (
            .O(N__33165),
            .I(N__33162));
    LocalMux I__5476 (
            .O(N__33162),
            .I(\serializer_mod_inst.shift_regZ0Z_35 ));
    InMux I__5475 (
            .O(N__33159),
            .I(N__33156));
    LocalMux I__5474 (
            .O(N__33156),
            .I(\serializer_mod_inst.shift_regZ0Z_76 ));
    InMux I__5473 (
            .O(N__33153),
            .I(N__33150));
    LocalMux I__5472 (
            .O(N__33150),
            .I(N__33147));
    Span4Mux_h I__5471 (
            .O(N__33147),
            .I(N__33144));
    Span4Mux_v I__5470 (
            .O(N__33144),
            .I(N__33141));
    Sp12to4 I__5469 (
            .O(N__33141),
            .I(N__33138));
    Odrv12 I__5468 (
            .O(N__33138),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_17));
    InMux I__5467 (
            .O(N__33135),
            .I(N__33132));
    LocalMux I__5466 (
            .O(N__33132),
            .I(N__33129));
    Span4Mux_v I__5465 (
            .O(N__33129),
            .I(N__33126));
    Odrv4 I__5464 (
            .O(N__33126),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_753 ));
    CascadeMux I__5463 (
            .O(N__33123),
            .I(N__33120));
    InMux I__5462 (
            .O(N__33120),
            .I(N__33117));
    LocalMux I__5461 (
            .O(N__33117),
            .I(N__33114));
    Span4Mux_h I__5460 (
            .O(N__33114),
            .I(N__33111));
    Span4Mux_v I__5459 (
            .O(N__33111),
            .I(N__33108));
    Span4Mux_h I__5458 (
            .O(N__33108),
            .I(N__33105));
    Odrv4 I__5457 (
            .O(N__33105),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_19));
    InMux I__5456 (
            .O(N__33102),
            .I(N__33099));
    LocalMux I__5455 (
            .O(N__33099),
            .I(N__33096));
    Span4Mux_v I__5454 (
            .O(N__33096),
            .I(N__33093));
    Span4Mux_h I__5453 (
            .O(N__33093),
            .I(N__33090));
    Odrv4 I__5452 (
            .O(N__33090),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_2));
    InMux I__5451 (
            .O(N__33087),
            .I(N__33084));
    LocalMux I__5450 (
            .O(N__33084),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_918 ));
    CascadeMux I__5449 (
            .O(N__33081),
            .I(N__33078));
    InMux I__5448 (
            .O(N__33078),
            .I(N__33075));
    LocalMux I__5447 (
            .O(N__33075),
            .I(N__33072));
    Span4Mux_v I__5446 (
            .O(N__33072),
            .I(N__33069));
    Span4Mux_v I__5445 (
            .O(N__33069),
            .I(N__33066));
    Span4Mux_h I__5444 (
            .O(N__33066),
            .I(N__33063));
    Odrv4 I__5443 (
            .O(N__33063),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_4 ));
    InMux I__5442 (
            .O(N__33060),
            .I(N__33057));
    LocalMux I__5441 (
            .O(N__33057),
            .I(N__33054));
    Odrv4 I__5440 (
            .O(N__33054),
            .I(\serializer_mod_inst.shift_regZ0Z_111 ));
    InMux I__5439 (
            .O(N__33051),
            .I(N__33048));
    LocalMux I__5438 (
            .O(N__33048),
            .I(\serializer_mod_inst.shift_regZ0Z_119 ));
    InMux I__5437 (
            .O(N__33045),
            .I(N__33042));
    LocalMux I__5436 (
            .O(N__33042),
            .I(\serializer_mod_inst.shift_regZ0Z_120 ));
    InMux I__5435 (
            .O(N__33039),
            .I(N__33036));
    LocalMux I__5434 (
            .O(N__33036),
            .I(\serializer_mod_inst.shift_regZ0Z_36 ));
    InMux I__5433 (
            .O(N__33033),
            .I(N__33030));
    LocalMux I__5432 (
            .O(N__33030),
            .I(\serializer_mod_inst.shift_regZ0Z_118 ));
    CascadeMux I__5431 (
            .O(N__33027),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_2_cascade_ ));
    InMux I__5430 (
            .O(N__33024),
            .I(N__33021));
    LocalMux I__5429 (
            .O(N__33021),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1950 ));
    CascadeMux I__5428 (
            .O(N__33018),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1949_cascade_ ));
    IoInMux I__5427 (
            .O(N__33015),
            .I(N__33012));
    LocalMux I__5426 (
            .O(N__33012),
            .I(N__33009));
    IoSpan4Mux I__5425 (
            .O(N__33009),
            .I(N__33006));
    Sp12to4 I__5424 (
            .O(N__33006),
            .I(N__33003));
    Span12Mux_h I__5423 (
            .O(N__33003),
            .I(N__33000));
    Odrv12 I__5422 (
            .O(N__33000),
            .I(stop_fpga2_c));
    InMux I__5421 (
            .O(N__32997),
            .I(N__32994));
    LocalMux I__5420 (
            .O(N__32994),
            .I(N__32989));
    InMux I__5419 (
            .O(N__32993),
            .I(N__32986));
    InMux I__5418 (
            .O(N__32992),
            .I(N__32983));
    Span4Mux_v I__5417 (
            .O(N__32989),
            .I(N__32977));
    LocalMux I__5416 (
            .O(N__32986),
            .I(N__32977));
    LocalMux I__5415 (
            .O(N__32983),
            .I(N__32974));
    InMux I__5414 (
            .O(N__32982),
            .I(N__32970));
    Span4Mux_h I__5413 (
            .O(N__32977),
            .I(N__32967));
    Span4Mux_h I__5412 (
            .O(N__32974),
            .I(N__32964));
    InMux I__5411 (
            .O(N__32973),
            .I(N__32961));
    LocalMux I__5410 (
            .O(N__32970),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_b ));
    Odrv4 I__5409 (
            .O(N__32967),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_b ));
    Odrv4 I__5408 (
            .O(N__32964),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_b ));
    LocalMux I__5407 (
            .O(N__32961),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_b ));
    InMux I__5406 (
            .O(N__32952),
            .I(N__32946));
    InMux I__5405 (
            .O(N__32951),
            .I(N__32943));
    InMux I__5404 (
            .O(N__32950),
            .I(N__32938));
    InMux I__5403 (
            .O(N__32949),
            .I(N__32938));
    LocalMux I__5402 (
            .O(N__32946),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847 ));
    LocalMux I__5401 (
            .O(N__32943),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847 ));
    LocalMux I__5400 (
            .O(N__32938),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847 ));
    InMux I__5399 (
            .O(N__32931),
            .I(N__32928));
    LocalMux I__5398 (
            .O(N__32928),
            .I(\serializer_mod_inst.shift_regZ0Z_112 ));
    CascadeMux I__5397 (
            .O(N__32925),
            .I(N__32922));
    InMux I__5396 (
            .O(N__32922),
            .I(N__32919));
    LocalMux I__5395 (
            .O(N__32919),
            .I(N__32916));
    Span4Mux_v I__5394 (
            .O(N__32916),
            .I(N__32913));
    Span4Mux_v I__5393 (
            .O(N__32913),
            .I(N__32910));
    Span4Mux_v I__5392 (
            .O(N__32910),
            .I(N__32907));
    Odrv4 I__5391 (
            .O(N__32907),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_2 ));
    InMux I__5390 (
            .O(N__32904),
            .I(N__32896));
    InMux I__5389 (
            .O(N__32903),
            .I(N__32885));
    InMux I__5388 (
            .O(N__32902),
            .I(N__32885));
    InMux I__5387 (
            .O(N__32901),
            .I(N__32885));
    InMux I__5386 (
            .O(N__32900),
            .I(N__32885));
    InMux I__5385 (
            .O(N__32899),
            .I(N__32885));
    LocalMux I__5384 (
            .O(N__32896),
            .I(N__32878));
    LocalMux I__5383 (
            .O(N__32885),
            .I(N__32878));
    InMux I__5382 (
            .O(N__32884),
            .I(N__32875));
    InMux I__5381 (
            .O(N__32883),
            .I(N__32872));
    Odrv4 I__5380 (
            .O(N__32878),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_a ));
    LocalMux I__5379 (
            .O(N__32875),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_a ));
    LocalMux I__5378 (
            .O(N__32872),
            .I(\cemf_module_64ch_ctrl_inst1.end_conf_a ));
    CascadeMux I__5377 (
            .O(N__32865),
            .I(\cemf_module_64ch_ctrl_inst1.N_1817_0_cascade_ ));
    CascadeMux I__5376 (
            .O(N__32862),
            .I(N__32859));
    InMux I__5375 (
            .O(N__32859),
            .I(N__32852));
    InMux I__5374 (
            .O(N__32858),
            .I(N__32843));
    InMux I__5373 (
            .O(N__32857),
            .I(N__32843));
    InMux I__5372 (
            .O(N__32856),
            .I(N__32843));
    InMux I__5371 (
            .O(N__32855),
            .I(N__32843));
    LocalMux I__5370 (
            .O(N__32852),
            .I(\cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2 ));
    LocalMux I__5369 (
            .O(N__32843),
            .I(\cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2 ));
    InMux I__5368 (
            .O(N__32838),
            .I(N__32835));
    LocalMux I__5367 (
            .O(N__32835),
            .I(N__32832));
    Span4Mux_v I__5366 (
            .O(N__32832),
            .I(N__32829));
    Odrv4 I__5365 (
            .O(N__32829),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2_8 ));
    CascadeMux I__5364 (
            .O(N__32826),
            .I(N__32822));
    InMux I__5363 (
            .O(N__32825),
            .I(N__32819));
    InMux I__5362 (
            .O(N__32822),
            .I(N__32814));
    LocalMux I__5361 (
            .O(N__32819),
            .I(N__32811));
    InMux I__5360 (
            .O(N__32818),
            .I(N__32806));
    InMux I__5359 (
            .O(N__32817),
            .I(N__32806));
    LocalMux I__5358 (
            .O(N__32814),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845 ));
    Odrv4 I__5357 (
            .O(N__32811),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845 ));
    LocalMux I__5356 (
            .O(N__32806),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845 ));
    CascadeMux I__5355 (
            .O(N__32799),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_0_1_cascade_ ));
    InMux I__5354 (
            .O(N__32796),
            .I(N__32793));
    LocalMux I__5353 (
            .O(N__32793),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1873_0 ));
    InMux I__5352 (
            .O(N__32790),
            .I(N__32787));
    LocalMux I__5351 (
            .O(N__32787),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1874_0 ));
    InMux I__5350 (
            .O(N__32784),
            .I(N__32777));
    InMux I__5349 (
            .O(N__32783),
            .I(N__32777));
    InMux I__5348 (
            .O(N__32782),
            .I(N__32774));
    LocalMux I__5347 (
            .O(N__32777),
            .I(N__32771));
    LocalMux I__5346 (
            .O(N__32774),
            .I(N__32767));
    Span4Mux_v I__5345 (
            .O(N__32771),
            .I(N__32764));
    InMux I__5344 (
            .O(N__32770),
            .I(N__32761));
    Span4Mux_v I__5343 (
            .O(N__32767),
            .I(N__32758));
    Odrv4 I__5342 (
            .O(N__32764),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0 ));
    LocalMux I__5341 (
            .O(N__32761),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0 ));
    Odrv4 I__5340 (
            .O(N__32758),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0 ));
    InMux I__5339 (
            .O(N__32751),
            .I(N__32745));
    InMux I__5338 (
            .O(N__32750),
            .I(N__32745));
    LocalMux I__5337 (
            .O(N__32745),
            .I(N__32740));
    ClkMux I__5336 (
            .O(N__32744),
            .I(N__32733));
    ClkMux I__5335 (
            .O(N__32743),
            .I(N__32733));
    Glb2LocalMux I__5334 (
            .O(N__32740),
            .I(N__32733));
    GlobalMux I__5333 (
            .O(N__32733),
            .I(N__32730));
    gio2CtrlBuf I__5332 (
            .O(N__32730),
            .I(s_sda_i_g));
    InMux I__5331 (
            .O(N__32727),
            .I(N__32724));
    LocalMux I__5330 (
            .O(N__32724),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1392 ));
    CascadeMux I__5329 (
            .O(N__32721),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1381_0_cascade_ ));
    CascadeMux I__5328 (
            .O(N__32718),
            .I(N__32715));
    InMux I__5327 (
            .O(N__32715),
            .I(N__32712));
    LocalMux I__5326 (
            .O(N__32712),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392 ));
    InMux I__5325 (
            .O(N__32709),
            .I(N__32706));
    LocalMux I__5324 (
            .O(N__32706),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_i_2_2 ));
    CascadeMux I__5323 (
            .O(N__32703),
            .I(N__32699));
    InMux I__5322 (
            .O(N__32702),
            .I(N__32693));
    InMux I__5321 (
            .O(N__32699),
            .I(N__32688));
    InMux I__5320 (
            .O(N__32698),
            .I(N__32688));
    InMux I__5319 (
            .O(N__32697),
            .I(N__32685));
    InMux I__5318 (
            .O(N__32696),
            .I(N__32682));
    LocalMux I__5317 (
            .O(N__32693),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16 ));
    LocalMux I__5316 (
            .O(N__32688),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16 ));
    LocalMux I__5315 (
            .O(N__32685),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16 ));
    LocalMux I__5314 (
            .O(N__32682),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16 ));
    InMux I__5313 (
            .O(N__32673),
            .I(N__32668));
    InMux I__5312 (
            .O(N__32672),
            .I(N__32661));
    InMux I__5311 (
            .O(N__32671),
            .I(N__32661));
    LocalMux I__5310 (
            .O(N__32668),
            .I(N__32658));
    InMux I__5309 (
            .O(N__32667),
            .I(N__32653));
    InMux I__5308 (
            .O(N__32666),
            .I(N__32653));
    LocalMux I__5307 (
            .O(N__32661),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17 ));
    Odrv4 I__5306 (
            .O(N__32658),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17 ));
    LocalMux I__5305 (
            .O(N__32653),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17 ));
    InMux I__5304 (
            .O(N__32646),
            .I(N__32643));
    LocalMux I__5303 (
            .O(N__32643),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_18 ));
    CascadeMux I__5302 (
            .O(N__32640),
            .I(N__32637));
    InMux I__5301 (
            .O(N__32637),
            .I(N__32626));
    InMux I__5300 (
            .O(N__32636),
            .I(N__32626));
    InMux I__5299 (
            .O(N__32635),
            .I(N__32621));
    InMux I__5298 (
            .O(N__32634),
            .I(N__32621));
    InMux I__5297 (
            .O(N__32633),
            .I(N__32618));
    InMux I__5296 (
            .O(N__32632),
            .I(N__32613));
    InMux I__5295 (
            .O(N__32631),
            .I(N__32613));
    LocalMux I__5294 (
            .O(N__32626),
            .I(N__32606));
    LocalMux I__5293 (
            .O(N__32621),
            .I(N__32606));
    LocalMux I__5292 (
            .O(N__32618),
            .I(N__32606));
    LocalMux I__5291 (
            .O(N__32613),
            .I(N__32603));
    Span4Mux_v I__5290 (
            .O(N__32606),
            .I(N__32599));
    Span4Mux_v I__5289 (
            .O(N__32603),
            .I(N__32596));
    InMux I__5288 (
            .O(N__32602),
            .I(N__32593));
    Span4Mux_h I__5287 (
            .O(N__32599),
            .I(N__32588));
    Span4Mux_h I__5286 (
            .O(N__32596),
            .I(N__32585));
    LocalMux I__5285 (
            .O(N__32593),
            .I(N__32582));
    InMux I__5284 (
            .O(N__32592),
            .I(N__32577));
    InMux I__5283 (
            .O(N__32591),
            .I(N__32577));
    Odrv4 I__5282 (
            .O(N__32588),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0 ));
    Odrv4 I__5281 (
            .O(N__32585),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0 ));
    Odrv4 I__5280 (
            .O(N__32582),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0 ));
    LocalMux I__5279 (
            .O(N__32577),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0 ));
    InMux I__5278 (
            .O(N__32568),
            .I(N__32561));
    InMux I__5277 (
            .O(N__32567),
            .I(N__32561));
    InMux I__5276 (
            .O(N__32566),
            .I(N__32558));
    LocalMux I__5275 (
            .O(N__32561),
            .I(N__32552));
    LocalMux I__5274 (
            .O(N__32558),
            .I(N__32552));
    InMux I__5273 (
            .O(N__32557),
            .I(N__32549));
    Span4Mux_v I__5272 (
            .O(N__32552),
            .I(N__32546));
    LocalMux I__5271 (
            .O(N__32549),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1 ));
    Odrv4 I__5270 (
            .O(N__32546),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1 ));
    InMux I__5269 (
            .O(N__32541),
            .I(N__32529));
    InMux I__5268 (
            .O(N__32540),
            .I(N__32529));
    InMux I__5267 (
            .O(N__32539),
            .I(N__32529));
    InMux I__5266 (
            .O(N__32538),
            .I(N__32529));
    LocalMux I__5265 (
            .O(N__32529),
            .I(N__32526));
    Span4Mux_v I__5264 (
            .O(N__32526),
            .I(N__32523));
    Odrv4 I__5263 (
            .O(N__32523),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_11_0_i_0_1 ));
    CascadeMux I__5262 (
            .O(N__32520),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_1394_cascade_ ));
    CEMux I__5261 (
            .O(N__32517),
            .I(N__32513));
    CEMux I__5260 (
            .O(N__32516),
            .I(N__32509));
    LocalMux I__5259 (
            .O(N__32513),
            .I(N__32506));
    CEMux I__5258 (
            .O(N__32512),
            .I(N__32503));
    LocalMux I__5257 (
            .O(N__32509),
            .I(N__32500));
    Span4Mux_v I__5256 (
            .O(N__32506),
            .I(N__32497));
    LocalMux I__5255 (
            .O(N__32503),
            .I(N__32494));
    Span4Mux_h I__5254 (
            .O(N__32500),
            .I(N__32491));
    Sp12to4 I__5253 (
            .O(N__32497),
            .I(N__32485));
    Span4Mux_v I__5252 (
            .O(N__32494),
            .I(N__32482));
    Span4Mux_h I__5251 (
            .O(N__32491),
            .I(N__32479));
    CEMux I__5250 (
            .O(N__32490),
            .I(N__32476));
    CEMux I__5249 (
            .O(N__32489),
            .I(N__32473));
    CEMux I__5248 (
            .O(N__32488),
            .I(N__32470));
    Span12Mux_h I__5247 (
            .O(N__32485),
            .I(N__32465));
    Sp12to4 I__5246 (
            .O(N__32482),
            .I(N__32465));
    Span4Mux_v I__5245 (
            .O(N__32479),
            .I(N__32462));
    LocalMux I__5244 (
            .O(N__32476),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ));
    LocalMux I__5243 (
            .O(N__32473),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ));
    LocalMux I__5242 (
            .O(N__32470),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ));
    Odrv12 I__5241 (
            .O(N__32465),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ));
    Odrv4 I__5240 (
            .O(N__32462),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ));
    InMux I__5239 (
            .O(N__32451),
            .I(N__32448));
    LocalMux I__5238 (
            .O(N__32448),
            .I(N__32445));
    Span4Mux_h I__5237 (
            .O(N__32445),
            .I(N__32442));
    Span4Mux_h I__5236 (
            .O(N__32442),
            .I(N__32439));
    Span4Mux_v I__5235 (
            .O(N__32439),
            .I(N__32436));
    Odrv4 I__5234 (
            .O(N__32436),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_16));
    CascadeMux I__5233 (
            .O(N__32433),
            .I(N__32430));
    InMux I__5232 (
            .O(N__32430),
            .I(N__32427));
    LocalMux I__5231 (
            .O(N__32427),
            .I(N__32424));
    Span4Mux_v I__5230 (
            .O(N__32424),
            .I(N__32421));
    Span4Mux_h I__5229 (
            .O(N__32421),
            .I(N__32418));
    Span4Mux_h I__5228 (
            .O(N__32418),
            .I(N__32415));
    Odrv4 I__5227 (
            .O(N__32415),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_18));
    InMux I__5226 (
            .O(N__32412),
            .I(N__32409));
    LocalMux I__5225 (
            .O(N__32409),
            .I(N__32406));
    Span4Mux_v I__5224 (
            .O(N__32406),
            .I(N__32403));
    Odrv4 I__5223 (
            .O(N__32403),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1911 ));
    InMux I__5222 (
            .O(N__32400),
            .I(N__32397));
    LocalMux I__5221 (
            .O(N__32397),
            .I(N__32394));
    Span4Mux_v I__5220 (
            .O(N__32394),
            .I(N__32391));
    Span4Mux_h I__5219 (
            .O(N__32391),
            .I(N__32388));
    Odrv4 I__5218 (
            .O(N__32388),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_8));
    CascadeMux I__5217 (
            .O(N__32385),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0_cascade_ ));
    InMux I__5216 (
            .O(N__32382),
            .I(N__32379));
    LocalMux I__5215 (
            .O(N__32379),
            .I(N__32376));
    Span4Mux_h I__5214 (
            .O(N__32376),
            .I(N__32373));
    Span4Mux_v I__5213 (
            .O(N__32373),
            .I(N__32370));
    Span4Mux_v I__5212 (
            .O(N__32370),
            .I(N__32367));
    Odrv4 I__5211 (
            .O(N__32367),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1920 ));
    InMux I__5210 (
            .O(N__32364),
            .I(N__32357));
    InMux I__5209 (
            .O(N__32363),
            .I(N__32350));
    InMux I__5208 (
            .O(N__32362),
            .I(N__32350));
    InMux I__5207 (
            .O(N__32361),
            .I(N__32350));
    InMux I__5206 (
            .O(N__32360),
            .I(N__32347));
    LocalMux I__5205 (
            .O(N__32357),
            .I(N__32344));
    LocalMux I__5204 (
            .O(N__32350),
            .I(N__32341));
    LocalMux I__5203 (
            .O(N__32347),
            .I(N__32338));
    Span4Mux_h I__5202 (
            .O(N__32344),
            .I(N__32331));
    Span4Mux_h I__5201 (
            .O(N__32341),
            .I(N__32331));
    Span4Mux_h I__5200 (
            .O(N__32338),
            .I(N__32328));
    InMux I__5199 (
            .O(N__32337),
            .I(N__32323));
    InMux I__5198 (
            .O(N__32336),
            .I(N__32323));
    Span4Mux_v I__5197 (
            .O(N__32331),
            .I(N__32320));
    Odrv4 I__5196 (
            .O(N__32328),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable));
    LocalMux I__5195 (
            .O(N__32323),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable));
    Odrv4 I__5194 (
            .O(N__32320),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable));
    InMux I__5193 (
            .O(N__32313),
            .I(N__32306));
    InMux I__5192 (
            .O(N__32312),
            .I(N__32306));
    InMux I__5191 (
            .O(N__32311),
            .I(N__32303));
    LocalMux I__5190 (
            .O(N__32306),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0 ));
    LocalMux I__5189 (
            .O(N__32303),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0 ));
    InMux I__5188 (
            .O(N__32298),
            .I(N__32294));
    InMux I__5187 (
            .O(N__32297),
            .I(N__32291));
    LocalMux I__5186 (
            .O(N__32294),
            .I(N__32288));
    LocalMux I__5185 (
            .O(N__32291),
            .I(N__32285));
    Span4Mux_h I__5184 (
            .O(N__32288),
            .I(N__32280));
    Span4Mux_v I__5183 (
            .O(N__32285),
            .I(N__32280));
    Odrv4 I__5182 (
            .O(N__32280),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m20_0_a2_4_1 ));
    CascadeMux I__5181 (
            .O(N__32277),
            .I(N__32273));
    CascadeMux I__5180 (
            .O(N__32276),
            .I(N__32268));
    InMux I__5179 (
            .O(N__32273),
            .I(N__32265));
    InMux I__5178 (
            .O(N__32272),
            .I(N__32260));
    InMux I__5177 (
            .O(N__32271),
            .I(N__32260));
    InMux I__5176 (
            .O(N__32268),
            .I(N__32257));
    LocalMux I__5175 (
            .O(N__32265),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13 ));
    LocalMux I__5174 (
            .O(N__32260),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13 ));
    LocalMux I__5173 (
            .O(N__32257),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13 ));
    IoInMux I__5172 (
            .O(N__32250),
            .I(N__32247));
    LocalMux I__5171 (
            .O(N__32247),
            .I(N__32244));
    Span4Mux_s2_h I__5170 (
            .O(N__32244),
            .I(N__32241));
    Span4Mux_h I__5169 (
            .O(N__32241),
            .I(N__32238));
    Span4Mux_h I__5168 (
            .O(N__32238),
            .I(N__32235));
    Span4Mux_h I__5167 (
            .O(N__32235),
            .I(N__32232));
    Odrv4 I__5166 (
            .O(N__32232),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa ));
    CascadeMux I__5165 (
            .O(N__32229),
            .I(N__32226));
    InMux I__5164 (
            .O(N__32226),
            .I(N__32223));
    LocalMux I__5163 (
            .O(N__32223),
            .I(N__32219));
    InMux I__5162 (
            .O(N__32222),
            .I(N__32216));
    Span12Mux_h I__5161 (
            .O(N__32219),
            .I(N__32213));
    LocalMux I__5160 (
            .O(N__32216),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_5));
    Odrv12 I__5159 (
            .O(N__32213),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_5));
    CascadeMux I__5158 (
            .O(N__32208),
            .I(N__32204));
    InMux I__5157 (
            .O(N__32207),
            .I(N__32201));
    InMux I__5156 (
            .O(N__32204),
            .I(N__32198));
    LocalMux I__5155 (
            .O(N__32201),
            .I(N__32194));
    LocalMux I__5154 (
            .O(N__32198),
            .I(N__32191));
    InMux I__5153 (
            .O(N__32197),
            .I(N__32188));
    Span4Mux_v I__5152 (
            .O(N__32194),
            .I(N__32185));
    Span12Mux_v I__5151 (
            .O(N__32191),
            .I(N__32182));
    LocalMux I__5150 (
            .O(N__32188),
            .I(N__32177));
    Span4Mux_h I__5149 (
            .O(N__32185),
            .I(N__32177));
    Odrv12 I__5148 (
            .O(N__32182),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_5));
    Odrv4 I__5147 (
            .O(N__32177),
            .I(cemf_module_64ch_ctrl_inst1_data_interrupts_5));
    CascadeMux I__5146 (
            .O(N__32172),
            .I(N__32167));
    InMux I__5145 (
            .O(N__32171),
            .I(N__32164));
    InMux I__5144 (
            .O(N__32170),
            .I(N__32161));
    InMux I__5143 (
            .O(N__32167),
            .I(N__32158));
    LocalMux I__5142 (
            .O(N__32164),
            .I(N__32155));
    LocalMux I__5141 (
            .O(N__32161),
            .I(N__32152));
    LocalMux I__5140 (
            .O(N__32158),
            .I(N__32149));
    Odrv12 I__5139 (
            .O(N__32155),
            .I(cemf_module_64ch_ctrl_inst1_data_config_5));
    Odrv4 I__5138 (
            .O(N__32152),
            .I(cemf_module_64ch_ctrl_inst1_data_config_5));
    Odrv4 I__5137 (
            .O(N__32149),
            .I(cemf_module_64ch_ctrl_inst1_data_config_5));
    CascadeMux I__5136 (
            .O(N__32142),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_5_cascade_ ));
    InMux I__5135 (
            .O(N__32139),
            .I(N__32136));
    LocalMux I__5134 (
            .O(N__32136),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRLZ0Z7 ));
    InMux I__5133 (
            .O(N__32133),
            .I(N__32130));
    LocalMux I__5132 (
            .O(N__32130),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_5 ));
    InMux I__5131 (
            .O(N__32127),
            .I(N__32124));
    LocalMux I__5130 (
            .O(N__32124),
            .I(N__32120));
    InMux I__5129 (
            .O(N__32123),
            .I(N__32117));
    Span4Mux_h I__5128 (
            .O(N__32120),
            .I(N__32114));
    LocalMux I__5127 (
            .O(N__32117),
            .I(N__32111));
    Span4Mux_h I__5126 (
            .O(N__32114),
            .I(N__32105));
    Span4Mux_h I__5125 (
            .O(N__32111),
            .I(N__32105));
    InMux I__5124 (
            .O(N__32110),
            .I(N__32102));
    Odrv4 I__5123 (
            .O(N__32105),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_5));
    LocalMux I__5122 (
            .O(N__32102),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_5));
    InMux I__5121 (
            .O(N__32097),
            .I(N__32094));
    LocalMux I__5120 (
            .O(N__32094),
            .I(N__32091));
    Span4Mux_v I__5119 (
            .O(N__32091),
            .I(N__32088));
    Span4Mux_h I__5118 (
            .O(N__32088),
            .I(N__32085));
    Sp12to4 I__5117 (
            .O(N__32085),
            .I(N__32082));
    Span12Mux_h I__5116 (
            .O(N__32082),
            .I(N__32077));
    InMux I__5115 (
            .O(N__32081),
            .I(N__32072));
    InMux I__5114 (
            .O(N__32080),
            .I(N__32072));
    Odrv12 I__5113 (
            .O(N__32077),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_14));
    LocalMux I__5112 (
            .O(N__32072),
            .I(cemf_module_64ch_ctrl_inst1_data_clkctrovf_14));
    CascadeMux I__5111 (
            .O(N__32067),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_242_cascade_ ));
    InMux I__5110 (
            .O(N__32064),
            .I(N__32061));
    LocalMux I__5109 (
            .O(N__32061),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_6 ));
    InMux I__5108 (
            .O(N__32058),
            .I(N__32052));
    InMux I__5107 (
            .O(N__32057),
            .I(N__32052));
    LocalMux I__5106 (
            .O(N__32052),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_7 ));
    InMux I__5105 (
            .O(N__32049),
            .I(N__32046));
    LocalMux I__5104 (
            .O(N__32046),
            .I(N__32043));
    Odrv4 I__5103 (
            .O(N__32043),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_6 ));
    CascadeMux I__5102 (
            .O(N__32040),
            .I(N__32036));
    InMux I__5101 (
            .O(N__32039),
            .I(N__32031));
    InMux I__5100 (
            .O(N__32036),
            .I(N__32031));
    LocalMux I__5099 (
            .O(N__32031),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_6));
    InMux I__5098 (
            .O(N__32028),
            .I(N__32025));
    LocalMux I__5097 (
            .O(N__32025),
            .I(N__32022));
    Span4Mux_h I__5096 (
            .O(N__32022),
            .I(N__32019));
    Span4Mux_v I__5095 (
            .O(N__32019),
            .I(N__32016));
    Odrv4 I__5094 (
            .O(N__32016),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_283 ));
    CascadeMux I__5093 (
            .O(N__32013),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_20_cascade_ ));
    CascadeMux I__5092 (
            .O(N__32010),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_20_cascade_ ));
    InMux I__5091 (
            .O(N__32007),
            .I(N__32004));
    LocalMux I__5090 (
            .O(N__32004),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_20 ));
    InMux I__5089 (
            .O(N__32001),
            .I(N__31998));
    LocalMux I__5088 (
            .O(N__31998),
            .I(N__31995));
    Span4Mux_v I__5087 (
            .O(N__31995),
            .I(N__31992));
    Odrv4 I__5086 (
            .O(N__31992),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_6 ));
    InMux I__5085 (
            .O(N__31989),
            .I(N__31986));
    LocalMux I__5084 (
            .O(N__31986),
            .I(N__31982));
    InMux I__5083 (
            .O(N__31985),
            .I(N__31978));
    Span4Mux_h I__5082 (
            .O(N__31982),
            .I(N__31975));
    InMux I__5081 (
            .O(N__31981),
            .I(N__31972));
    LocalMux I__5080 (
            .O(N__31978),
            .I(cemf_module_64ch_ctrl_inst1_data_config_6));
    Odrv4 I__5079 (
            .O(N__31975),
            .I(cemf_module_64ch_ctrl_inst1_data_config_6));
    LocalMux I__5078 (
            .O(N__31972),
            .I(cemf_module_64ch_ctrl_inst1_data_config_6));
    CascadeMux I__5077 (
            .O(N__31965),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_6_cascade_ ));
    CascadeMux I__5076 (
            .O(N__31962),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SLZ0Z7_cascade_ ));
    InMux I__5075 (
            .O(N__31959),
            .I(N__31956));
    LocalMux I__5074 (
            .O(N__31956),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRLZ0Z7 ));
    InMux I__5073 (
            .O(N__31953),
            .I(N__31950));
    LocalMux I__5072 (
            .O(N__31950),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6 ));
    InMux I__5071 (
            .O(N__31947),
            .I(N__31944));
    LocalMux I__5070 (
            .O(N__31944),
            .I(N__31941));
    Odrv4 I__5069 (
            .O(N__31941),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_5 ));
    CascadeMux I__5068 (
            .O(N__31938),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6_cascade_ ));
    InMux I__5067 (
            .O(N__31935),
            .I(N__31932));
    LocalMux I__5066 (
            .O(N__31932),
            .I(N__31929));
    Span4Mux_v I__5065 (
            .O(N__31929),
            .I(N__31926));
    Span4Mux_h I__5064 (
            .O(N__31926),
            .I(N__31923));
    Span4Mux_h I__5063 (
            .O(N__31923),
            .I(N__31920));
    Span4Mux_v I__5062 (
            .O(N__31920),
            .I(N__31917));
    Odrv4 I__5061 (
            .O(N__31917),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_11));
    CascadeMux I__5060 (
            .O(N__31914),
            .I(N__31911));
    InMux I__5059 (
            .O(N__31911),
            .I(N__31908));
    LocalMux I__5058 (
            .O(N__31908),
            .I(N__31905));
    Span4Mux_v I__5057 (
            .O(N__31905),
            .I(N__31902));
    Span4Mux_v I__5056 (
            .O(N__31902),
            .I(N__31899));
    Sp12to4 I__5055 (
            .O(N__31899),
            .I(N__31896));
    Odrv12 I__5054 (
            .O(N__31896),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_11));
    CascadeMux I__5053 (
            .O(N__31893),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_11_cascade_ ));
    InMux I__5052 (
            .O(N__31890),
            .I(N__31887));
    LocalMux I__5051 (
            .O(N__31887),
            .I(N__31884));
    Span4Mux_v I__5050 (
            .O(N__31884),
            .I(N__31881));
    Span4Mux_h I__5049 (
            .O(N__31881),
            .I(N__31878));
    Span4Mux_h I__5048 (
            .O(N__31878),
            .I(N__31875));
    Odrv4 I__5047 (
            .O(N__31875),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_11));
    InMux I__5046 (
            .O(N__31872),
            .I(N__31869));
    LocalMux I__5045 (
            .O(N__31869),
            .I(N__31866));
    Span4Mux_v I__5044 (
            .O(N__31866),
            .I(N__31863));
    Span4Mux_h I__5043 (
            .O(N__31863),
            .I(N__31860));
    Odrv4 I__5042 (
            .O(N__31860),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_819 ));
    CascadeMux I__5041 (
            .O(N__31857),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_11_cascade_ ));
    InMux I__5040 (
            .O(N__31854),
            .I(N__31851));
    LocalMux I__5039 (
            .O(N__31851),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_11 ));
    InMux I__5038 (
            .O(N__31848),
            .I(N__31845));
    LocalMux I__5037 (
            .O(N__31845),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_11 ));
    CascadeMux I__5036 (
            .O(N__31842),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_11_cascade_ ));
    InMux I__5035 (
            .O(N__31839),
            .I(N__31836));
    LocalMux I__5034 (
            .O(N__31836),
            .I(N__31833));
    Span4Mux_h I__5033 (
            .O(N__31833),
            .I(N__31830));
    Span4Mux_h I__5032 (
            .O(N__31830),
            .I(N__31827));
    Span4Mux_v I__5031 (
            .O(N__31827),
            .I(N__31824));
    Odrv4 I__5030 (
            .O(N__31824),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_19));
    InMux I__5029 (
            .O(N__31821),
            .I(N__31818));
    LocalMux I__5028 (
            .O(N__31818),
            .I(N__31815));
    Span4Mux_h I__5027 (
            .O(N__31815),
            .I(N__31812));
    Span4Mux_h I__5026 (
            .O(N__31812),
            .I(N__31809));
    Span4Mux_v I__5025 (
            .O(N__31809),
            .I(N__31806));
    Odrv4 I__5024 (
            .O(N__31806),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_20));
    CascadeMux I__5023 (
            .O(N__31803),
            .I(N__31800));
    InMux I__5022 (
            .O(N__31800),
            .I(N__31797));
    LocalMux I__5021 (
            .O(N__31797),
            .I(N__31794));
    Span4Mux_v I__5020 (
            .O(N__31794),
            .I(N__31791));
    Span4Mux_h I__5019 (
            .O(N__31791),
            .I(N__31788));
    Odrv4 I__5018 (
            .O(N__31788),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_20));
    CascadeMux I__5017 (
            .O(N__31785),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_20_cascade_ ));
    InMux I__5016 (
            .O(N__31782),
            .I(N__31779));
    LocalMux I__5015 (
            .O(N__31779),
            .I(N__31776));
    Span4Mux_h I__5014 (
            .O(N__31776),
            .I(N__31773));
    Span4Mux_h I__5013 (
            .O(N__31773),
            .I(N__31770));
    Span4Mux_h I__5012 (
            .O(N__31770),
            .I(N__31767));
    Odrv4 I__5011 (
            .O(N__31767),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_20));
    CascadeMux I__5010 (
            .O(N__31764),
            .I(N__31761));
    InMux I__5009 (
            .O(N__31761),
            .I(N__31758));
    LocalMux I__5008 (
            .O(N__31758),
            .I(N__31755));
    Span4Mux_h I__5007 (
            .O(N__31755),
            .I(N__31752));
    Span4Mux_h I__5006 (
            .O(N__31752),
            .I(N__31749));
    Odrv4 I__5005 (
            .O(N__31749),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_2));
    CascadeMux I__5004 (
            .O(N__31746),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_2_cascade_ ));
    CascadeMux I__5003 (
            .O(N__31743),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_2_cascade_ ));
    InMux I__5002 (
            .O(N__31740),
            .I(N__31737));
    LocalMux I__5001 (
            .O(N__31737),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_2 ));
    InMux I__5000 (
            .O(N__31734),
            .I(N__31731));
    LocalMux I__4999 (
            .O(N__31731),
            .I(N__31728));
    Span4Mux_h I__4998 (
            .O(N__31728),
            .I(N__31725));
    Span4Mux_v I__4997 (
            .O(N__31725),
            .I(N__31722));
    Span4Mux_v I__4996 (
            .O(N__31722),
            .I(N__31719));
    Odrv4 I__4995 (
            .O(N__31719),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_10));
    CascadeMux I__4994 (
            .O(N__31716),
            .I(N__31713));
    InMux I__4993 (
            .O(N__31713),
            .I(N__31710));
    LocalMux I__4992 (
            .O(N__31710),
            .I(N__31707));
    Span4Mux_v I__4991 (
            .O(N__31707),
            .I(N__31704));
    Span4Mux_h I__4990 (
            .O(N__31704),
            .I(N__31701));
    Odrv4 I__4989 (
            .O(N__31701),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_10));
    CascadeMux I__4988 (
            .O(N__31698),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_10_cascade_ ));
    InMux I__4987 (
            .O(N__31695),
            .I(N__31692));
    LocalMux I__4986 (
            .O(N__31692),
            .I(N__31689));
    Span4Mux_h I__4985 (
            .O(N__31689),
            .I(N__31686));
    Span4Mux_h I__4984 (
            .O(N__31686),
            .I(N__31683));
    Span4Mux_v I__4983 (
            .O(N__31683),
            .I(N__31680));
    Odrv4 I__4982 (
            .O(N__31680),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_10));
    InMux I__4981 (
            .O(N__31677),
            .I(N__31674));
    LocalMux I__4980 (
            .O(N__31674),
            .I(N__31671));
    Odrv12 I__4979 (
            .O(N__31671),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_830 ));
    CascadeMux I__4978 (
            .O(N__31668),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_10_cascade_ ));
    InMux I__4977 (
            .O(N__31665),
            .I(N__31662));
    LocalMux I__4976 (
            .O(N__31662),
            .I(N__31659));
    Span4Mux_h I__4975 (
            .O(N__31659),
            .I(N__31656));
    Odrv4 I__4974 (
            .O(N__31656),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_10 ));
    CascadeMux I__4973 (
            .O(N__31653),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_10_cascade_ ));
    InMux I__4972 (
            .O(N__31650),
            .I(N__31647));
    LocalMux I__4971 (
            .O(N__31647),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_10 ));
    InMux I__4970 (
            .O(N__31644),
            .I(N__31641));
    LocalMux I__4969 (
            .O(N__31641),
            .I(N__31638));
    Span4Mux_v I__4968 (
            .O(N__31638),
            .I(N__31635));
    Span4Mux_v I__4967 (
            .O(N__31635),
            .I(N__31632));
    Sp12to4 I__4966 (
            .O(N__31632),
            .I(N__31629));
    Odrv12 I__4965 (
            .O(N__31629),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_18));
    CascadeMux I__4964 (
            .O(N__31626),
            .I(N__31623));
    InMux I__4963 (
            .O(N__31623),
            .I(N__31620));
    LocalMux I__4962 (
            .O(N__31620),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_18 ));
    InMux I__4961 (
            .O(N__31617),
            .I(N__31614));
    LocalMux I__4960 (
            .O(N__31614),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_3 ));
    InMux I__4959 (
            .O(N__31611),
            .I(N__31608));
    LocalMux I__4958 (
            .O(N__31608),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_2 ));
    InMux I__4957 (
            .O(N__31605),
            .I(N__31602));
    LocalMux I__4956 (
            .O(N__31602),
            .I(N__31599));
    Odrv12 I__4955 (
            .O(N__31599),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_275_0 ));
    CascadeMux I__4954 (
            .O(N__31596),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_275_0_cascade_ ));
    CascadeMux I__4953 (
            .O(N__31593),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_2_cascade_ ));
    CascadeMux I__4952 (
            .O(N__31590),
            .I(N__31586));
    InMux I__4951 (
            .O(N__31589),
            .I(N__31583));
    InMux I__4950 (
            .O(N__31586),
            .I(N__31580));
    LocalMux I__4949 (
            .O(N__31583),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_59 ));
    LocalMux I__4948 (
            .O(N__31580),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.N_59 ));
    InMux I__4947 (
            .O(N__31575),
            .I(N__31572));
    LocalMux I__4946 (
            .O(N__31572),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_2 ));
    InMux I__4945 (
            .O(N__31569),
            .I(N__31566));
    LocalMux I__4944 (
            .O(N__31566),
            .I(N__31563));
    Span4Mux_v I__4943 (
            .O(N__31563),
            .I(N__31560));
    Span4Mux_h I__4942 (
            .O(N__31560),
            .I(N__31557));
    Span4Mux_h I__4941 (
            .O(N__31557),
            .I(N__31554));
    Odrv4 I__4940 (
            .O(N__31554),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_2));
    InMux I__4939 (
            .O(N__31551),
            .I(N__31548));
    LocalMux I__4938 (
            .O(N__31548),
            .I(N__31545));
    Span4Mux_h I__4937 (
            .O(N__31545),
            .I(N__31542));
    Odrv4 I__4936 (
            .O(N__31542),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1945 ));
    CascadeMux I__4935 (
            .O(N__31539),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2_cascade_ ));
    InMux I__4934 (
            .O(N__31536),
            .I(N__31533));
    LocalMux I__4933 (
            .O(N__31533),
            .I(N__31530));
    Span4Mux_h I__4932 (
            .O(N__31530),
            .I(N__31527));
    Odrv4 I__4931 (
            .O(N__31527),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1844 ));
    IoInMux I__4930 (
            .O(N__31524),
            .I(N__31521));
    LocalMux I__4929 (
            .O(N__31521),
            .I(N__31518));
    Span4Mux_s1_h I__4928 (
            .O(N__31518),
            .I(N__31515));
    Span4Mux_h I__4927 (
            .O(N__31515),
            .I(N__31512));
    Span4Mux_h I__4926 (
            .O(N__31512),
            .I(N__31509));
    Span4Mux_h I__4925 (
            .O(N__31509),
            .I(N__31506));
    Odrv4 I__4924 (
            .O(N__31506),
            .I(N_528_0));
    InMux I__4923 (
            .O(N__31503),
            .I(N__31500));
    LocalMux I__4922 (
            .O(N__31500),
            .I(N__31497));
    Odrv4 I__4921 (
            .O(N__31497),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_0 ));
    InMux I__4920 (
            .O(N__31494),
            .I(N__31491));
    LocalMux I__4919 (
            .O(N__31491),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_2 ));
    InMux I__4918 (
            .O(N__31488),
            .I(N__31482));
    InMux I__4917 (
            .O(N__31487),
            .I(N__31482));
    LocalMux I__4916 (
            .O(N__31482),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_1 ));
    InMux I__4915 (
            .O(N__31479),
            .I(N__31474));
    InMux I__4914 (
            .O(N__31478),
            .I(N__31471));
    InMux I__4913 (
            .O(N__31477),
            .I(N__31468));
    LocalMux I__4912 (
            .O(N__31474),
            .I(N__31465));
    LocalMux I__4911 (
            .O(N__31471),
            .I(\cemf_module_64ch_ctrl_inst1.n_state41 ));
    LocalMux I__4910 (
            .O(N__31468),
            .I(\cemf_module_64ch_ctrl_inst1.n_state41 ));
    Odrv4 I__4909 (
            .O(N__31465),
            .I(\cemf_module_64ch_ctrl_inst1.n_state41 ));
    CascadeMux I__4908 (
            .O(N__31458),
            .I(N__31452));
    CascadeMux I__4907 (
            .O(N__31457),
            .I(N__31448));
    InMux I__4906 (
            .O(N__31456),
            .I(N__31445));
    CascadeMux I__4905 (
            .O(N__31455),
            .I(N__31442));
    InMux I__4904 (
            .O(N__31452),
            .I(N__31439));
    InMux I__4903 (
            .O(N__31451),
            .I(N__31436));
    InMux I__4902 (
            .O(N__31448),
            .I(N__31433));
    LocalMux I__4901 (
            .O(N__31445),
            .I(N__31430));
    InMux I__4900 (
            .O(N__31442),
            .I(N__31427));
    LocalMux I__4899 (
            .O(N__31439),
            .I(N__31418));
    LocalMux I__4898 (
            .O(N__31436),
            .I(N__31418));
    LocalMux I__4897 (
            .O(N__31433),
            .I(N__31418));
    Span4Mux_h I__4896 (
            .O(N__31430),
            .I(N__31418));
    LocalMux I__4895 (
            .O(N__31427),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_19 ));
    Odrv4 I__4894 (
            .O(N__31418),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_19 ));
    InMux I__4893 (
            .O(N__31413),
            .I(N__31410));
    LocalMux I__4892 (
            .O(N__31410),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_1 ));
    InMux I__4891 (
            .O(N__31407),
            .I(N__31404));
    LocalMux I__4890 (
            .O(N__31404),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_0 ));
    InMux I__4889 (
            .O(N__31401),
            .I(N__31398));
    LocalMux I__4888 (
            .O(N__31398),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_1 ));
    CascadeMux I__4887 (
            .O(N__31395),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1_cascade_ ));
    InMux I__4886 (
            .O(N__31392),
            .I(N__31389));
    LocalMux I__4885 (
            .O(N__31389),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_1 ));
    InMux I__4884 (
            .O(N__31386),
            .I(N__31378));
    InMux I__4883 (
            .O(N__31385),
            .I(N__31378));
    InMux I__4882 (
            .O(N__31384),
            .I(N__31375));
    InMux I__4881 (
            .O(N__31383),
            .I(N__31372));
    LocalMux I__4880 (
            .O(N__31378),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3 ));
    LocalMux I__4879 (
            .O(N__31375),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3 ));
    LocalMux I__4878 (
            .O(N__31372),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3 ));
    CascadeMux I__4877 (
            .O(N__31365),
            .I(N__31361));
    InMux I__4876 (
            .O(N__31364),
            .I(N__31358));
    InMux I__4875 (
            .O(N__31361),
            .I(N__31355));
    LocalMux I__4874 (
            .O(N__31358),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2 ));
    LocalMux I__4873 (
            .O(N__31355),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2 ));
    InMux I__4872 (
            .O(N__31350),
            .I(N__31347));
    LocalMux I__4871 (
            .O(N__31347),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_4 ));
    InMux I__4870 (
            .O(N__31344),
            .I(N__31340));
    CascadeMux I__4869 (
            .O(N__31343),
            .I(N__31337));
    LocalMux I__4868 (
            .O(N__31340),
            .I(N__31333));
    InMux I__4867 (
            .O(N__31337),
            .I(N__31330));
    InMux I__4866 (
            .O(N__31336),
            .I(N__31327));
    Odrv12 I__4865 (
            .O(N__31333),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967 ));
    LocalMux I__4864 (
            .O(N__31330),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967 ));
    LocalMux I__4863 (
            .O(N__31327),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967 ));
    CascadeMux I__4862 (
            .O(N__31320),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_2_cascade_ ));
    CascadeMux I__4861 (
            .O(N__31317),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_3_cascade_ ));
    InMux I__4860 (
            .O(N__31314),
            .I(N__31311));
    LocalMux I__4859 (
            .O(N__31311),
            .I(N__31308));
    Span4Mux_v I__4858 (
            .O(N__31308),
            .I(N__31305));
    Odrv4 I__4857 (
            .O(N__31305),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2 ));
    CascadeMux I__4856 (
            .O(N__31302),
            .I(N__31298));
    InMux I__4855 (
            .O(N__31301),
            .I(N__31293));
    InMux I__4854 (
            .O(N__31298),
            .I(N__31293));
    LocalMux I__4853 (
            .O(N__31293),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_14 ));
    InMux I__4852 (
            .O(N__31290),
            .I(N__31287));
    LocalMux I__4851 (
            .O(N__31287),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_14 ));
    InMux I__4850 (
            .O(N__31284),
            .I(N__31275));
    InMux I__4849 (
            .O(N__31283),
            .I(N__31275));
    InMux I__4848 (
            .O(N__31282),
            .I(N__31268));
    InMux I__4847 (
            .O(N__31281),
            .I(N__31268));
    InMux I__4846 (
            .O(N__31280),
            .I(N__31268));
    LocalMux I__4845 (
            .O(N__31275),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12 ));
    LocalMux I__4844 (
            .O(N__31268),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12 ));
    InMux I__4843 (
            .O(N__31263),
            .I(N__31248));
    InMux I__4842 (
            .O(N__31262),
            .I(N__31248));
    InMux I__4841 (
            .O(N__31261),
            .I(N__31248));
    InMux I__4840 (
            .O(N__31260),
            .I(N__31241));
    InMux I__4839 (
            .O(N__31259),
            .I(N__31241));
    InMux I__4838 (
            .O(N__31258),
            .I(N__31241));
    InMux I__4837 (
            .O(N__31257),
            .I(N__31234));
    InMux I__4836 (
            .O(N__31256),
            .I(N__31234));
    InMux I__4835 (
            .O(N__31255),
            .I(N__31234));
    LocalMux I__4834 (
            .O(N__31248),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987 ));
    LocalMux I__4833 (
            .O(N__31241),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987 ));
    LocalMux I__4832 (
            .O(N__31234),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987 ));
    CascadeMux I__4831 (
            .O(N__31227),
            .I(N__31222));
    CascadeMux I__4830 (
            .O(N__31226),
            .I(N__31219));
    InMux I__4829 (
            .O(N__31225),
            .I(N__31215));
    InMux I__4828 (
            .O(N__31222),
            .I(N__31208));
    InMux I__4827 (
            .O(N__31219),
            .I(N__31208));
    InMux I__4826 (
            .O(N__31218),
            .I(N__31208));
    LocalMux I__4825 (
            .O(N__31215),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15 ));
    LocalMux I__4824 (
            .O(N__31208),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15 ));
    CascadeMux I__4823 (
            .O(N__31203),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967i_cascade_ ));
    InMux I__4822 (
            .O(N__31200),
            .I(N__31197));
    LocalMux I__4821 (
            .O(N__31197),
            .I(N__31194));
    Odrv4 I__4820 (
            .O(N__31194),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retZ0Z_13 ));
    InMux I__4819 (
            .O(N__31191),
            .I(N__31188));
    LocalMux I__4818 (
            .O(N__31188),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_276_reti ));
    CascadeMux I__4817 (
            .O(N__31185),
            .I(N__31181));
    InMux I__4816 (
            .O(N__31184),
            .I(N__31176));
    InMux I__4815 (
            .O(N__31181),
            .I(N__31176));
    LocalMux I__4814 (
            .O(N__31176),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_8_1 ));
    InMux I__4813 (
            .O(N__31173),
            .I(N__31168));
    InMux I__4812 (
            .O(N__31172),
            .I(N__31163));
    InMux I__4811 (
            .O(N__31171),
            .I(N__31163));
    LocalMux I__4810 (
            .O(N__31168),
            .I(N__31157));
    LocalMux I__4809 (
            .O(N__31163),
            .I(N__31154));
    InMux I__4808 (
            .O(N__31162),
            .I(N__31147));
    InMux I__4807 (
            .O(N__31161),
            .I(N__31147));
    InMux I__4806 (
            .O(N__31160),
            .I(N__31147));
    Odrv4 I__4805 (
            .O(N__31157),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8 ));
    Odrv4 I__4804 (
            .O(N__31154),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8 ));
    LocalMux I__4803 (
            .O(N__31147),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8 ));
    InMux I__4802 (
            .O(N__31140),
            .I(N__31134));
    InMux I__4801 (
            .O(N__31139),
            .I(N__31134));
    LocalMux I__4800 (
            .O(N__31134),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1 ));
    InMux I__4799 (
            .O(N__31131),
            .I(N__31128));
    LocalMux I__4798 (
            .O(N__31128),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_6 ));
    CascadeMux I__4797 (
            .O(N__31125),
            .I(N__31120));
    InMux I__4796 (
            .O(N__31124),
            .I(N__31116));
    InMux I__4795 (
            .O(N__31123),
            .I(N__31113));
    InMux I__4794 (
            .O(N__31120),
            .I(N__31108));
    InMux I__4793 (
            .O(N__31119),
            .I(N__31108));
    LocalMux I__4792 (
            .O(N__31116),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7 ));
    LocalMux I__4791 (
            .O(N__31113),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7 ));
    LocalMux I__4790 (
            .O(N__31108),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7 ));
    CascadeMux I__4789 (
            .O(N__31101),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.en_count_bits_0_i_a2_0_a2_1_cascade_ ));
    InMux I__4788 (
            .O(N__31098),
            .I(N__31095));
    LocalMux I__4787 (
            .O(N__31095),
            .I(N__31092));
    Span4Mux_v I__4786 (
            .O(N__31092),
            .I(N__31083));
    InMux I__4785 (
            .O(N__31091),
            .I(N__31078));
    InMux I__4784 (
            .O(N__31090),
            .I(N__31078));
    InMux I__4783 (
            .O(N__31089),
            .I(N__31071));
    InMux I__4782 (
            .O(N__31088),
            .I(N__31071));
    InMux I__4781 (
            .O(N__31087),
            .I(N__31071));
    InMux I__4780 (
            .O(N__31086),
            .I(N__31068));
    Span4Mux_h I__4779 (
            .O(N__31083),
            .I(N__31061));
    LocalMux I__4778 (
            .O(N__31078),
            .I(N__31061));
    LocalMux I__4777 (
            .O(N__31071),
            .I(N__31061));
    LocalMux I__4776 (
            .O(N__31068),
            .I(N__31056));
    Span4Mux_h I__4775 (
            .O(N__31061),
            .I(N__31056));
    Odrv4 I__4774 (
            .O(N__31056),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_277_0 ));
    InMux I__4773 (
            .O(N__31053),
            .I(N__31044));
    InMux I__4772 (
            .O(N__31052),
            .I(N__31044));
    InMux I__4771 (
            .O(N__31051),
            .I(N__31044));
    LocalMux I__4770 (
            .O(N__31044),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_19 ));
    InMux I__4769 (
            .O(N__31041),
            .I(N__31038));
    LocalMux I__4768 (
            .O(N__31038),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_18 ));
    InMux I__4767 (
            .O(N__31035),
            .I(N__31032));
    LocalMux I__4766 (
            .O(N__31032),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_13 ));
    InMux I__4765 (
            .O(N__31029),
            .I(N__31023));
    InMux I__4764 (
            .O(N__31028),
            .I(N__31020));
    InMux I__4763 (
            .O(N__31027),
            .I(N__31017));
    InMux I__4762 (
            .O(N__31026),
            .I(N__31014));
    LocalMux I__4761 (
            .O(N__31023),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11 ));
    LocalMux I__4760 (
            .O(N__31020),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11 ));
    LocalMux I__4759 (
            .O(N__31017),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11 ));
    LocalMux I__4758 (
            .O(N__31014),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11 ));
    SRMux I__4757 (
            .O(N__31005),
            .I(N__31002));
    LocalMux I__4756 (
            .O(N__31002),
            .I(N__30999));
    Span4Mux_v I__4755 (
            .O(N__30999),
            .I(N__30996));
    Span4Mux_h I__4754 (
            .O(N__30996),
            .I(N__30993));
    Odrv4 I__4753 (
            .O(N__30993),
            .I(\I2C_top_level_inst1.I2C_Control_StartUp_inst.N_8_i ));
    InMux I__4752 (
            .O(N__30990),
            .I(N__30986));
    InMux I__4751 (
            .O(N__30989),
            .I(N__30983));
    LocalMux I__4750 (
            .O(N__30986),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1 ));
    LocalMux I__4749 (
            .O(N__30983),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1 ));
    InMux I__4748 (
            .O(N__30978),
            .I(N__30975));
    LocalMux I__4747 (
            .O(N__30975),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0 ));
    CascadeMux I__4746 (
            .O(N__30972),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0_cascade_ ));
    InMux I__4745 (
            .O(N__30969),
            .I(N__30966));
    LocalMux I__4744 (
            .O(N__30966),
            .I(N__30963));
    Span4Mux_v I__4743 (
            .O(N__30963),
            .I(N__30959));
    InMux I__4742 (
            .O(N__30962),
            .I(N__30956));
    Span4Mux_h I__4741 (
            .O(N__30959),
            .I(N__30953));
    LocalMux I__4740 (
            .O(N__30956),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26 ));
    Odrv4 I__4739 (
            .O(N__30953),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26 ));
    CascadeMux I__4738 (
            .O(N__30948),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3Z0Z_0_cascade_ ));
    CascadeMux I__4737 (
            .O(N__30945),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1959_cascade_ ));
    CascadeMux I__4736 (
            .O(N__30942),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0_cascade_ ));
    CascadeMux I__4735 (
            .O(N__30939),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRLZ0Z7_cascade_ ));
    InMux I__4734 (
            .O(N__30936),
            .I(N__30933));
    LocalMux I__4733 (
            .O(N__30933),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3 ));
    CascadeMux I__4732 (
            .O(N__30930),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3_cascade_ ));
    InMux I__4731 (
            .O(N__30927),
            .I(N__30924));
    LocalMux I__4730 (
            .O(N__30924),
            .I(N__30921));
    Odrv4 I__4729 (
            .O(N__30921),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5 ));
    CascadeMux I__4728 (
            .O(N__30918),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5_cascade_ ));
    InMux I__4727 (
            .O(N__30915),
            .I(N__30912));
    LocalMux I__4726 (
            .O(N__30912),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_3 ));
    InMux I__4725 (
            .O(N__30909),
            .I(N__30906));
    LocalMux I__4724 (
            .O(N__30906),
            .I(N__30902));
    InMux I__4723 (
            .O(N__30905),
            .I(N__30899));
    Span4Mux_h I__4722 (
            .O(N__30902),
            .I(N__30896));
    LocalMux I__4721 (
            .O(N__30899),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4 ));
    Odrv4 I__4720 (
            .O(N__30896),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4 ));
    InMux I__4719 (
            .O(N__30891),
            .I(N__30888));
    LocalMux I__4718 (
            .O(N__30888),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_4 ));
    InMux I__4717 (
            .O(N__30885),
            .I(N__30882));
    LocalMux I__4716 (
            .O(N__30882),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_9 ));
    CascadeMux I__4715 (
            .O(N__30879),
            .I(N__30875));
    InMux I__4714 (
            .O(N__30878),
            .I(N__30870));
    InMux I__4713 (
            .O(N__30875),
            .I(N__30870));
    LocalMux I__4712 (
            .O(N__30870),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_9));
    InMux I__4711 (
            .O(N__30867),
            .I(N__30863));
    InMux I__4710 (
            .O(N__30866),
            .I(N__30860));
    LocalMux I__4709 (
            .O(N__30863),
            .I(N__30857));
    LocalMux I__4708 (
            .O(N__30860),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_22));
    Odrv12 I__4707 (
            .O(N__30857),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_22));
    CascadeMux I__4706 (
            .O(N__30852),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_13_cascade_ ));
    CascadeMux I__4705 (
            .O(N__30849),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GHZ0Z5_cascade_ ));
    InMux I__4704 (
            .O(N__30846),
            .I(N__30843));
    LocalMux I__4703 (
            .O(N__30843),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13 ));
    CascadeMux I__4702 (
            .O(N__30840),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13_cascade_ ));
    InMux I__4701 (
            .O(N__30837),
            .I(N__30834));
    LocalMux I__4700 (
            .O(N__30834),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3QZ0Z5 ));
    InMux I__4699 (
            .O(N__30831),
            .I(N__30828));
    LocalMux I__4698 (
            .O(N__30828),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4 ));
    CascadeMux I__4697 (
            .O(N__30825),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4_cascade_ ));
    InMux I__4696 (
            .O(N__30822),
            .I(N__30819));
    LocalMux I__4695 (
            .O(N__30819),
            .I(N__30816));
    Odrv4 I__4694 (
            .O(N__30816),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_4 ));
    InMux I__4693 (
            .O(N__30813),
            .I(N__30810));
    LocalMux I__4692 (
            .O(N__30810),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_13 ));
    CascadeMux I__4691 (
            .O(N__30807),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_3_cascade_ ));
    InMux I__4690 (
            .O(N__30804),
            .I(N__30801));
    LocalMux I__4689 (
            .O(N__30801),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_17 ));
    CascadeMux I__4688 (
            .O(N__30798),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_18_cascade_ ));
    CascadeMux I__4687 (
            .O(N__30795),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_18_cascade_ ));
    InMux I__4686 (
            .O(N__30792),
            .I(N__30789));
    LocalMux I__4685 (
            .O(N__30789),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_18 ));
    InMux I__4684 (
            .O(N__30786),
            .I(N__30783));
    LocalMux I__4683 (
            .O(N__30783),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_18 ));
    InMux I__4682 (
            .O(N__30780),
            .I(N__30777));
    LocalMux I__4681 (
            .O(N__30777),
            .I(N__30774));
    Odrv4 I__4680 (
            .O(N__30774),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_13 ));
    InMux I__4679 (
            .O(N__30771),
            .I(N__30768));
    LocalMux I__4678 (
            .O(N__30768),
            .I(N__30765));
    Span4Mux_v I__4677 (
            .O(N__30765),
            .I(N__30762));
    Odrv4 I__4676 (
            .O(N__30762),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_14 ));
    InMux I__4675 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__4674 (
            .O(N__30756),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_15 ));
    SRMux I__4673 (
            .O(N__30753),
            .I(N__30750));
    LocalMux I__4672 (
            .O(N__30750),
            .I(N__30747));
    Odrv4 I__4671 (
            .O(N__30747),
            .I(\I2C_top_level_inst1.I2C_Control_StartUp_inst.rst_neg_i ));
    InMux I__4670 (
            .O(N__30744),
            .I(N__30741));
    LocalMux I__4669 (
            .O(N__30741),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_22 ));
    InMux I__4668 (
            .O(N__30738),
            .I(N__30735));
    LocalMux I__4667 (
            .O(N__30735),
            .I(N__30732));
    Span4Mux_h I__4666 (
            .O(N__30732),
            .I(N__30729));
    Span4Mux_v I__4665 (
            .O(N__30729),
            .I(N__30726));
    Span4Mux_h I__4664 (
            .O(N__30726),
            .I(N__30723));
    Odrv4 I__4663 (
            .O(N__30723),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_2));
    InMux I__4662 (
            .O(N__30720),
            .I(N__30717));
    LocalMux I__4661 (
            .O(N__30717),
            .I(N__30714));
    Span12Mux_v I__4660 (
            .O(N__30714),
            .I(N__30711));
    Odrv12 I__4659 (
            .O(N__30711),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_13));
    CascadeMux I__4658 (
            .O(N__30708),
            .I(N__30705));
    InMux I__4657 (
            .O(N__30705),
            .I(N__30702));
    LocalMux I__4656 (
            .O(N__30702),
            .I(N__30699));
    Span4Mux_h I__4655 (
            .O(N__30699),
            .I(N__30696));
    Span4Mux_v I__4654 (
            .O(N__30696),
            .I(N__30693));
    Odrv4 I__4653 (
            .O(N__30693),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_13));
    CascadeMux I__4652 (
            .O(N__30690),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_13_cascade_ ));
    InMux I__4651 (
            .O(N__30687),
            .I(N__30684));
    LocalMux I__4650 (
            .O(N__30684),
            .I(N__30681));
    Span4Mux_h I__4649 (
            .O(N__30681),
            .I(N__30678));
    Span4Mux_h I__4648 (
            .O(N__30678),
            .I(N__30675));
    Odrv4 I__4647 (
            .O(N__30675),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_13));
    InMux I__4646 (
            .O(N__30672),
            .I(N__30669));
    LocalMux I__4645 (
            .O(N__30669),
            .I(N__30666));
    Span4Mux_v I__4644 (
            .O(N__30666),
            .I(N__30663));
    Span4Mux_v I__4643 (
            .O(N__30663),
            .I(N__30660));
    Odrv4 I__4642 (
            .O(N__30660),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_797 ));
    CascadeMux I__4641 (
            .O(N__30657),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_13_cascade_ ));
    InMux I__4640 (
            .O(N__30654),
            .I(N__30651));
    LocalMux I__4639 (
            .O(N__30651),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_13 ));
    CascadeMux I__4638 (
            .O(N__30648),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_13_cascade_ ));
    InMux I__4637 (
            .O(N__30645),
            .I(N__30642));
    LocalMux I__4636 (
            .O(N__30642),
            .I(N__30639));
    Span4Mux_h I__4635 (
            .O(N__30639),
            .I(N__30636));
    Span4Mux_h I__4634 (
            .O(N__30636),
            .I(N__30633));
    Odrv4 I__4633 (
            .O(N__30633),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_18));
    CascadeMux I__4632 (
            .O(N__30630),
            .I(N__30627));
    InMux I__4631 (
            .O(N__30627),
            .I(N__30624));
    LocalMux I__4630 (
            .O(N__30624),
            .I(N__30621));
    Span4Mux_h I__4629 (
            .O(N__30621),
            .I(N__30618));
    Span4Mux_h I__4628 (
            .O(N__30618),
            .I(N__30615));
    Span4Mux_h I__4627 (
            .O(N__30615),
            .I(N__30612));
    Odrv4 I__4626 (
            .O(N__30612),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_18));
    InMux I__4625 (
            .O(N__30609),
            .I(N__30603));
    InMux I__4624 (
            .O(N__30608),
            .I(N__30603));
    LocalMux I__4623 (
            .O(N__30603),
            .I(N__30600));
    Odrv4 I__4622 (
            .O(N__30600),
            .I(\cemf_module_64ch_ctrl_inst1.N_410_0 ));
    CascadeMux I__4621 (
            .O(N__30597),
            .I(N__30592));
    InMux I__4620 (
            .O(N__30596),
            .I(N__30589));
    InMux I__4619 (
            .O(N__30595),
            .I(N__30584));
    InMux I__4618 (
            .O(N__30592),
            .I(N__30584));
    LocalMux I__4617 (
            .O(N__30589),
            .I(N__30581));
    LocalMux I__4616 (
            .O(N__30584),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_7 ));
    Odrv4 I__4615 (
            .O(N__30581),
            .I(\cemf_module_64ch_ctrl_inst1.c_state_7 ));
    InMux I__4614 (
            .O(N__30576),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0 ));
    InMux I__4613 (
            .O(N__30573),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1 ));
    InMux I__4612 (
            .O(N__30570),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_2 ));
    InMux I__4611 (
            .O(N__30567),
            .I(N__30564));
    LocalMux I__4610 (
            .O(N__30564),
            .I(\I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetterZ0 ));
    CascadeMux I__4609 (
            .O(N__30561),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1_cascade_ ));
    InMux I__4608 (
            .O(N__30558),
            .I(N__30549));
    InMux I__4607 (
            .O(N__30557),
            .I(N__30549));
    InMux I__4606 (
            .O(N__30556),
            .I(N__30542));
    InMux I__4605 (
            .O(N__30555),
            .I(N__30542));
    InMux I__4604 (
            .O(N__30554),
            .I(N__30542));
    LocalMux I__4603 (
            .O(N__30549),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4 ));
    LocalMux I__4602 (
            .O(N__30542),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4 ));
    InMux I__4601 (
            .O(N__30537),
            .I(N__30534));
    LocalMux I__4600 (
            .O(N__30534),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1 ));
    CascadeMux I__4599 (
            .O(N__30531),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_2_cascade_ ));
    CascadeMux I__4598 (
            .O(N__30528),
            .I(N__30525));
    InMux I__4597 (
            .O(N__30525),
            .I(N__30522));
    LocalMux I__4596 (
            .O(N__30522),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_9 ));
    InMux I__4595 (
            .O(N__30519),
            .I(N__30516));
    LocalMux I__4594 (
            .O(N__30516),
            .I(N__30510));
    InMux I__4593 (
            .O(N__30515),
            .I(N__30507));
    InMux I__4592 (
            .O(N__30514),
            .I(N__30504));
    InMux I__4591 (
            .O(N__30513),
            .I(N__30501));
    Span4Mux_v I__4590 (
            .O(N__30510),
            .I(N__30498));
    LocalMux I__4589 (
            .O(N__30507),
            .I(N__30495));
    LocalMux I__4588 (
            .O(N__30504),
            .I(N__30492));
    LocalMux I__4587 (
            .O(N__30501),
            .I(N__30489));
    Span4Mux_h I__4586 (
            .O(N__30498),
            .I(N__30484));
    Span4Mux_v I__4585 (
            .O(N__30495),
            .I(N__30484));
    Odrv4 I__4584 (
            .O(N__30492),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9 ));
    Odrv4 I__4583 (
            .O(N__30489),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9 ));
    Odrv4 I__4582 (
            .O(N__30484),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9 ));
    InMux I__4581 (
            .O(N__30477),
            .I(N__30464));
    InMux I__4580 (
            .O(N__30476),
            .I(N__30464));
    InMux I__4579 (
            .O(N__30475),
            .I(N__30464));
    CascadeMux I__4578 (
            .O(N__30474),
            .I(N__30455));
    InMux I__4577 (
            .O(N__30473),
            .I(N__30452));
    InMux I__4576 (
            .O(N__30472),
            .I(N__30449));
    CascadeMux I__4575 (
            .O(N__30471),
            .I(N__30446));
    LocalMux I__4574 (
            .O(N__30464),
            .I(N__30443));
    InMux I__4573 (
            .O(N__30463),
            .I(N__30430));
    InMux I__4572 (
            .O(N__30462),
            .I(N__30430));
    InMux I__4571 (
            .O(N__30461),
            .I(N__30430));
    InMux I__4570 (
            .O(N__30460),
            .I(N__30430));
    InMux I__4569 (
            .O(N__30459),
            .I(N__30430));
    InMux I__4568 (
            .O(N__30458),
            .I(N__30430));
    InMux I__4567 (
            .O(N__30455),
            .I(N__30427));
    LocalMux I__4566 (
            .O(N__30452),
            .I(N__30424));
    LocalMux I__4565 (
            .O(N__30449),
            .I(N__30421));
    InMux I__4564 (
            .O(N__30446),
            .I(N__30418));
    Span4Mux_v I__4563 (
            .O(N__30443),
            .I(N__30413));
    LocalMux I__4562 (
            .O(N__30430),
            .I(N__30413));
    LocalMux I__4561 (
            .O(N__30427),
            .I(N__30410));
    Span4Mux_v I__4560 (
            .O(N__30424),
            .I(N__30405));
    Span4Mux_v I__4559 (
            .O(N__30421),
            .I(N__30405));
    LocalMux I__4558 (
            .O(N__30418),
            .I(N__30402));
    Span4Mux_h I__4557 (
            .O(N__30413),
            .I(N__30397));
    Span4Mux_v I__4556 (
            .O(N__30410),
            .I(N__30397));
    Span4Mux_h I__4555 (
            .O(N__30405),
            .I(N__30394));
    Span4Mux_h I__4554 (
            .O(N__30402),
            .I(N__30391));
    Span4Mux_h I__4553 (
            .O(N__30397),
            .I(N__30388));
    Odrv4 I__4552 (
            .O(N__30394),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10 ));
    Odrv4 I__4551 (
            .O(N__30391),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10 ));
    Odrv4 I__4550 (
            .O(N__30388),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10 ));
    InMux I__4549 (
            .O(N__30381),
            .I(N__30374));
    InMux I__4548 (
            .O(N__30380),
            .I(N__30374));
    InMux I__4547 (
            .O(N__30379),
            .I(N__30371));
    LocalMux I__4546 (
            .O(N__30374),
            .I(N__30368));
    LocalMux I__4545 (
            .O(N__30371),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9 ));
    Odrv4 I__4544 (
            .O(N__30368),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9 ));
    InMux I__4543 (
            .O(N__30363),
            .I(N__30360));
    LocalMux I__4542 (
            .O(N__30360),
            .I(N__30357));
    Odrv4 I__4541 (
            .O(N__30357),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_10 ));
    InMux I__4540 (
            .O(N__30354),
            .I(N__30351));
    LocalMux I__4539 (
            .O(N__30351),
            .I(N__30346));
    InMux I__4538 (
            .O(N__30350),
            .I(N__30341));
    InMux I__4537 (
            .O(N__30349),
            .I(N__30341));
    Odrv12 I__4536 (
            .O(N__30346),
            .I(\cemf_module_64ch_ctrl_inst1.N_68_0 ));
    LocalMux I__4535 (
            .O(N__30341),
            .I(\cemf_module_64ch_ctrl_inst1.N_68_0 ));
    InMux I__4534 (
            .O(N__30336),
            .I(N__30332));
    InMux I__4533 (
            .O(N__30335),
            .I(N__30329));
    LocalMux I__4532 (
            .O(N__30332),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4 ));
    LocalMux I__4531 (
            .O(N__30329),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4 ));
    InMux I__4530 (
            .O(N__30324),
            .I(N__30320));
    InMux I__4529 (
            .O(N__30323),
            .I(N__30317));
    LocalMux I__4528 (
            .O(N__30320),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3 ));
    LocalMux I__4527 (
            .O(N__30317),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3 ));
    InMux I__4526 (
            .O(N__30312),
            .I(N__30308));
    InMux I__4525 (
            .O(N__30311),
            .I(N__30305));
    LocalMux I__4524 (
            .O(N__30308),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2 ));
    LocalMux I__4523 (
            .O(N__30305),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2 ));
    InMux I__4522 (
            .O(N__30300),
            .I(N__30296));
    InMux I__4521 (
            .O(N__30299),
            .I(N__30293));
    LocalMux I__4520 (
            .O(N__30296),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1 ));
    LocalMux I__4519 (
            .O(N__30293),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1 ));
    CascadeMux I__4518 (
            .O(N__30288),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ns_i_a2_1_1_3_cascade_ ));
    InMux I__4517 (
            .O(N__30285),
            .I(N__30281));
    InMux I__4516 (
            .O(N__30284),
            .I(N__30278));
    LocalMux I__4515 (
            .O(N__30281),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0 ));
    LocalMux I__4514 (
            .O(N__30278),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0 ));
    CascadeMux I__4513 (
            .O(N__30273),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987_cascade_ ));
    InMux I__4512 (
            .O(N__30270),
            .I(N__30267));
    LocalMux I__4511 (
            .O(N__30267),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_2 ));
    CascadeMux I__4510 (
            .O(N__30264),
            .I(N__30261));
    InMux I__4509 (
            .O(N__30261),
            .I(N__30256));
    InMux I__4508 (
            .O(N__30260),
            .I(N__30251));
    InMux I__4507 (
            .O(N__30259),
            .I(N__30251));
    LocalMux I__4506 (
            .O(N__30256),
            .I(N__30246));
    LocalMux I__4505 (
            .O(N__30251),
            .I(N__30246));
    Odrv4 I__4504 (
            .O(N__30246),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_0 ));
    InMux I__4503 (
            .O(N__30243),
            .I(N__30239));
    InMux I__4502 (
            .O(N__30242),
            .I(N__30235));
    LocalMux I__4501 (
            .O(N__30239),
            .I(N__30232));
    InMux I__4500 (
            .O(N__30238),
            .I(N__30229));
    LocalMux I__4499 (
            .O(N__30235),
            .I(N__30226));
    Odrv12 I__4498 (
            .O(N__30232),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291 ));
    LocalMux I__4497 (
            .O(N__30229),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291 ));
    Odrv4 I__4496 (
            .O(N__30226),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291 ));
    InMux I__4495 (
            .O(N__30219),
            .I(N__30216));
    LocalMux I__4494 (
            .O(N__30216),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_5 ));
    CascadeMux I__4493 (
            .O(N__30213),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_o3_i_a2_1_1_cascade_ ));
    InMux I__4492 (
            .O(N__30210),
            .I(N__30207));
    LocalMux I__4491 (
            .O(N__30207),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_6 ));
    InMux I__4490 (
            .O(N__30204),
            .I(N__30195));
    InMux I__4489 (
            .O(N__30203),
            .I(N__30195));
    InMux I__4488 (
            .O(N__30202),
            .I(N__30195));
    LocalMux I__4487 (
            .O(N__30195),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_5 ));
    InMux I__4486 (
            .O(N__30192),
            .I(N__30189));
    LocalMux I__4485 (
            .O(N__30189),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_10 ));
    InMux I__4484 (
            .O(N__30186),
            .I(N__30183));
    LocalMux I__4483 (
            .O(N__30183),
            .I(N__30180));
    Span12Mux_v I__4482 (
            .O(N__30180),
            .I(N__30177));
    Odrv12 I__4481 (
            .O(N__30177),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_4));
    InMux I__4480 (
            .O(N__30174),
            .I(N__30171));
    LocalMux I__4479 (
            .O(N__30171),
            .I(N__30168));
    Span4Mux_h I__4478 (
            .O(N__30168),
            .I(N__30165));
    Odrv4 I__4477 (
            .O(N__30165),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_896 ));
    CascadeMux I__4476 (
            .O(N__30162),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_291_reti_cascade_ ));
    InMux I__4475 (
            .O(N__30159),
            .I(N__30156));
    LocalMux I__4474 (
            .O(N__30156),
            .I(N__30153));
    Odrv4 I__4473 (
            .O(N__30153),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_276i ));
    InMux I__4472 (
            .O(N__30150),
            .I(N__30147));
    LocalMux I__4471 (
            .O(N__30147),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_retZ0Z_4 ));
    CascadeMux I__4470 (
            .O(N__30144),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_4_0_cascade_ ));
    InMux I__4469 (
            .O(N__30141),
            .I(N__30138));
    LocalMux I__4468 (
            .O(N__30138),
            .I(N__30134));
    InMux I__4467 (
            .O(N__30137),
            .I(N__30131));
    Span4Mux_h I__4466 (
            .O(N__30134),
            .I(N__30128));
    LocalMux I__4465 (
            .O(N__30131),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283 ));
    Odrv4 I__4464 (
            .O(N__30128),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283 ));
    InMux I__4463 (
            .O(N__30123),
            .I(N__30118));
    CascadeMux I__4462 (
            .O(N__30122),
            .I(N__30115));
    InMux I__4461 (
            .O(N__30121),
            .I(N__30112));
    LocalMux I__4460 (
            .O(N__30118),
            .I(N__30109));
    InMux I__4459 (
            .O(N__30115),
            .I(N__30106));
    LocalMux I__4458 (
            .O(N__30112),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10 ));
    Odrv4 I__4457 (
            .O(N__30109),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10 ));
    LocalMux I__4456 (
            .O(N__30106),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10 ));
    CascadeMux I__4455 (
            .O(N__30099),
            .I(N__30096));
    InMux I__4454 (
            .O(N__30096),
            .I(N__30093));
    LocalMux I__4453 (
            .O(N__30093),
            .I(N__30090));
    Span4Mux_h I__4452 (
            .O(N__30090),
            .I(N__30087));
    Odrv4 I__4451 (
            .O(N__30087),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287 ));
    CascadeMux I__4450 (
            .O(N__30084),
            .I(N__30078));
    InMux I__4449 (
            .O(N__30083),
            .I(N__30074));
    InMux I__4448 (
            .O(N__30082),
            .I(N__30071));
    InMux I__4447 (
            .O(N__30081),
            .I(N__30068));
    InMux I__4446 (
            .O(N__30078),
            .I(N__30063));
    InMux I__4445 (
            .O(N__30077),
            .I(N__30063));
    LocalMux I__4444 (
            .O(N__30074),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11 ));
    LocalMux I__4443 (
            .O(N__30071),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11 ));
    LocalMux I__4442 (
            .O(N__30068),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11 ));
    LocalMux I__4441 (
            .O(N__30063),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11 ));
    CascadeMux I__4440 (
            .O(N__30054),
            .I(N__30049));
    InMux I__4439 (
            .O(N__30053),
            .I(N__30046));
    InMux I__4438 (
            .O(N__30052),
            .I(N__30041));
    InMux I__4437 (
            .O(N__30049),
            .I(N__30041));
    LocalMux I__4436 (
            .O(N__30046),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14 ));
    LocalMux I__4435 (
            .O(N__30041),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14 ));
    InMux I__4434 (
            .O(N__30036),
            .I(N__30030));
    CascadeMux I__4433 (
            .O(N__30035),
            .I(N__30027));
    InMux I__4432 (
            .O(N__30034),
            .I(N__30023));
    InMux I__4431 (
            .O(N__30033),
            .I(N__30020));
    LocalMux I__4430 (
            .O(N__30030),
            .I(N__30017));
    InMux I__4429 (
            .O(N__30027),
            .I(N__30012));
    InMux I__4428 (
            .O(N__30026),
            .I(N__30012));
    LocalMux I__4427 (
            .O(N__30023),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15 ));
    LocalMux I__4426 (
            .O(N__30020),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15 ));
    Odrv4 I__4425 (
            .O(N__30017),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15 ));
    LocalMux I__4424 (
            .O(N__30012),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15 ));
    CascadeMux I__4423 (
            .O(N__30003),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_2_0_cascade_ ));
    InMux I__4422 (
            .O(N__30000),
            .I(N__29996));
    InMux I__4421 (
            .O(N__29999),
            .I(N__29993));
    LocalMux I__4420 (
            .O(N__29996),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286 ));
    LocalMux I__4419 (
            .O(N__29993),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286 ));
    CascadeMux I__4418 (
            .O(N__29988),
            .I(N__29983));
    InMux I__4417 (
            .O(N__29987),
            .I(N__29976));
    InMux I__4416 (
            .O(N__29986),
            .I(N__29976));
    InMux I__4415 (
            .O(N__29983),
            .I(N__29976));
    LocalMux I__4414 (
            .O(N__29976),
            .I(N__29973));
    Odrv4 I__4413 (
            .O(N__29973),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_0_0 ));
    CascadeMux I__4412 (
            .O(N__29970),
            .I(N__29965));
    CascadeMux I__4411 (
            .O(N__29969),
            .I(N__29962));
    CascadeMux I__4410 (
            .O(N__29968),
            .I(N__29959));
    InMux I__4409 (
            .O(N__29965),
            .I(N__29952));
    InMux I__4408 (
            .O(N__29962),
            .I(N__29952));
    InMux I__4407 (
            .O(N__29959),
            .I(N__29943));
    InMux I__4406 (
            .O(N__29958),
            .I(N__29943));
    InMux I__4405 (
            .O(N__29957),
            .I(N__29943));
    LocalMux I__4404 (
            .O(N__29952),
            .I(N__29937));
    InMux I__4403 (
            .O(N__29951),
            .I(N__29932));
    InMux I__4402 (
            .O(N__29950),
            .I(N__29932));
    LocalMux I__4401 (
            .O(N__29943),
            .I(N__29929));
    InMux I__4400 (
            .O(N__29942),
            .I(N__29924));
    InMux I__4399 (
            .O(N__29941),
            .I(N__29924));
    CascadeMux I__4398 (
            .O(N__29940),
            .I(N__29921));
    Span4Mux_v I__4397 (
            .O(N__29937),
            .I(N__29913));
    LocalMux I__4396 (
            .O(N__29932),
            .I(N__29913));
    Span4Mux_v I__4395 (
            .O(N__29929),
            .I(N__29913));
    LocalMux I__4394 (
            .O(N__29924),
            .I(N__29910));
    InMux I__4393 (
            .O(N__29921),
            .I(N__29905));
    InMux I__4392 (
            .O(N__29920),
            .I(N__29905));
    Span4Mux_h I__4391 (
            .O(N__29913),
            .I(N__29900));
    Span4Mux_v I__4390 (
            .O(N__29910),
            .I(N__29900));
    LocalMux I__4389 (
            .O(N__29905),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0 ));
    Odrv4 I__4388 (
            .O(N__29900),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0 ));
    CascadeMux I__4387 (
            .O(N__29895),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_6_cascade_ ));
    CascadeMux I__4386 (
            .O(N__29892),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3QZ0Z5_cascade_ ));
    InMux I__4385 (
            .O(N__29889),
            .I(N__29885));
    InMux I__4384 (
            .O(N__29888),
            .I(N__29882));
    LocalMux I__4383 (
            .O(N__29885),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6 ));
    LocalMux I__4382 (
            .O(N__29882),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6 ));
    InMux I__4381 (
            .O(N__29877),
            .I(N__29874));
    LocalMux I__4380 (
            .O(N__29874),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3QZ0Z5 ));
    InMux I__4379 (
            .O(N__29871),
            .I(N__29868));
    LocalMux I__4378 (
            .O(N__29868),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5 ));
    CascadeMux I__4377 (
            .O(N__29865),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5_cascade_ ));
    InMux I__4376 (
            .O(N__29862),
            .I(N__29859));
    LocalMux I__4375 (
            .O(N__29859),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_5 ));
    InMux I__4374 (
            .O(N__29856),
            .I(N__29852));
    InMux I__4373 (
            .O(N__29855),
            .I(N__29849));
    LocalMux I__4372 (
            .O(N__29852),
            .I(N__29846));
    LocalMux I__4371 (
            .O(N__29849),
            .I(\cemf_module_64ch_ctrl_inst1.N_1615 ));
    Odrv12 I__4370 (
            .O(N__29846),
            .I(\cemf_module_64ch_ctrl_inst1.N_1615 ));
    CascadeMux I__4369 (
            .O(N__29841),
            .I(N_1614_cascade_));
    InMux I__4368 (
            .O(N__29838),
            .I(N__29835));
    LocalMux I__4367 (
            .O(N__29835),
            .I(N__29832));
    Span4Mux_v I__4366 (
            .O(N__29832),
            .I(N__29829));
    Span4Mux_h I__4365 (
            .O(N__29829),
            .I(N__29826));
    Odrv4 I__4364 (
            .O(N__29826),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_28));
    InMux I__4363 (
            .O(N__29823),
            .I(N__29820));
    LocalMux I__4362 (
            .O(N__29820),
            .I(N__29817));
    Odrv12 I__4361 (
            .O(N__29817),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_643 ));
    InMux I__4360 (
            .O(N__29814),
            .I(N__29811));
    LocalMux I__4359 (
            .O(N__29811),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_5 ));
    InMux I__4358 (
            .O(N__29808),
            .I(N__29805));
    LocalMux I__4357 (
            .O(N__29805),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_6 ));
    InMux I__4356 (
            .O(N__29802),
            .I(N__29799));
    LocalMux I__4355 (
            .O(N__29799),
            .I(N__29796));
    Span4Mux_v I__4354 (
            .O(N__29796),
            .I(N__29793));
    Span4Mux_h I__4353 (
            .O(N__29793),
            .I(N__29790));
    Span4Mux_v I__4352 (
            .O(N__29790),
            .I(N__29787));
    Span4Mux_v I__4351 (
            .O(N__29787),
            .I(N__29784));
    Odrv4 I__4350 (
            .O(N__29784),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_6));
    CascadeMux I__4349 (
            .O(N__29781),
            .I(N__29778));
    InMux I__4348 (
            .O(N__29778),
            .I(N__29775));
    LocalMux I__4347 (
            .O(N__29775),
            .I(N__29772));
    Span4Mux_v I__4346 (
            .O(N__29772),
            .I(N__29769));
    Span4Mux_v I__4345 (
            .O(N__29769),
            .I(N__29766));
    Span4Mux_h I__4344 (
            .O(N__29766),
            .I(N__29763));
    Odrv4 I__4343 (
            .O(N__29763),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_6));
    InMux I__4342 (
            .O(N__29760),
            .I(N__29757));
    LocalMux I__4341 (
            .O(N__29757),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_6 ));
    InMux I__4340 (
            .O(N__29754),
            .I(N__29751));
    LocalMux I__4339 (
            .O(N__29751),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_9 ));
    CascadeMux I__4338 (
            .O(N__29748),
            .I(N__29745));
    InMux I__4337 (
            .O(N__29745),
            .I(N__29742));
    LocalMux I__4336 (
            .O(N__29742),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_841 ));
    CascadeMux I__4335 (
            .O(N__29739),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_9_cascade_ ));
    InMux I__4334 (
            .O(N__29736),
            .I(N__29733));
    LocalMux I__4333 (
            .O(N__29733),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_9 ));
    InMux I__4332 (
            .O(N__29730),
            .I(N__29727));
    LocalMux I__4331 (
            .O(N__29727),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_9 ));
    InMux I__4330 (
            .O(N__29724),
            .I(N__29721));
    LocalMux I__4329 (
            .O(N__29721),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_9 ));
    CascadeMux I__4328 (
            .O(N__29718),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_5_cascade_ ));
    CascadeMux I__4327 (
            .O(N__29715),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_4_cascade_ ));
    InMux I__4326 (
            .O(N__29712),
            .I(N__29709));
    LocalMux I__4325 (
            .O(N__29709),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_4 ));
    InMux I__4324 (
            .O(N__29706),
            .I(N__29703));
    LocalMux I__4323 (
            .O(N__29703),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_4 ));
    CascadeMux I__4322 (
            .O(N__29700),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_4_cascade_ ));
    InMux I__4321 (
            .O(N__29697),
            .I(N__29694));
    LocalMux I__4320 (
            .O(N__29694),
            .I(N__29691));
    Span4Mux_v I__4319 (
            .O(N__29691),
            .I(N__29686));
    InMux I__4318 (
            .O(N__29690),
            .I(N__29681));
    InMux I__4317 (
            .O(N__29689),
            .I(N__29681));
    Odrv4 I__4316 (
            .O(N__29686),
            .I(cemf_module_64ch_ctrl_inst1_data_config_4));
    LocalMux I__4315 (
            .O(N__29681),
            .I(cemf_module_64ch_ctrl_inst1_data_config_4));
    CascadeMux I__4314 (
            .O(N__29676),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRLZ0Z7_cascade_ ));
    CascadeMux I__4313 (
            .O(N__29673),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_6_cascade_ ));
    InMux I__4312 (
            .O(N__29670),
            .I(N__29667));
    LocalMux I__4311 (
            .O(N__29667),
            .I(N__29664));
    Odrv12 I__4310 (
            .O(N__29664),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_6 ));
    InMux I__4309 (
            .O(N__29661),
            .I(N__29658));
    LocalMux I__4308 (
            .O(N__29658),
            .I(N__29655));
    Span4Mux_v I__4307 (
            .O(N__29655),
            .I(N__29652));
    Odrv4 I__4306 (
            .O(N__29652),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_775 ));
    CascadeMux I__4305 (
            .O(N__29649),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_15_cascade_ ));
    CascadeMux I__4304 (
            .O(N__29646),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_15_cascade_ ));
    InMux I__4303 (
            .O(N__29643),
            .I(N__29640));
    LocalMux I__4302 (
            .O(N__29640),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_15 ));
    InMux I__4301 (
            .O(N__29637),
            .I(N__29634));
    LocalMux I__4300 (
            .O(N__29634),
            .I(N__29631));
    Span4Mux_v I__4299 (
            .O(N__29631),
            .I(N__29628));
    Span4Mux_h I__4298 (
            .O(N__29628),
            .I(N__29625));
    Odrv4 I__4297 (
            .O(N__29625),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_23));
    InMux I__4296 (
            .O(N__29622),
            .I(N__29619));
    LocalMux I__4295 (
            .O(N__29619),
            .I(N__29616));
    Span4Mux_h I__4294 (
            .O(N__29616),
            .I(N__29613));
    Span4Mux_h I__4293 (
            .O(N__29613),
            .I(N__29610));
    Span4Mux_v I__4292 (
            .O(N__29610),
            .I(N__29607));
    Odrv4 I__4291 (
            .O(N__29607),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_17));
    CascadeMux I__4290 (
            .O(N__29604),
            .I(N__29601));
    InMux I__4289 (
            .O(N__29601),
            .I(N__29598));
    LocalMux I__4288 (
            .O(N__29598),
            .I(N__29595));
    Span4Mux_v I__4287 (
            .O(N__29595),
            .I(N__29592));
    Sp12to4 I__4286 (
            .O(N__29592),
            .I(N__29589));
    Odrv12 I__4285 (
            .O(N__29589),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_17));
    CascadeMux I__4284 (
            .O(N__29586),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_17_cascade_ ));
    InMux I__4283 (
            .O(N__29583),
            .I(N__29580));
    LocalMux I__4282 (
            .O(N__29580),
            .I(N__29577));
    Span4Mux_v I__4281 (
            .O(N__29577),
            .I(N__29574));
    Span4Mux_h I__4280 (
            .O(N__29574),
            .I(N__29571));
    Odrv4 I__4279 (
            .O(N__29571),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_17));
    CascadeMux I__4278 (
            .O(N__29568),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_17_cascade_ ));
    CascadeMux I__4277 (
            .O(N__29565),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_17_cascade_ ));
    InMux I__4276 (
            .O(N__29562),
            .I(N__29559));
    LocalMux I__4275 (
            .O(N__29559),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_17 ));
    InMux I__4274 (
            .O(N__29556),
            .I(N__29553));
    LocalMux I__4273 (
            .O(N__29553),
            .I(N__29550));
    Span4Mux_h I__4272 (
            .O(N__29550),
            .I(N__29547));
    Span4Mux_v I__4271 (
            .O(N__29547),
            .I(N__29544));
    Span4Mux_h I__4270 (
            .O(N__29544),
            .I(N__29541));
    Odrv4 I__4269 (
            .O(N__29541),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_25));
    InMux I__4268 (
            .O(N__29538),
            .I(N__29535));
    LocalMux I__4267 (
            .O(N__29535),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_22 ));
    InMux I__4266 (
            .O(N__29532),
            .I(N__29529));
    LocalMux I__4265 (
            .O(N__29529),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_22 ));
    InMux I__4264 (
            .O(N__29526),
            .I(N__29523));
    LocalMux I__4263 (
            .O(N__29523),
            .I(N__29520));
    Span12Mux_v I__4262 (
            .O(N__29520),
            .I(N__29517));
    Odrv12 I__4261 (
            .O(N__29517),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_28));
    CascadeMux I__4260 (
            .O(N__29514),
            .I(N__29511));
    InMux I__4259 (
            .O(N__29511),
            .I(N__29508));
    LocalMux I__4258 (
            .O(N__29508),
            .I(N__29505));
    Span4Mux_v I__4257 (
            .O(N__29505),
            .I(N__29502));
    Span4Mux_h I__4256 (
            .O(N__29502),
            .I(N__29499));
    Odrv4 I__4255 (
            .O(N__29499),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_28));
    CascadeMux I__4254 (
            .O(N__29496),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_28_cascade_ ));
    InMux I__4253 (
            .O(N__29493),
            .I(N__29490));
    LocalMux I__4252 (
            .O(N__29490),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_28 ));
    CascadeMux I__4251 (
            .O(N__29487),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_28_cascade_ ));
    InMux I__4250 (
            .O(N__29484),
            .I(N__29481));
    LocalMux I__4249 (
            .O(N__29481),
            .I(N__29478));
    Span4Mux_h I__4248 (
            .O(N__29478),
            .I(N__29475));
    Odrv4 I__4247 (
            .O(N__29475),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_28 ));
    InMux I__4246 (
            .O(N__29472),
            .I(N__29469));
    LocalMux I__4245 (
            .O(N__29469),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_28 ));
    InMux I__4244 (
            .O(N__29466),
            .I(N__29463));
    LocalMux I__4243 (
            .O(N__29463),
            .I(N__29460));
    Span4Mux_v I__4242 (
            .O(N__29460),
            .I(N__29457));
    Span4Mux_h I__4241 (
            .O(N__29457),
            .I(N__29454));
    Span4Mux_v I__4240 (
            .O(N__29454),
            .I(N__29451));
    Odrv4 I__4239 (
            .O(N__29451),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_15));
    CascadeMux I__4238 (
            .O(N__29448),
            .I(N__29445));
    InMux I__4237 (
            .O(N__29445),
            .I(N__29442));
    LocalMux I__4236 (
            .O(N__29442),
            .I(N__29439));
    Span4Mux_v I__4235 (
            .O(N__29439),
            .I(N__29436));
    Span4Mux_h I__4234 (
            .O(N__29436),
            .I(N__29433));
    Odrv4 I__4233 (
            .O(N__29433),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_15));
    CascadeMux I__4232 (
            .O(N__29430),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_15_cascade_ ));
    InMux I__4231 (
            .O(N__29427),
            .I(N__29424));
    LocalMux I__4230 (
            .O(N__29424),
            .I(N__29421));
    Span4Mux_h I__4229 (
            .O(N__29421),
            .I(N__29418));
    Span4Mux_h I__4228 (
            .O(N__29418),
            .I(N__29415));
    Odrv4 I__4227 (
            .O(N__29415),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_15));
    InMux I__4226 (
            .O(N__29412),
            .I(N__29409));
    LocalMux I__4225 (
            .O(N__29409),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un40_0_a2_4_a2_0 ));
    InMux I__4224 (
            .O(N__29406),
            .I(N__29402));
    InMux I__4223 (
            .O(N__29405),
            .I(N__29399));
    LocalMux I__4222 (
            .O(N__29402),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0 ));
    LocalMux I__4221 (
            .O(N__29399),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0 ));
    InMux I__4220 (
            .O(N__29394),
            .I(N__29382));
    InMux I__4219 (
            .O(N__29393),
            .I(N__29382));
    InMux I__4218 (
            .O(N__29392),
            .I(N__29382));
    InMux I__4217 (
            .O(N__29391),
            .I(N__29377));
    InMux I__4216 (
            .O(N__29390),
            .I(N__29377));
    InMux I__4215 (
            .O(N__29389),
            .I(N__29374));
    LocalMux I__4214 (
            .O(N__29382),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17 ));
    LocalMux I__4213 (
            .O(N__29377),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17 ));
    LocalMux I__4212 (
            .O(N__29374),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17 ));
    InMux I__4211 (
            .O(N__29367),
            .I(N__29360));
    InMux I__4210 (
            .O(N__29366),
            .I(N__29353));
    InMux I__4209 (
            .O(N__29365),
            .I(N__29353));
    InMux I__4208 (
            .O(N__29364),
            .I(N__29353));
    InMux I__4207 (
            .O(N__29363),
            .I(N__29350));
    LocalMux I__4206 (
            .O(N__29360),
            .I(N__29347));
    LocalMux I__4205 (
            .O(N__29353),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16 ));
    LocalMux I__4204 (
            .O(N__29350),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16 ));
    Odrv4 I__4203 (
            .O(N__29347),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16 ));
    IoInMux I__4202 (
            .O(N__29340),
            .I(N__29337));
    LocalMux I__4201 (
            .O(N__29337),
            .I(N__29334));
    IoSpan4Mux I__4200 (
            .O(N__29334),
            .I(N__29331));
    Span4Mux_s3_h I__4199 (
            .O(N__29331),
            .I(N__29328));
    Span4Mux_h I__4198 (
            .O(N__29328),
            .I(N__29325));
    Span4Mux_h I__4197 (
            .O(N__29325),
            .I(N__29322));
    Odrv4 I__4196 (
            .O(N__29322),
            .I(sda_o));
    CascadeMux I__4195 (
            .O(N__29319),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_22_cascade_ ));
    InMux I__4194 (
            .O(N__29316),
            .I(N__29313));
    LocalMux I__4193 (
            .O(N__29313),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_22 ));
    InMux I__4192 (
            .O(N__29310),
            .I(N__29307));
    LocalMux I__4191 (
            .O(N__29307),
            .I(N__29304));
    Span4Mux_v I__4190 (
            .O(N__29304),
            .I(N__29301));
    Span4Mux_h I__4189 (
            .O(N__29301),
            .I(N__29298));
    Odrv4 I__4188 (
            .O(N__29298),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_22));
    CascadeMux I__4187 (
            .O(N__29295),
            .I(N__29292));
    InMux I__4186 (
            .O(N__29292),
            .I(N__29289));
    LocalMux I__4185 (
            .O(N__29289),
            .I(N__29286));
    Span4Mux_v I__4184 (
            .O(N__29286),
            .I(N__29283));
    Span4Mux_h I__4183 (
            .O(N__29283),
            .I(N__29280));
    Odrv4 I__4182 (
            .O(N__29280),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_22));
    InMux I__4181 (
            .O(N__29277),
            .I(N__29274));
    LocalMux I__4180 (
            .O(N__29274),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_22 ));
    InMux I__4179 (
            .O(N__29271),
            .I(bfn_12_20_0_));
    InMux I__4178 (
            .O(N__29268),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0 ));
    InMux I__4177 (
            .O(N__29265),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1 ));
    InMux I__4176 (
            .O(N__29262),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2 ));
    InMux I__4175 (
            .O(N__29259),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_3 ));
    InMux I__4174 (
            .O(N__29256),
            .I(N__29253));
    LocalMux I__4173 (
            .O(N__29253),
            .I(\cemf_module_64ch_ctrl_inst1.en_ch_cnt_0_a2_0_a2_1 ));
    InMux I__4172 (
            .O(N__29250),
            .I(N__29247));
    LocalMux I__4171 (
            .O(N__29247),
            .I(N__29244));
    Span4Mux_h I__4170 (
            .O(N__29244),
            .I(N__29241));
    Span4Mux_h I__4169 (
            .O(N__29241),
            .I(N__29238));
    Odrv4 I__4168 (
            .O(N__29238),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1867_0 ));
    InMux I__4167 (
            .O(N__29235),
            .I(N__29229));
    InMux I__4166 (
            .O(N__29234),
            .I(N__29229));
    LocalMux I__4165 (
            .O(N__29229),
            .I(N__29226));
    Span4Mux_h I__4164 (
            .O(N__29226),
            .I(N__29216));
    InMux I__4163 (
            .O(N__29225),
            .I(N__29209));
    InMux I__4162 (
            .O(N__29224),
            .I(N__29209));
    InMux I__4161 (
            .O(N__29223),
            .I(N__29209));
    InMux I__4160 (
            .O(N__29222),
            .I(N__29204));
    InMux I__4159 (
            .O(N__29221),
            .I(N__29204));
    InMux I__4158 (
            .O(N__29220),
            .I(N__29199));
    InMux I__4157 (
            .O(N__29219),
            .I(N__29199));
    Odrv4 I__4156 (
            .O(N__29216),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996 ));
    LocalMux I__4155 (
            .O(N__29209),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996 ));
    LocalMux I__4154 (
            .O(N__29204),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996 ));
    LocalMux I__4153 (
            .O(N__29199),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996 ));
    InMux I__4152 (
            .O(N__29190),
            .I(N__29186));
    InMux I__4151 (
            .O(N__29189),
            .I(N__29183));
    LocalMux I__4150 (
            .O(N__29186),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1 ));
    LocalMux I__4149 (
            .O(N__29183),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1 ));
    InMux I__4148 (
            .O(N__29178),
            .I(N__29172));
    InMux I__4147 (
            .O(N__29177),
            .I(N__29172));
    LocalMux I__4146 (
            .O(N__29172),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_13 ));
    InMux I__4145 (
            .O(N__29169),
            .I(N__29157));
    InMux I__4144 (
            .O(N__29168),
            .I(N__29157));
    InMux I__4143 (
            .O(N__29167),
            .I(N__29157));
    InMux I__4142 (
            .O(N__29166),
            .I(N__29157));
    LocalMux I__4141 (
            .O(N__29157),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_12 ));
    InMux I__4140 (
            .O(N__29154),
            .I(N__29151));
    LocalMux I__4139 (
            .O(N__29151),
            .I(N__29148));
    Span4Mux_v I__4138 (
            .O(N__29148),
            .I(N__29142));
    InMux I__4137 (
            .O(N__29147),
            .I(N__29135));
    InMux I__4136 (
            .O(N__29146),
            .I(N__29135));
    InMux I__4135 (
            .O(N__29145),
            .I(N__29135));
    Odrv4 I__4134 (
            .O(N__29142),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4 ));
    LocalMux I__4133 (
            .O(N__29135),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4 ));
    InMux I__4132 (
            .O(N__29130),
            .I(N__29126));
    InMux I__4131 (
            .O(N__29129),
            .I(N__29123));
    LocalMux I__4130 (
            .O(N__29126),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4 ));
    LocalMux I__4129 (
            .O(N__29123),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4 ));
    InMux I__4128 (
            .O(N__29118),
            .I(N__29114));
    InMux I__4127 (
            .O(N__29117),
            .I(N__29111));
    LocalMux I__4126 (
            .O(N__29114),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3 ));
    LocalMux I__4125 (
            .O(N__29111),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3 ));
    InMux I__4124 (
            .O(N__29106),
            .I(N__29103));
    LocalMux I__4123 (
            .O(N__29103),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_i_a2_1_1_3 ));
    InMux I__4122 (
            .O(N__29100),
            .I(N__29096));
    InMux I__4121 (
            .O(N__29099),
            .I(N__29092));
    LocalMux I__4120 (
            .O(N__29096),
            .I(N__29089));
    InMux I__4119 (
            .O(N__29095),
            .I(N__29086));
    LocalMux I__4118 (
            .O(N__29092),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16 ));
    Odrv4 I__4117 (
            .O(N__29089),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16 ));
    LocalMux I__4116 (
            .O(N__29086),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16 ));
    InMux I__4115 (
            .O(N__29079),
            .I(N__29076));
    LocalMux I__4114 (
            .O(N__29076),
            .I(N__29071));
    InMux I__4113 (
            .O(N__29075),
            .I(N__29066));
    InMux I__4112 (
            .O(N__29074),
            .I(N__29066));
    Odrv4 I__4111 (
            .O(N__29071),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8 ));
    LocalMux I__4110 (
            .O(N__29066),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8 ));
    InMux I__4109 (
            .O(N__29061),
            .I(N__29057));
    InMux I__4108 (
            .O(N__29060),
            .I(N__29054));
    LocalMux I__4107 (
            .O(N__29057),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1 ));
    LocalMux I__4106 (
            .O(N__29054),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1 ));
    InMux I__4105 (
            .O(N__29049),
            .I(N__29045));
    InMux I__4104 (
            .O(N__29048),
            .I(N__29042));
    LocalMux I__4103 (
            .O(N__29045),
            .I(N__29038));
    LocalMux I__4102 (
            .O(N__29042),
            .I(N__29034));
    CascadeMux I__4101 (
            .O(N__29041),
            .I(N__29030));
    Span4Mux_h I__4100 (
            .O(N__29038),
            .I(N__29027));
    InMux I__4099 (
            .O(N__29037),
            .I(N__29024));
    Span4Mux_h I__4098 (
            .O(N__29034),
            .I(N__29021));
    InMux I__4097 (
            .O(N__29033),
            .I(N__29016));
    InMux I__4096 (
            .O(N__29030),
            .I(N__29016));
    Odrv4 I__4095 (
            .O(N__29027),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17 ));
    LocalMux I__4094 (
            .O(N__29024),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17 ));
    Odrv4 I__4093 (
            .O(N__29021),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17 ));
    LocalMux I__4092 (
            .O(N__29016),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17 ));
    CascadeMux I__4091 (
            .O(N__29007),
            .I(N__29003));
    CascadeMux I__4090 (
            .O(N__29006),
            .I(N__29000));
    InMux I__4089 (
            .O(N__29003),
            .I(N__28996));
    InMux I__4088 (
            .O(N__29000),
            .I(N__28992));
    InMux I__4087 (
            .O(N__28999),
            .I(N__28989));
    LocalMux I__4086 (
            .O(N__28996),
            .I(N__28986));
    InMux I__4085 (
            .O(N__28995),
            .I(N__28983));
    LocalMux I__4084 (
            .O(N__28992),
            .I(N__28980));
    LocalMux I__4083 (
            .O(N__28989),
            .I(N__28977));
    Span12Mux_v I__4082 (
            .O(N__28986),
            .I(N__28974));
    LocalMux I__4081 (
            .O(N__28983),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5 ));
    Odrv4 I__4080 (
            .O(N__28980),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5 ));
    Odrv4 I__4079 (
            .O(N__28977),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5 ));
    Odrv12 I__4078 (
            .O(N__28974),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5 ));
    InMux I__4077 (
            .O(N__28965),
            .I(N__28962));
    LocalMux I__4076 (
            .O(N__28962),
            .I(N__28959));
    Span4Mux_h I__4075 (
            .O(N__28959),
            .I(N__28953));
    InMux I__4074 (
            .O(N__28958),
            .I(N__28946));
    InMux I__4073 (
            .O(N__28957),
            .I(N__28946));
    InMux I__4072 (
            .O(N__28956),
            .I(N__28946));
    Odrv4 I__4071 (
            .O(N__28953),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9 ));
    LocalMux I__4070 (
            .O(N__28946),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9 ));
    InMux I__4069 (
            .O(N__28941),
            .I(N__28938));
    LocalMux I__4068 (
            .O(N__28938),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_18 ));
    InMux I__4067 (
            .O(N__28935),
            .I(N__28932));
    LocalMux I__4066 (
            .O(N__28932),
            .I(N__28929));
    Span4Mux_v I__4065 (
            .O(N__28929),
            .I(N__28926));
    Span4Mux_h I__4064 (
            .O(N__28926),
            .I(N__28923));
    Odrv4 I__4063 (
            .O(N__28923),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_18 ));
    CascadeMux I__4062 (
            .O(N__28920),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286_cascade_ ));
    InMux I__4061 (
            .O(N__28917),
            .I(N__28914));
    LocalMux I__4060 (
            .O(N__28914),
            .I(N__28911));
    Span4Mux_h I__4059 (
            .O(N__28911),
            .I(N__28905));
    InMux I__4058 (
            .O(N__28910),
            .I(N__28902));
    InMux I__4057 (
            .O(N__28909),
            .I(N__28897));
    InMux I__4056 (
            .O(N__28908),
            .I(N__28897));
    Odrv4 I__4055 (
            .O(N__28905),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3 ));
    LocalMux I__4054 (
            .O(N__28902),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3 ));
    LocalMux I__4053 (
            .O(N__28897),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3 ));
    CascadeMux I__4052 (
            .O(N__28890),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15Z0Z_0_cascade_ ));
    InMux I__4051 (
            .O(N__28887),
            .I(N__28883));
    InMux I__4050 (
            .O(N__28886),
            .I(N__28880));
    LocalMux I__4049 (
            .O(N__28883),
            .I(N__28875));
    LocalMux I__4048 (
            .O(N__28880),
            .I(N__28875));
    Span4Mux_h I__4047 (
            .O(N__28875),
            .I(N__28871));
    InMux I__4046 (
            .O(N__28874),
            .I(N__28868));
    Odrv4 I__4045 (
            .O(N__28871),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7 ));
    LocalMux I__4044 (
            .O(N__28868),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7 ));
    InMux I__4043 (
            .O(N__28863),
            .I(N__28858));
    InMux I__4042 (
            .O(N__28862),
            .I(N__28853));
    InMux I__4041 (
            .O(N__28861),
            .I(N__28853));
    LocalMux I__4040 (
            .O(N__28858),
            .I(N__28850));
    LocalMux I__4039 (
            .O(N__28853),
            .I(N__28844));
    Span4Mux_h I__4038 (
            .O(N__28850),
            .I(N__28841));
    InMux I__4037 (
            .O(N__28849),
            .I(N__28834));
    InMux I__4036 (
            .O(N__28848),
            .I(N__28834));
    InMux I__4035 (
            .O(N__28847),
            .I(N__28834));
    Span4Mux_h I__4034 (
            .O(N__28844),
            .I(N__28831));
    Span4Mux_h I__4033 (
            .O(N__28841),
            .I(N__28826));
    LocalMux I__4032 (
            .O(N__28834),
            .I(N__28826));
    Odrv4 I__4031 (
            .O(N__28831),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0 ));
    Odrv4 I__4030 (
            .O(N__28826),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0 ));
    InMux I__4029 (
            .O(N__28821),
            .I(N__28812));
    InMux I__4028 (
            .O(N__28820),
            .I(N__28812));
    InMux I__4027 (
            .O(N__28819),
            .I(N__28812));
    LocalMux I__4026 (
            .O(N__28812),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_19 ));
    InMux I__4025 (
            .O(N__28809),
            .I(N__28806));
    LocalMux I__4024 (
            .O(N__28806),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_13 ));
    CascadeMux I__4023 (
            .O(N__28803),
            .I(N__28800));
    InMux I__4022 (
            .O(N__28800),
            .I(N__28797));
    LocalMux I__4021 (
            .O(N__28797),
            .I(N__28793));
    InMux I__4020 (
            .O(N__28796),
            .I(N__28790));
    Span12Mux_s9_v I__4019 (
            .O(N__28793),
            .I(N__28787));
    LocalMux I__4018 (
            .O(N__28790),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_8));
    Odrv12 I__4017 (
            .O(N__28787),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_8));
    CascadeMux I__4016 (
            .O(N__28782),
            .I(N__28779));
    InMux I__4015 (
            .O(N__28779),
            .I(N__28776));
    LocalMux I__4014 (
            .O(N__28776),
            .I(N__28773));
    Span4Mux_v I__4013 (
            .O(N__28773),
            .I(N__28770));
    Span4Mux_h I__4012 (
            .O(N__28770),
            .I(N__28767));
    Odrv4 I__4011 (
            .O(N__28767),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_0));
    CascadeMux I__4010 (
            .O(N__28764),
            .I(N__28761));
    InMux I__4009 (
            .O(N__28761),
            .I(N__28758));
    LocalMux I__4008 (
            .O(N__28758),
            .I(N__28755));
    Span12Mux_v I__4007 (
            .O(N__28755),
            .I(N__28752));
    Odrv12 I__4006 (
            .O(N__28752),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_11));
    InMux I__4005 (
            .O(N__28749),
            .I(N__28746));
    LocalMux I__4004 (
            .O(N__28746),
            .I(N__28743));
    Span4Mux_h I__4003 (
            .O(N__28743),
            .I(N__28740));
    Span4Mux_h I__4002 (
            .O(N__28740),
            .I(N__28737));
    Span4Mux_v I__4001 (
            .O(N__28737),
            .I(N__28734));
    Odrv4 I__4000 (
            .O(N__28734),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_12));
    CascadeMux I__3999 (
            .O(N__28731),
            .I(N__28728));
    InMux I__3998 (
            .O(N__28728),
            .I(N__28725));
    LocalMux I__3997 (
            .O(N__28725),
            .I(N__28722));
    Span4Mux_v I__3996 (
            .O(N__28722),
            .I(N__28719));
    Span4Mux_v I__3995 (
            .O(N__28719),
            .I(N__28716));
    Odrv4 I__3994 (
            .O(N__28716),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_13));
    InMux I__3993 (
            .O(N__28713),
            .I(N__28710));
    LocalMux I__3992 (
            .O(N__28710),
            .I(N__28707));
    Span4Mux_v I__3991 (
            .O(N__28707),
            .I(N__28704));
    Span4Mux_v I__3990 (
            .O(N__28704),
            .I(N__28701));
    Odrv4 I__3989 (
            .O(N__28701),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_14));
    InMux I__3988 (
            .O(N__28698),
            .I(N__28695));
    LocalMux I__3987 (
            .O(N__28695),
            .I(N__28692));
    Span4Mux_v I__3986 (
            .O(N__28692),
            .I(N__28689));
    Odrv4 I__3985 (
            .O(N__28689),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_786 ));
    CascadeMux I__3984 (
            .O(N__28686),
            .I(N__28683));
    InMux I__3983 (
            .O(N__28683),
            .I(N__28680));
    LocalMux I__3982 (
            .O(N__28680),
            .I(N__28677));
    Span4Mux_v I__3981 (
            .O(N__28677),
            .I(N__28674));
    Span4Mux_h I__3980 (
            .O(N__28674),
            .I(N__28671));
    Span4Mux_v I__3979 (
            .O(N__28671),
            .I(N__28668));
    Odrv4 I__3978 (
            .O(N__28668),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_15));
    InMux I__3977 (
            .O(N__28665),
            .I(N__28662));
    LocalMux I__3976 (
            .O(N__28662),
            .I(N__28659));
    Odrv12 I__3975 (
            .O(N__28659),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_20));
    CascadeMux I__3974 (
            .O(N__28656),
            .I(N__28653));
    InMux I__3973 (
            .O(N__28653),
            .I(N__28650));
    LocalMux I__3972 (
            .O(N__28650),
            .I(N__28647));
    Span4Mux_v I__3971 (
            .O(N__28647),
            .I(N__28644));
    Span4Mux_h I__3970 (
            .O(N__28644),
            .I(N__28641));
    Span4Mux_v I__3969 (
            .O(N__28641),
            .I(N__28638));
    Odrv4 I__3968 (
            .O(N__28638),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_9));
    InMux I__3967 (
            .O(N__28635),
            .I(N__28632));
    LocalMux I__3966 (
            .O(N__28632),
            .I(N__28629));
    Span12Mux_h I__3965 (
            .O(N__28629),
            .I(N__28626));
    Span12Mux_v I__3964 (
            .O(N__28626),
            .I(N__28623));
    Odrv12 I__3963 (
            .O(N__28623),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_4));
    CascadeMux I__3962 (
            .O(N__28620),
            .I(N__28617));
    InMux I__3961 (
            .O(N__28617),
            .I(N__28614));
    LocalMux I__3960 (
            .O(N__28614),
            .I(N__28611));
    Span4Mux_v I__3959 (
            .O(N__28611),
            .I(N__28608));
    Span4Mux_v I__3958 (
            .O(N__28608),
            .I(N__28605));
    Odrv4 I__3957 (
            .O(N__28605),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_4));
    InMux I__3956 (
            .O(N__28602),
            .I(N__28599));
    LocalMux I__3955 (
            .O(N__28599),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_4 ));
    InMux I__3954 (
            .O(N__28596),
            .I(N__28593));
    LocalMux I__3953 (
            .O(N__28593),
            .I(N__28590));
    Span4Mux_h I__3952 (
            .O(N__28590),
            .I(N__28587));
    Odrv4 I__3951 (
            .O(N__28587),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_9));
    InMux I__3950 (
            .O(N__28584),
            .I(N__28580));
    InMux I__3949 (
            .O(N__28583),
            .I(N__28577));
    LocalMux I__3948 (
            .O(N__28580),
            .I(N__28574));
    LocalMux I__3947 (
            .O(N__28577),
            .I(N__28569));
    Span4Mux_v I__3946 (
            .O(N__28574),
            .I(N__28569));
    Odrv4 I__3945 (
            .O(N__28569),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_30));
    CascadeMux I__3944 (
            .O(N__28566),
            .I(N__28563));
    InMux I__3943 (
            .O(N__28563),
            .I(N__28559));
    CascadeMux I__3942 (
            .O(N__28562),
            .I(N__28556));
    LocalMux I__3941 (
            .O(N__28559),
            .I(N__28553));
    InMux I__3940 (
            .O(N__28556),
            .I(N__28550));
    Span4Mux_v I__3939 (
            .O(N__28553),
            .I(N__28547));
    LocalMux I__3938 (
            .O(N__28550),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_4));
    Odrv4 I__3937 (
            .O(N__28547),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_4));
    InMux I__3936 (
            .O(N__28542),
            .I(N__28539));
    LocalMux I__3935 (
            .O(N__28539),
            .I(N__28536));
    Span4Mux_h I__3934 (
            .O(N__28536),
            .I(N__28533));
    Span4Mux_v I__3933 (
            .O(N__28533),
            .I(N__28530));
    Odrv4 I__3932 (
            .O(N__28530),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_9));
    InMux I__3931 (
            .O(N__28527),
            .I(N__28524));
    LocalMux I__3930 (
            .O(N__28524),
            .I(N__28521));
    Span4Mux_v I__3929 (
            .O(N__28521),
            .I(N__28518));
    Span4Mux_h I__3928 (
            .O(N__28518),
            .I(N__28515));
    Odrv4 I__3927 (
            .O(N__28515),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_29));
    InMux I__3926 (
            .O(N__28512),
            .I(N__28509));
    LocalMux I__3925 (
            .O(N__28509),
            .I(N__28506));
    Span4Mux_h I__3924 (
            .O(N__28506),
            .I(N__28503));
    Odrv4 I__3923 (
            .O(N__28503),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_3));
    CascadeMux I__3922 (
            .O(N__28500),
            .I(N__28497));
    InMux I__3921 (
            .O(N__28497),
            .I(N__28494));
    LocalMux I__3920 (
            .O(N__28494),
            .I(N__28491));
    Odrv4 I__3919 (
            .O(N__28491),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_907 ));
    CascadeMux I__3918 (
            .O(N__28488),
            .I(N__28485));
    InMux I__3917 (
            .O(N__28485),
            .I(N__28482));
    LocalMux I__3916 (
            .O(N__28482),
            .I(N__28479));
    Span4Mux_h I__3915 (
            .O(N__28479),
            .I(N__28476));
    Span4Mux_h I__3914 (
            .O(N__28476),
            .I(N__28473));
    Odrv4 I__3913 (
            .O(N__28473),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_30));
    InMux I__3912 (
            .O(N__28470),
            .I(N__28467));
    LocalMux I__3911 (
            .O(N__28467),
            .I(N__28464));
    Odrv4 I__3910 (
            .O(N__28464),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_621 ));
    InMux I__3909 (
            .O(N__28461),
            .I(N__28458));
    LocalMux I__3908 (
            .O(N__28458),
            .I(N__28455));
    Span4Mux_h I__3907 (
            .O(N__28455),
            .I(N__28452));
    Odrv4 I__3906 (
            .O(N__28452),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_31));
    InMux I__3905 (
            .O(N__28449),
            .I(N__28446));
    LocalMux I__3904 (
            .O(N__28446),
            .I(N__28443));
    Span4Mux_h I__3903 (
            .O(N__28443),
            .I(N__28440));
    Odrv4 I__3902 (
            .O(N__28440),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_610 ));
    CascadeMux I__3901 (
            .O(N__28437),
            .I(N__28434));
    InMux I__3900 (
            .O(N__28434),
            .I(N__28431));
    LocalMux I__3899 (
            .O(N__28431),
            .I(N__28428));
    Span4Mux_h I__3898 (
            .O(N__28428),
            .I(N__28425));
    Odrv4 I__3897 (
            .O(N__28425),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_1));
    InMux I__3896 (
            .O(N__28422),
            .I(N__28419));
    LocalMux I__3895 (
            .O(N__28419),
            .I(N__28416));
    Span4Mux_v I__3894 (
            .O(N__28416),
            .I(N__28413));
    Odrv4 I__3893 (
            .O(N__28413),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316 ));
    InMux I__3892 (
            .O(N__28410),
            .I(N__28407));
    LocalMux I__3891 (
            .O(N__28407),
            .I(N__28404));
    Span4Mux_v I__3890 (
            .O(N__28404),
            .I(N__28401));
    Span4Mux_h I__3889 (
            .O(N__28401),
            .I(N__28398));
    Sp12to4 I__3888 (
            .O(N__28398),
            .I(N__28395));
    Odrv12 I__3887 (
            .O(N__28395),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_5));
    CascadeMux I__3886 (
            .O(N__28392),
            .I(N__28389));
    InMux I__3885 (
            .O(N__28389),
            .I(N__28386));
    LocalMux I__3884 (
            .O(N__28386),
            .I(N__28383));
    Span4Mux_h I__3883 (
            .O(N__28383),
            .I(N__28380));
    Odrv4 I__3882 (
            .O(N__28380),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_885 ));
    CascadeMux I__3881 (
            .O(N__28377),
            .I(N__28374));
    InMux I__3880 (
            .O(N__28374),
            .I(N__28371));
    LocalMux I__3879 (
            .O(N__28371),
            .I(N__28368));
    Span4Mux_v I__3878 (
            .O(N__28368),
            .I(N__28365));
    Span4Mux_h I__3877 (
            .O(N__28365),
            .I(N__28362));
    Odrv4 I__3876 (
            .O(N__28362),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_6));
    CascadeMux I__3875 (
            .O(N__28359),
            .I(N__28356));
    InMux I__3874 (
            .O(N__28356),
            .I(N__28353));
    LocalMux I__3873 (
            .O(N__28353),
            .I(N__28350));
    Odrv4 I__3872 (
            .O(N__28350),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_874 ));
    InMux I__3871 (
            .O(N__28347),
            .I(N__28344));
    LocalMux I__3870 (
            .O(N__28344),
            .I(N__28341));
    Span4Mux_v I__3869 (
            .O(N__28341),
            .I(N__28338));
    Span4Mux_h I__3868 (
            .O(N__28338),
            .I(N__28335));
    Span4Mux_v I__3867 (
            .O(N__28335),
            .I(N__28332));
    Span4Mux_v I__3866 (
            .O(N__28332),
            .I(N__28329));
    Odrv4 I__3865 (
            .O(N__28329),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_9));
    CascadeMux I__3864 (
            .O(N__28326),
            .I(N__28322));
    InMux I__3863 (
            .O(N__28325),
            .I(N__28314));
    InMux I__3862 (
            .O(N__28322),
            .I(N__28314));
    InMux I__3861 (
            .O(N__28321),
            .I(N__28314));
    LocalMux I__3860 (
            .O(N__28314),
            .I(cemf_module_64ch_ctrl_inst1_data_clkstopmask_4));
    InMux I__3859 (
            .O(N__28311),
            .I(N__28308));
    LocalMux I__3858 (
            .O(N__28308),
            .I(N__28305));
    Span4Mux_v I__3857 (
            .O(N__28305),
            .I(N__28302));
    Odrv4 I__3856 (
            .O(N__28302),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_26));
    InMux I__3855 (
            .O(N__28299),
            .I(N__28296));
    LocalMux I__3854 (
            .O(N__28296),
            .I(N__28293));
    Span4Mux_v I__3853 (
            .O(N__28293),
            .I(N__28290));
    Span4Mux_h I__3852 (
            .O(N__28290),
            .I(N__28287));
    Span4Mux_v I__3851 (
            .O(N__28287),
            .I(N__28284));
    Odrv4 I__3850 (
            .O(N__28284),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_26));
    CascadeMux I__3849 (
            .O(N__28281),
            .I(N__28278));
    InMux I__3848 (
            .O(N__28278),
            .I(N__28275));
    LocalMux I__3847 (
            .O(N__28275),
            .I(N__28272));
    Span4Mux_v I__3846 (
            .O(N__28272),
            .I(N__28269));
    Span4Mux_h I__3845 (
            .O(N__28269),
            .I(N__28266));
    Odrv4 I__3844 (
            .O(N__28266),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_26));
    InMux I__3843 (
            .O(N__28263),
            .I(N__28260));
    LocalMux I__3842 (
            .O(N__28260),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_0_26 ));
    CascadeMux I__3841 (
            .O(N__28257),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_1_26_cascade_ ));
    InMux I__3840 (
            .O(N__28254),
            .I(N__28251));
    LocalMux I__3839 (
            .O(N__28251),
            .I(N__28248));
    Span12Mux_h I__3838 (
            .O(N__28248),
            .I(N__28245));
    Odrv12 I__3837 (
            .O(N__28245),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_26));
    InMux I__3836 (
            .O(N__28242),
            .I(N__28239));
    LocalMux I__3835 (
            .O(N__28239),
            .I(N__28236));
    Span4Mux_h I__3834 (
            .O(N__28236),
            .I(N__28233));
    Span4Mux_h I__3833 (
            .O(N__28233),
            .I(N__28230));
    Odrv4 I__3832 (
            .O(N__28230),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_21));
    CascadeMux I__3831 (
            .O(N__28227),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_30_cascade_ ));
    InMux I__3830 (
            .O(N__28224),
            .I(N__28221));
    LocalMux I__3829 (
            .O(N__28221),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_30 ));
    CascadeMux I__3828 (
            .O(N__28218),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_30_cascade_ ));
    InMux I__3827 (
            .O(N__28215),
            .I(N__28212));
    LocalMux I__3826 (
            .O(N__28212),
            .I(N__28209));
    Odrv4 I__3825 (
            .O(N__28209),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_30 ));
    InMux I__3824 (
            .O(N__28206),
            .I(N__28203));
    LocalMux I__3823 (
            .O(N__28203),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_30 ));
    InMux I__3822 (
            .O(N__28200),
            .I(N__28197));
    LocalMux I__3821 (
            .O(N__28197),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_30 ));
    CascadeMux I__3820 (
            .O(N__28194),
            .I(N__28191));
    InMux I__3819 (
            .O(N__28191),
            .I(N__28188));
    LocalMux I__3818 (
            .O(N__28188),
            .I(N__28185));
    Odrv4 I__3817 (
            .O(N__28185),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_30));
    InMux I__3816 (
            .O(N__28182),
            .I(N__28178));
    InMux I__3815 (
            .O(N__28181),
            .I(N__28175));
    LocalMux I__3814 (
            .O(N__28178),
            .I(N__28171));
    LocalMux I__3813 (
            .O(N__28175),
            .I(N__28168));
    InMux I__3812 (
            .O(N__28174),
            .I(N__28165));
    Span4Mux_v I__3811 (
            .O(N__28171),
            .I(N__28162));
    Span12Mux_v I__3810 (
            .O(N__28168),
            .I(N__28159));
    LocalMux I__3809 (
            .O(N__28165),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_31));
    Odrv4 I__3808 (
            .O(N__28162),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_31));
    Odrv12 I__3807 (
            .O(N__28159),
            .I(cemf_module_64ch_ctrl_inst1_s_data_system_o_31));
    InMux I__3806 (
            .O(N__28152),
            .I(N__28149));
    LocalMux I__3805 (
            .O(N__28149),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_31 ));
    CascadeMux I__3804 (
            .O(N__28146),
            .I(N__28143));
    InMux I__3803 (
            .O(N__28143),
            .I(N__28140));
    LocalMux I__3802 (
            .O(N__28140),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_31));
    InMux I__3801 (
            .O(N__28137),
            .I(N__28134));
    LocalMux I__3800 (
            .O(N__28134),
            .I(N__28131));
    Span4Mux_v I__3799 (
            .O(N__28131),
            .I(N__28128));
    Odrv4 I__3798 (
            .O(N__28128),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_4 ));
    InMux I__3797 (
            .O(N__28125),
            .I(N__28122));
    LocalMux I__3796 (
            .O(N__28122),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_8 ));
    InMux I__3795 (
            .O(N__28119),
            .I(N__28116));
    LocalMux I__3794 (
            .O(N__28116),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_8 ));
    CascadeMux I__3793 (
            .O(N__28113),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_8_cascade_ ));
    InMux I__3792 (
            .O(N__28110),
            .I(N__28107));
    LocalMux I__3791 (
            .O(N__28107),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_8 ));
    InMux I__3790 (
            .O(N__28104),
            .I(N__28101));
    LocalMux I__3789 (
            .O(N__28101),
            .I(N__28098));
    Span4Mux_v I__3788 (
            .O(N__28098),
            .I(N__28095));
    Span4Mux_v I__3787 (
            .O(N__28095),
            .I(N__28092));
    Odrv4 I__3786 (
            .O(N__28092),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_14));
    CascadeMux I__3785 (
            .O(N__28089),
            .I(N__28086));
    InMux I__3784 (
            .O(N__28086),
            .I(N__28083));
    LocalMux I__3783 (
            .O(N__28083),
            .I(N__28080));
    Span4Mux_v I__3782 (
            .O(N__28080),
            .I(N__28077));
    Span4Mux_h I__3781 (
            .O(N__28077),
            .I(N__28074));
    Odrv4 I__3780 (
            .O(N__28074),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_14));
    CascadeMux I__3779 (
            .O(N__28071),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_14_cascade_ ));
    InMux I__3778 (
            .O(N__28068),
            .I(N__28065));
    LocalMux I__3777 (
            .O(N__28065),
            .I(N__28062));
    Span4Mux_h I__3776 (
            .O(N__28062),
            .I(N__28059));
    Span4Mux_v I__3775 (
            .O(N__28059),
            .I(N__28056));
    Odrv4 I__3774 (
            .O(N__28056),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_14));
    CascadeMux I__3773 (
            .O(N__28053),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_14_cascade_ ));
    CascadeMux I__3772 (
            .O(N__28050),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_14_cascade_ ));
    InMux I__3771 (
            .O(N__28047),
            .I(N__28044));
    LocalMux I__3770 (
            .O(N__28044),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_14 ));
    InMux I__3769 (
            .O(N__28041),
            .I(N__28038));
    LocalMux I__3768 (
            .O(N__28038),
            .I(N__28035));
    Span4Mux_h I__3767 (
            .O(N__28035),
            .I(N__28032));
    Span4Mux_v I__3766 (
            .O(N__28032),
            .I(N__28029));
    Odrv4 I__3765 (
            .O(N__28029),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_22));
    InMux I__3764 (
            .O(N__28026),
            .I(N__28023));
    LocalMux I__3763 (
            .O(N__28023),
            .I(N__28020));
    Span4Mux_v I__3762 (
            .O(N__28020),
            .I(N__28017));
    Span4Mux_v I__3761 (
            .O(N__28017),
            .I(N__28014));
    Odrv4 I__3760 (
            .O(N__28014),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_30));
    CascadeMux I__3759 (
            .O(N__28011),
            .I(N__28008));
    InMux I__3758 (
            .O(N__28008),
            .I(N__28005));
    LocalMux I__3757 (
            .O(N__28005),
            .I(N__28002));
    Span4Mux_v I__3756 (
            .O(N__28002),
            .I(N__27999));
    Odrv4 I__3755 (
            .O(N__27999),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_30));
    InMux I__3754 (
            .O(N__27996),
            .I(N__27993));
    LocalMux I__3753 (
            .O(N__27993),
            .I(N__27990));
    Span4Mux_v I__3752 (
            .O(N__27990),
            .I(N__27987));
    Span4Mux_v I__3751 (
            .O(N__27987),
            .I(N__27984));
    IoSpan4Mux I__3750 (
            .O(N__27984),
            .I(N__27981));
    Odrv4 I__3749 (
            .O(N__27981),
            .I(sync_50hz_c));
    InMux I__3748 (
            .O(N__27978),
            .I(N__27974));
    InMux I__3747 (
            .O(N__27977),
            .I(N__27971));
    LocalMux I__3746 (
            .O(N__27974),
            .I(\cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0 ));
    LocalMux I__3745 (
            .O(N__27971),
            .I(\cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0 ));
    InMux I__3744 (
            .O(N__27966),
            .I(N__27962));
    InMux I__3743 (
            .O(N__27965),
            .I(N__27959));
    LocalMux I__3742 (
            .O(N__27962),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config ));
    LocalMux I__3741 (
            .O(N__27959),
            .I(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config ));
    CascadeMux I__3740 (
            .O(N__27954),
            .I(\cemf_module_64ch_ctrl_inst1.N_410_0_cascade_ ));
    CascadeMux I__3739 (
            .O(N__27951),
            .I(\cemf_module_64ch_ctrl_inst1.N_68_0_cascade_ ));
    InMux I__3738 (
            .O(N__27948),
            .I(N__27945));
    LocalMux I__3737 (
            .O(N__27945),
            .I(N__27942));
    Span4Mux_v I__3736 (
            .O(N__27942),
            .I(N__27939));
    Span4Mux_h I__3735 (
            .O(N__27939),
            .I(N__27936));
    Odrv4 I__3734 (
            .O(N__27936),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_8));
    CascadeMux I__3733 (
            .O(N__27933),
            .I(N__27930));
    InMux I__3732 (
            .O(N__27930),
            .I(N__27927));
    LocalMux I__3731 (
            .O(N__27927),
            .I(N__27924));
    Span4Mux_v I__3730 (
            .O(N__27924),
            .I(N__27921));
    Span4Mux_h I__3729 (
            .O(N__27921),
            .I(N__27918));
    Odrv4 I__3728 (
            .O(N__27918),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_8));
    CascadeMux I__3727 (
            .O(N__27915),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_8_cascade_ ));
    InMux I__3726 (
            .O(N__27912),
            .I(N__27908));
    InMux I__3725 (
            .O(N__27911),
            .I(N__27905));
    LocalMux I__3724 (
            .O(N__27908),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2 ));
    LocalMux I__3723 (
            .O(N__27905),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2 ));
    InMux I__3722 (
            .O(N__27900),
            .I(N__27897));
    LocalMux I__3721 (
            .O(N__27897),
            .I(N__27894));
    Span4Mux_h I__3720 (
            .O(N__27894),
            .I(N__27891));
    Odrv4 I__3719 (
            .O(N__27891),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_1 ));
    CascadeMux I__3718 (
            .O(N__27888),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287_cascade_ ));
    InMux I__3717 (
            .O(N__27885),
            .I(N__27881));
    InMux I__3716 (
            .O(N__27884),
            .I(N__27878));
    LocalMux I__3715 (
            .O(N__27881),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0 ));
    LocalMux I__3714 (
            .O(N__27878),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0 ));
    InMux I__3713 (
            .O(N__27873),
            .I(bfn_11_19_0_));
    InMux I__3712 (
            .O(N__27870),
            .I(N__27866));
    InMux I__3711 (
            .O(N__27869),
            .I(N__27863));
    LocalMux I__3710 (
            .O(N__27866),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1 ));
    LocalMux I__3709 (
            .O(N__27863),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1 ));
    InMux I__3708 (
            .O(N__27858),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0 ));
    CascadeMux I__3707 (
            .O(N__27855),
            .I(N__27851));
    InMux I__3706 (
            .O(N__27854),
            .I(N__27848));
    InMux I__3705 (
            .O(N__27851),
            .I(N__27845));
    LocalMux I__3704 (
            .O(N__27848),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2 ));
    LocalMux I__3703 (
            .O(N__27845),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2 ));
    InMux I__3702 (
            .O(N__27840),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1 ));
    InMux I__3701 (
            .O(N__27837),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2 ));
    InMux I__3700 (
            .O(N__27834),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_3 ));
    InMux I__3699 (
            .O(N__27831),
            .I(N__27828));
    LocalMux I__3698 (
            .O(N__27828),
            .I(N__27824));
    CascadeMux I__3697 (
            .O(N__27827),
            .I(N__27818));
    Span4Mux_v I__3696 (
            .O(N__27824),
            .I(N__27814));
    InMux I__3695 (
            .O(N__27823),
            .I(N__27803));
    InMux I__3694 (
            .O(N__27822),
            .I(N__27803));
    InMux I__3693 (
            .O(N__27821),
            .I(N__27803));
    InMux I__3692 (
            .O(N__27818),
            .I(N__27803));
    InMux I__3691 (
            .O(N__27817),
            .I(N__27803));
    Odrv4 I__3690 (
            .O(N__27814),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0 ));
    LocalMux I__3689 (
            .O(N__27803),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0 ));
    CascadeMux I__3688 (
            .O(N__27798),
            .I(N__27795));
    InMux I__3687 (
            .O(N__27795),
            .I(N__27792));
    LocalMux I__3686 (
            .O(N__27792),
            .I(N__27789));
    Span4Mux_v I__3685 (
            .O(N__27789),
            .I(N__27765));
    InMux I__3684 (
            .O(N__27788),
            .I(N__27762));
    InMux I__3683 (
            .O(N__27787),
            .I(N__27745));
    InMux I__3682 (
            .O(N__27786),
            .I(N__27745));
    InMux I__3681 (
            .O(N__27785),
            .I(N__27745));
    InMux I__3680 (
            .O(N__27784),
            .I(N__27745));
    InMux I__3679 (
            .O(N__27783),
            .I(N__27745));
    InMux I__3678 (
            .O(N__27782),
            .I(N__27745));
    InMux I__3677 (
            .O(N__27781),
            .I(N__27745));
    InMux I__3676 (
            .O(N__27780),
            .I(N__27745));
    InMux I__3675 (
            .O(N__27779),
            .I(N__27728));
    InMux I__3674 (
            .O(N__27778),
            .I(N__27728));
    InMux I__3673 (
            .O(N__27777),
            .I(N__27728));
    InMux I__3672 (
            .O(N__27776),
            .I(N__27728));
    InMux I__3671 (
            .O(N__27775),
            .I(N__27728));
    InMux I__3670 (
            .O(N__27774),
            .I(N__27728));
    InMux I__3669 (
            .O(N__27773),
            .I(N__27728));
    InMux I__3668 (
            .O(N__27772),
            .I(N__27728));
    InMux I__3667 (
            .O(N__27771),
            .I(N__27719));
    InMux I__3666 (
            .O(N__27770),
            .I(N__27719));
    InMux I__3665 (
            .O(N__27769),
            .I(N__27719));
    InMux I__3664 (
            .O(N__27768),
            .I(N__27719));
    Odrv4 I__3663 (
            .O(N__27765),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ));
    LocalMux I__3662 (
            .O(N__27762),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ));
    LocalMux I__3661 (
            .O(N__27745),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ));
    LocalMux I__3660 (
            .O(N__27728),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ));
    LocalMux I__3659 (
            .O(N__27719),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ));
    CEMux I__3658 (
            .O(N__27708),
            .I(N__27704));
    CEMux I__3657 (
            .O(N__27707),
            .I(N__27701));
    LocalMux I__3656 (
            .O(N__27704),
            .I(N__27698));
    LocalMux I__3655 (
            .O(N__27701),
            .I(N__27695));
    Odrv4 I__3654 (
            .O(N__27698),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i ));
    Odrv4 I__3653 (
            .O(N__27695),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i ));
    CascadeMux I__3652 (
            .O(N__27690),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996_cascade_ ));
    InMux I__3651 (
            .O(N__27687),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1 ));
    InMux I__3650 (
            .O(N__27684),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2 ));
    InMux I__3649 (
            .O(N__27681),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_3 ));
    InMux I__3648 (
            .O(N__27678),
            .I(N__27675));
    LocalMux I__3647 (
            .O(N__27675),
            .I(N__27672));
    Span4Mux_h I__3646 (
            .O(N__27672),
            .I(N__27669));
    Odrv4 I__3645 (
            .O(N__27669),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2 ));
    InMux I__3644 (
            .O(N__27666),
            .I(N__27662));
    InMux I__3643 (
            .O(N__27665),
            .I(N__27659));
    LocalMux I__3642 (
            .O(N__27662),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4 ));
    LocalMux I__3641 (
            .O(N__27659),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4 ));
    InMux I__3640 (
            .O(N__27654),
            .I(N__27650));
    InMux I__3639 (
            .O(N__27653),
            .I(N__27647));
    LocalMux I__3638 (
            .O(N__27650),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2 ));
    LocalMux I__3637 (
            .O(N__27647),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2 ));
    CascadeMux I__3636 (
            .O(N__27642),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2_cascade_ ));
    InMux I__3635 (
            .O(N__27639),
            .I(N__27635));
    InMux I__3634 (
            .O(N__27638),
            .I(N__27632));
    LocalMux I__3633 (
            .O(N__27635),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1 ));
    LocalMux I__3632 (
            .O(N__27632),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1 ));
    InMux I__3631 (
            .O(N__27627),
            .I(N__27623));
    InMux I__3630 (
            .O(N__27626),
            .I(N__27620));
    LocalMux I__3629 (
            .O(N__27623),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3 ));
    LocalMux I__3628 (
            .O(N__27620),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3 ));
    CascadeMux I__3627 (
            .O(N__27615),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m7_3_cascade_ ));
    InMux I__3626 (
            .O(N__27612),
            .I(N__27608));
    InMux I__3625 (
            .O(N__27611),
            .I(N__27605));
    LocalMux I__3624 (
            .O(N__27608),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0 ));
    LocalMux I__3623 (
            .O(N__27605),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0 ));
    InMux I__3622 (
            .O(N__27600),
            .I(N__27591));
    InMux I__3621 (
            .O(N__27599),
            .I(N__27591));
    InMux I__3620 (
            .O(N__27598),
            .I(N__27584));
    InMux I__3619 (
            .O(N__27597),
            .I(N__27584));
    InMux I__3618 (
            .O(N__27596),
            .I(N__27584));
    LocalMux I__3617 (
            .O(N__27591),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2 ));
    LocalMux I__3616 (
            .O(N__27584),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2 ));
    InMux I__3615 (
            .O(N__27579),
            .I(N__27573));
    InMux I__3614 (
            .O(N__27578),
            .I(N__27573));
    LocalMux I__3613 (
            .O(N__27573),
            .I(N__27569));
    InMux I__3612 (
            .O(N__27572),
            .I(N__27564));
    Span4Mux_v I__3611 (
            .O(N__27569),
            .I(N__27561));
    InMux I__3610 (
            .O(N__27568),
            .I(N__27556));
    InMux I__3609 (
            .O(N__27567),
            .I(N__27556));
    LocalMux I__3608 (
            .O(N__27564),
            .I(N__27553));
    Sp12to4 I__3607 (
            .O(N__27561),
            .I(N__27548));
    LocalMux I__3606 (
            .O(N__27556),
            .I(N__27548));
    Span4Mux_v I__3605 (
            .O(N__27553),
            .I(N__27545));
    Odrv12 I__3604 (
            .O(N__27548),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46 ));
    Odrv4 I__3603 (
            .O(N__27545),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46 ));
    InMux I__3602 (
            .O(N__27540),
            .I(N__27537));
    LocalMux I__3601 (
            .O(N__27537),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_3 ));
    CascadeMux I__3600 (
            .O(N__27534),
            .I(N__27531));
    InMux I__3599 (
            .O(N__27531),
            .I(N__27528));
    LocalMux I__3598 (
            .O(N__27528),
            .I(N__27525));
    Span4Mux_h I__3597 (
            .O(N__27525),
            .I(N__27522));
    Odrv4 I__3596 (
            .O(N__27522),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_3));
    InMux I__3595 (
            .O(N__27519),
            .I(N__27516));
    LocalMux I__3594 (
            .O(N__27516),
            .I(N__27513));
    Odrv4 I__3593 (
            .O(N__27513),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3 ));
    InMux I__3592 (
            .O(N__27510),
            .I(N__27507));
    LocalMux I__3591 (
            .O(N__27507),
            .I(N__27504));
    Span4Mux_h I__3590 (
            .O(N__27504),
            .I(N__27501));
    Odrv4 I__3589 (
            .O(N__27501),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_4));
    CascadeMux I__3588 (
            .O(N__27498),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_cascade_ ));
    InMux I__3587 (
            .O(N__27495),
            .I(N__27492));
    LocalMux I__3586 (
            .O(N__27492),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_5 ));
    InMux I__3585 (
            .O(N__27489),
            .I(N__27486));
    LocalMux I__3584 (
            .O(N__27486),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_4 ));
    CascadeMux I__3583 (
            .O(N__27483),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_4_cascade_ ));
    InMux I__3582 (
            .O(N__27480),
            .I(N__27477));
    LocalMux I__3581 (
            .O(N__27477),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_4 ));
    InMux I__3580 (
            .O(N__27474),
            .I(bfn_11_15_0_));
    InMux I__3579 (
            .O(N__27471),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0 ));
    CascadeMux I__3578 (
            .O(N__27468),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_31_cascade_ ));
    InMux I__3577 (
            .O(N__27465),
            .I(N__27462));
    LocalMux I__3576 (
            .O(N__27462),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_31 ));
    CascadeMux I__3575 (
            .O(N__27459),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_31_cascade_ ));
    InMux I__3574 (
            .O(N__27456),
            .I(N__27453));
    LocalMux I__3573 (
            .O(N__27453),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_31 ));
    InMux I__3572 (
            .O(N__27450),
            .I(N__27447));
    LocalMux I__3571 (
            .O(N__27447),
            .I(N__27444));
    Span4Mux_v I__3570 (
            .O(N__27444),
            .I(N__27441));
    Odrv4 I__3569 (
            .O(N__27441),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_27));
    InMux I__3568 (
            .O(N__27438),
            .I(N__27435));
    LocalMux I__3567 (
            .O(N__27435),
            .I(N__27432));
    Span4Mux_h I__3566 (
            .O(N__27432),
            .I(N__27429));
    Odrv4 I__3565 (
            .O(N__27429),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_28));
    InMux I__3564 (
            .O(N__27426),
            .I(N__27423));
    LocalMux I__3563 (
            .O(N__27423),
            .I(N__27420));
    Span4Mux_h I__3562 (
            .O(N__27420),
            .I(N__27417));
    Odrv4 I__3561 (
            .O(N__27417),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_29));
    InMux I__3560 (
            .O(N__27414),
            .I(N__27411));
    LocalMux I__3559 (
            .O(N__27411),
            .I(N__27408));
    Span4Mux_v I__3558 (
            .O(N__27408),
            .I(N__27405));
    Odrv4 I__3557 (
            .O(N__27405),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_30));
    InMux I__3556 (
            .O(N__27402),
            .I(N__27399));
    LocalMux I__3555 (
            .O(N__27399),
            .I(N__27396));
    Span4Mux_h I__3554 (
            .O(N__27396),
            .I(N__27393));
    Odrv4 I__3553 (
            .O(N__27393),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_31));
    InMux I__3552 (
            .O(N__27390),
            .I(N__27387));
    LocalMux I__3551 (
            .O(N__27387),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_31 ));
    InMux I__3550 (
            .O(N__27384),
            .I(N__27381));
    LocalMux I__3549 (
            .O(N__27381),
            .I(N__27378));
    Span4Mux_v I__3548 (
            .O(N__27378),
            .I(N__27375));
    Odrv4 I__3547 (
            .O(N__27375),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_1 ));
    CascadeMux I__3546 (
            .O(N__27372),
            .I(N__27369));
    InMux I__3545 (
            .O(N__27369),
            .I(N__27366));
    LocalMux I__3544 (
            .O(N__27366),
            .I(N__27363));
    Odrv4 I__3543 (
            .O(N__27363),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_10));
    CascadeMux I__3542 (
            .O(N__27360),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_3_cascade_ ));
    InMux I__3541 (
            .O(N__27357),
            .I(N__27354));
    LocalMux I__3540 (
            .O(N__27354),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_3 ));
    InMux I__3539 (
            .O(N__27351),
            .I(N__27348));
    LocalMux I__3538 (
            .O(N__27348),
            .I(N__27345));
    Span4Mux_v I__3537 (
            .O(N__27345),
            .I(N__27342));
    Span4Mux_v I__3536 (
            .O(N__27342),
            .I(N__27339));
    Odrv4 I__3535 (
            .O(N__27339),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_3));
    CascadeMux I__3534 (
            .O(N__27336),
            .I(N__27333));
    InMux I__3533 (
            .O(N__27333),
            .I(N__27330));
    LocalMux I__3532 (
            .O(N__27330),
            .I(N__27327));
    Span12Mux_h I__3531 (
            .O(N__27327),
            .I(N__27324));
    Odrv12 I__3530 (
            .O(N__27324),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_3));
    CascadeMux I__3529 (
            .O(N__27321),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_3_cascade_ ));
    InMux I__3528 (
            .O(N__27318),
            .I(N__27315));
    LocalMux I__3527 (
            .O(N__27315),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_3 ));
    InMux I__3526 (
            .O(N__27312),
            .I(N__27309));
    LocalMux I__3525 (
            .O(N__27309),
            .I(N__27306));
    Span12Mux_h I__3524 (
            .O(N__27306),
            .I(N__27303));
    Odrv12 I__3523 (
            .O(N__27303),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_31));
    CascadeMux I__3522 (
            .O(N__27300),
            .I(N__27297));
    InMux I__3521 (
            .O(N__27297),
            .I(N__27294));
    LocalMux I__3520 (
            .O(N__27294),
            .I(N__27291));
    Span4Mux_v I__3519 (
            .O(N__27291),
            .I(N__27288));
    Odrv4 I__3518 (
            .O(N__27288),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_31));
    InMux I__3517 (
            .O(N__27285),
            .I(N__27282));
    LocalMux I__3516 (
            .O(N__27282),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_18 ));
    InMux I__3515 (
            .O(N__27279),
            .I(N__27276));
    LocalMux I__3514 (
            .O(N__27276),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_19 ));
    InMux I__3513 (
            .O(N__27273),
            .I(N__27270));
    LocalMux I__3512 (
            .O(N__27270),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_16 ));
    InMux I__3511 (
            .O(N__27267),
            .I(N__27264));
    LocalMux I__3510 (
            .O(N__27264),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_17 ));
    InMux I__3509 (
            .O(N__27261),
            .I(N__27258));
    LocalMux I__3508 (
            .O(N__27258),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_11 ));
    InMux I__3507 (
            .O(N__27255),
            .I(N__27252));
    LocalMux I__3506 (
            .O(N__27252),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_8 ));
    InMux I__3505 (
            .O(N__27249),
            .I(N__27246));
    LocalMux I__3504 (
            .O(N__27246),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_9 ));
    InMux I__3503 (
            .O(N__27243),
            .I(N__27240));
    LocalMux I__3502 (
            .O(N__27240),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_10 ));
    CEMux I__3501 (
            .O(N__27237),
            .I(N__27232));
    CEMux I__3500 (
            .O(N__27236),
            .I(N__27229));
    CEMux I__3499 (
            .O(N__27235),
            .I(N__27226));
    LocalMux I__3498 (
            .O(N__27232),
            .I(N__27223));
    LocalMux I__3497 (
            .O(N__27229),
            .I(N__27220));
    LocalMux I__3496 (
            .O(N__27226),
            .I(N__27217));
    Odrv4 I__3495 (
            .O(N__27223),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i ));
    Odrv4 I__3494 (
            .O(N__27220),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i ));
    Odrv4 I__3493 (
            .O(N__27217),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i ));
    InMux I__3492 (
            .O(N__27210),
            .I(N__27204));
    InMux I__3491 (
            .O(N__27209),
            .I(N__27199));
    InMux I__3490 (
            .O(N__27208),
            .I(N__27199));
    InMux I__3489 (
            .O(N__27207),
            .I(N__27196));
    LocalMux I__3488 (
            .O(N__27204),
            .I(N__27190));
    LocalMux I__3487 (
            .O(N__27199),
            .I(N__27187));
    LocalMux I__3486 (
            .O(N__27196),
            .I(N__27184));
    InMux I__3485 (
            .O(N__27195),
            .I(N__27177));
    InMux I__3484 (
            .O(N__27194),
            .I(N__27177));
    InMux I__3483 (
            .O(N__27193),
            .I(N__27174));
    Span4Mux_v I__3482 (
            .O(N__27190),
            .I(N__27169));
    Span4Mux_v I__3481 (
            .O(N__27187),
            .I(N__27169));
    Span4Mux_h I__3480 (
            .O(N__27184),
            .I(N__27166));
    InMux I__3479 (
            .O(N__27183),
            .I(N__27161));
    InMux I__3478 (
            .O(N__27182),
            .I(N__27161));
    LocalMux I__3477 (
            .O(N__27177),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ));
    LocalMux I__3476 (
            .O(N__27174),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ));
    Odrv4 I__3475 (
            .O(N__27169),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ));
    Odrv4 I__3474 (
            .O(N__27166),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ));
    LocalMux I__3473 (
            .O(N__27161),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ));
    CascadeMux I__3472 (
            .O(N__27150),
            .I(N__27128));
    InMux I__3471 (
            .O(N__27149),
            .I(N__27125));
    InMux I__3470 (
            .O(N__27148),
            .I(N__27114));
    InMux I__3469 (
            .O(N__27147),
            .I(N__27114));
    InMux I__3468 (
            .O(N__27146),
            .I(N__27114));
    InMux I__3467 (
            .O(N__27145),
            .I(N__27114));
    InMux I__3466 (
            .O(N__27144),
            .I(N__27114));
    InMux I__3465 (
            .O(N__27143),
            .I(N__27111));
    InMux I__3464 (
            .O(N__27142),
            .I(N__27108));
    InMux I__3463 (
            .O(N__27141),
            .I(N__27098));
    InMux I__3462 (
            .O(N__27140),
            .I(N__27098));
    InMux I__3461 (
            .O(N__27139),
            .I(N__27098));
    InMux I__3460 (
            .O(N__27138),
            .I(N__27098));
    InMux I__3459 (
            .O(N__27137),
            .I(N__27083));
    InMux I__3458 (
            .O(N__27136),
            .I(N__27083));
    InMux I__3457 (
            .O(N__27135),
            .I(N__27083));
    InMux I__3456 (
            .O(N__27134),
            .I(N__27083));
    InMux I__3455 (
            .O(N__27133),
            .I(N__27083));
    InMux I__3454 (
            .O(N__27132),
            .I(N__27083));
    InMux I__3453 (
            .O(N__27131),
            .I(N__27083));
    InMux I__3452 (
            .O(N__27128),
            .I(N__27080));
    LocalMux I__3451 (
            .O(N__27125),
            .I(N__27073));
    LocalMux I__3450 (
            .O(N__27114),
            .I(N__27073));
    LocalMux I__3449 (
            .O(N__27111),
            .I(N__27073));
    LocalMux I__3448 (
            .O(N__27108),
            .I(N__27070));
    InMux I__3447 (
            .O(N__27107),
            .I(N__27065));
    LocalMux I__3446 (
            .O(N__27098),
            .I(N__27060));
    LocalMux I__3445 (
            .O(N__27083),
            .I(N__27060));
    LocalMux I__3444 (
            .O(N__27080),
            .I(N__27055));
    Span4Mux_h I__3443 (
            .O(N__27073),
            .I(N__27055));
    Span4Mux_h I__3442 (
            .O(N__27070),
            .I(N__27052));
    InMux I__3441 (
            .O(N__27069),
            .I(N__27047));
    InMux I__3440 (
            .O(N__27068),
            .I(N__27047));
    LocalMux I__3439 (
            .O(N__27065),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ));
    Odrv12 I__3438 (
            .O(N__27060),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ));
    Odrv4 I__3437 (
            .O(N__27055),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ));
    Odrv4 I__3436 (
            .O(N__27052),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ));
    LocalMux I__3435 (
            .O(N__27047),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ));
    CascadeMux I__3434 (
            .O(N__27036),
            .I(N__27032));
    InMux I__3433 (
            .O(N__27035),
            .I(N__27027));
    InMux I__3432 (
            .O(N__27032),
            .I(N__27027));
    LocalMux I__3431 (
            .O(N__27027),
            .I(N__27024));
    Odrv12 I__3430 (
            .O(N__27024),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_391 ));
    InMux I__3429 (
            .O(N__27021),
            .I(N__27018));
    LocalMux I__3428 (
            .O(N__27018),
            .I(N__27015));
    Odrv4 I__3427 (
            .O(N__27015),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_8 ));
    InMux I__3426 (
            .O(N__27012),
            .I(N__27009));
    LocalMux I__3425 (
            .O(N__27009),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_11 ));
    InMux I__3424 (
            .O(N__27006),
            .I(N__27003));
    LocalMux I__3423 (
            .O(N__27003),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_12 ));
    InMux I__3422 (
            .O(N__27000),
            .I(N__26991));
    InMux I__3421 (
            .O(N__26999),
            .I(N__26983));
    InMux I__3420 (
            .O(N__26998),
            .I(N__26983));
    InMux I__3419 (
            .O(N__26997),
            .I(N__26983));
    InMux I__3418 (
            .O(N__26996),
            .I(N__26977));
    InMux I__3417 (
            .O(N__26995),
            .I(N__26977));
    InMux I__3416 (
            .O(N__26994),
            .I(N__26973));
    LocalMux I__3415 (
            .O(N__26991),
            .I(N__26970));
    InMux I__3414 (
            .O(N__26990),
            .I(N__26967));
    LocalMux I__3413 (
            .O(N__26983),
            .I(N__26964));
    InMux I__3412 (
            .O(N__26982),
            .I(N__26961));
    LocalMux I__3411 (
            .O(N__26977),
            .I(N__26958));
    InMux I__3410 (
            .O(N__26976),
            .I(N__26955));
    LocalMux I__3409 (
            .O(N__26973),
            .I(N__26948));
    Span4Mux_v I__3408 (
            .O(N__26970),
            .I(N__26948));
    LocalMux I__3407 (
            .O(N__26967),
            .I(N__26948));
    Odrv4 I__3406 (
            .O(N__26964),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ));
    LocalMux I__3405 (
            .O(N__26961),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ));
    Odrv12 I__3404 (
            .O(N__26958),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ));
    LocalMux I__3403 (
            .O(N__26955),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ));
    Odrv4 I__3402 (
            .O(N__26948),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ));
    InMux I__3401 (
            .O(N__26937),
            .I(N__26934));
    LocalMux I__3400 (
            .O(N__26934),
            .I(N__26928));
    InMux I__3399 (
            .O(N__26933),
            .I(N__26925));
    InMux I__3398 (
            .O(N__26932),
            .I(N__26920));
    InMux I__3397 (
            .O(N__26931),
            .I(N__26917));
    Span4Mux_h I__3396 (
            .O(N__26928),
            .I(N__26914));
    LocalMux I__3395 (
            .O(N__26925),
            .I(N__26911));
    InMux I__3394 (
            .O(N__26924),
            .I(N__26906));
    InMux I__3393 (
            .O(N__26923),
            .I(N__26906));
    LocalMux I__3392 (
            .O(N__26920),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ));
    LocalMux I__3391 (
            .O(N__26917),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ));
    Odrv4 I__3390 (
            .O(N__26914),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ));
    Odrv12 I__3389 (
            .O(N__26911),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ));
    LocalMux I__3388 (
            .O(N__26906),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ));
    CascadeMux I__3387 (
            .O(N__26895),
            .I(N__26890));
    InMux I__3386 (
            .O(N__26894),
            .I(N__26883));
    InMux I__3385 (
            .O(N__26893),
            .I(N__26883));
    InMux I__3384 (
            .O(N__26890),
            .I(N__26878));
    InMux I__3383 (
            .O(N__26889),
            .I(N__26878));
    InMux I__3382 (
            .O(N__26888),
            .I(N__26875));
    LocalMux I__3381 (
            .O(N__26883),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i ));
    LocalMux I__3380 (
            .O(N__26878),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i ));
    LocalMux I__3379 (
            .O(N__26875),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i ));
    InMux I__3378 (
            .O(N__26868),
            .I(N__26865));
    LocalMux I__3377 (
            .O(N__26865),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_12 ));
    InMux I__3376 (
            .O(N__26862),
            .I(N__26859));
    LocalMux I__3375 (
            .O(N__26859),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_13 ));
    InMux I__3374 (
            .O(N__26856),
            .I(N__26853));
    LocalMux I__3373 (
            .O(N__26853),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_14 ));
    InMux I__3372 (
            .O(N__26850),
            .I(N__26847));
    LocalMux I__3371 (
            .O(N__26847),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_15 ));
    InMux I__3370 (
            .O(N__26844),
            .I(N__26841));
    LocalMux I__3369 (
            .O(N__26841),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_14 ));
    InMux I__3368 (
            .O(N__26838),
            .I(N__26835));
    LocalMux I__3367 (
            .O(N__26835),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_21 ));
    InMux I__3366 (
            .O(N__26832),
            .I(N__26829));
    LocalMux I__3365 (
            .O(N__26829),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_20 ));
    InMux I__3364 (
            .O(N__26826),
            .I(N__26823));
    LocalMux I__3363 (
            .O(N__26823),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_9 ));
    InMux I__3362 (
            .O(N__26820),
            .I(N__26817));
    LocalMux I__3361 (
            .O(N__26817),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_8 ));
    InMux I__3360 (
            .O(N__26814),
            .I(N__26811));
    LocalMux I__3359 (
            .O(N__26811),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_10 ));
    InMux I__3358 (
            .O(N__26808),
            .I(N__26805));
    LocalMux I__3357 (
            .O(N__26805),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_22 ));
    InMux I__3356 (
            .O(N__26802),
            .I(N__26799));
    LocalMux I__3355 (
            .O(N__26799),
            .I(N__26796));
    Span4Mux_v I__3354 (
            .O(N__26796),
            .I(N__26793));
    Odrv4 I__3353 (
            .O(N__26793),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.dout_op ));
    InMux I__3352 (
            .O(N__26790),
            .I(N__26787));
    LocalMux I__3351 (
            .O(N__26787),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_18 ));
    InMux I__3350 (
            .O(N__26784),
            .I(N__26781));
    LocalMux I__3349 (
            .O(N__26781),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_19 ));
    InMux I__3348 (
            .O(N__26778),
            .I(N__26775));
    LocalMux I__3347 (
            .O(N__26775),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_6 ));
    InMux I__3346 (
            .O(N__26772),
            .I(N__26769));
    LocalMux I__3345 (
            .O(N__26769),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_17 ));
    InMux I__3344 (
            .O(N__26766),
            .I(N__26763));
    LocalMux I__3343 (
            .O(N__26763),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_16 ));
    InMux I__3342 (
            .O(N__26760),
            .I(N__26757));
    LocalMux I__3341 (
            .O(N__26757),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_15 ));
    InMux I__3340 (
            .O(N__26754),
            .I(N__26751));
    LocalMux I__3339 (
            .O(N__26751),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_13 ));
    CascadeMux I__3338 (
            .O(N__26748),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_5_cascade_ ));
    InMux I__3337 (
            .O(N__26745),
            .I(N__26742));
    LocalMux I__3336 (
            .O(N__26742),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_5 ));
    InMux I__3335 (
            .O(N__26739),
            .I(N__26736));
    LocalMux I__3334 (
            .O(N__26736),
            .I(N__26733));
    Span4Mux_h I__3333 (
            .O(N__26733),
            .I(N__26730));
    Sp12to4 I__3332 (
            .O(N__26730),
            .I(N__26727));
    Odrv12 I__3331 (
            .O(N__26727),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_5));
    CascadeMux I__3330 (
            .O(N__26724),
            .I(N__26721));
    InMux I__3329 (
            .O(N__26721),
            .I(N__26718));
    LocalMux I__3328 (
            .O(N__26718),
            .I(N__26715));
    Span4Mux_v I__3327 (
            .O(N__26715),
            .I(N__26712));
    Span4Mux_v I__3326 (
            .O(N__26712),
            .I(N__26709));
    Odrv4 I__3325 (
            .O(N__26709),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_5));
    CascadeMux I__3324 (
            .O(N__26706),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_5_cascade_ ));
    InMux I__3323 (
            .O(N__26703),
            .I(N__26700));
    LocalMux I__3322 (
            .O(N__26700),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_5 ));
    InMux I__3321 (
            .O(N__26697),
            .I(N__26694));
    LocalMux I__3320 (
            .O(N__26694),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6 ));
    InMux I__3319 (
            .O(N__26691),
            .I(N__26688));
    LocalMux I__3318 (
            .O(N__26688),
            .I(N__26685));
    Odrv12 I__3317 (
            .O(N__26685),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_6 ));
    InMux I__3316 (
            .O(N__26682),
            .I(N__26679));
    LocalMux I__3315 (
            .O(N__26679),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_5 ));
    CascadeMux I__3314 (
            .O(N__26676),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283_cascade_ ));
    InMux I__3313 (
            .O(N__26673),
            .I(N__26669));
    InMux I__3312 (
            .O(N__26672),
            .I(N__26666));
    LocalMux I__3311 (
            .O(N__26669),
            .I(N__26662));
    LocalMux I__3310 (
            .O(N__26666),
            .I(N__26659));
    InMux I__3309 (
            .O(N__26665),
            .I(N__26656));
    Span4Mux_s3_v I__3308 (
            .O(N__26662),
            .I(N__26652));
    Span4Mux_v I__3307 (
            .O(N__26659),
            .I(N__26647));
    LocalMux I__3306 (
            .O(N__26656),
            .I(N__26647));
    InMux I__3305 (
            .O(N__26655),
            .I(N__26644));
    Odrv4 I__3304 (
            .O(N__26652),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0 ));
    Odrv4 I__3303 (
            .O(N__26647),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0 ));
    LocalMux I__3302 (
            .O(N__26644),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0 ));
    CEMux I__3301 (
            .O(N__26637),
            .I(N__26633));
    CEMux I__3300 (
            .O(N__26636),
            .I(N__26630));
    LocalMux I__3299 (
            .O(N__26633),
            .I(N__26627));
    LocalMux I__3298 (
            .O(N__26630),
            .I(N__26624));
    Span4Mux_h I__3297 (
            .O(N__26627),
            .I(N__26621));
    Span4Mux_h I__3296 (
            .O(N__26624),
            .I(N__26618));
    Odrv4 I__3295 (
            .O(N__26621),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0 ));
    Odrv4 I__3294 (
            .O(N__26618),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0 ));
    InMux I__3293 (
            .O(N__26613),
            .I(N__26610));
    LocalMux I__3292 (
            .O(N__26610),
            .I(N__26607));
    Span12Mux_v I__3291 (
            .O(N__26607),
            .I(N__26604));
    Odrv12 I__3290 (
            .O(N__26604),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_1));
    CascadeMux I__3289 (
            .O(N__26601),
            .I(N__26598));
    InMux I__3288 (
            .O(N__26598),
            .I(N__26595));
    LocalMux I__3287 (
            .O(N__26595),
            .I(N__26592));
    Span4Mux_v I__3286 (
            .O(N__26592),
            .I(N__26589));
    Odrv4 I__3285 (
            .O(N__26589),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_1));
    CascadeMux I__3284 (
            .O(N__26586),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_1_cascade_ ));
    InMux I__3283 (
            .O(N__26583),
            .I(N__26580));
    LocalMux I__3282 (
            .O(N__26580),
            .I(N__26577));
    Span4Mux_h I__3281 (
            .O(N__26577),
            .I(N__26574));
    Odrv4 I__3280 (
            .O(N__26574),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_1));
    CascadeMux I__3279 (
            .O(N__26571),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_1_cascade_ ));
    CascadeMux I__3278 (
            .O(N__26568),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_1_cascade_ ));
    InMux I__3277 (
            .O(N__26565),
            .I(N__26562));
    LocalMux I__3276 (
            .O(N__26562),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_1 ));
    InMux I__3275 (
            .O(N__26559),
            .I(N__26556));
    LocalMux I__3274 (
            .O(N__26556),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5 ));
    InMux I__3273 (
            .O(N__26553),
            .I(N__26549));
    InMux I__3272 (
            .O(N__26552),
            .I(N__26545));
    LocalMux I__3271 (
            .O(N__26549),
            .I(N__26542));
    InMux I__3270 (
            .O(N__26548),
            .I(N__26539));
    LocalMux I__3269 (
            .O(N__26545),
            .I(N__26535));
    Span4Mux_v I__3268 (
            .O(N__26542),
            .I(N__26530));
    LocalMux I__3267 (
            .O(N__26539),
            .I(N__26530));
    InMux I__3266 (
            .O(N__26538),
            .I(N__26527));
    Span4Mux_h I__3265 (
            .O(N__26535),
            .I(N__26524));
    Span4Mux_v I__3264 (
            .O(N__26530),
            .I(N__26519));
    LocalMux I__3263 (
            .O(N__26527),
            .I(N__26519));
    Odrv4 I__3262 (
            .O(N__26524),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0 ));
    Odrv4 I__3261 (
            .O(N__26519),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0 ));
    InMux I__3260 (
            .O(N__26514),
            .I(N__26511));
    LocalMux I__3259 (
            .O(N__26511),
            .I(N__26506));
    InMux I__3258 (
            .O(N__26510),
            .I(N__26503));
    InMux I__3257 (
            .O(N__26509),
            .I(N__26499));
    Span4Mux_h I__3256 (
            .O(N__26506),
            .I(N__26496));
    LocalMux I__3255 (
            .O(N__26503),
            .I(N__26493));
    InMux I__3254 (
            .O(N__26502),
            .I(N__26490));
    LocalMux I__3253 (
            .O(N__26499),
            .I(N__26487));
    Span4Mux_v I__3252 (
            .O(N__26496),
            .I(N__26482));
    Span4Mux_h I__3251 (
            .O(N__26493),
            .I(N__26482));
    LocalMux I__3250 (
            .O(N__26490),
            .I(N__26479));
    Span4Mux_h I__3249 (
            .O(N__26487),
            .I(N__26472));
    Span4Mux_v I__3248 (
            .O(N__26482),
            .I(N__26472));
    Span4Mux_h I__3247 (
            .O(N__26479),
            .I(N__26472));
    Odrv4 I__3246 (
            .O(N__26472),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_455_0 ));
    InMux I__3245 (
            .O(N__26469),
            .I(N__26466));
    LocalMux I__3244 (
            .O(N__26466),
            .I(N__26461));
    InMux I__3243 (
            .O(N__26465),
            .I(N__26458));
    InMux I__3242 (
            .O(N__26464),
            .I(N__26454));
    Span4Mux_h I__3241 (
            .O(N__26461),
            .I(N__26451));
    LocalMux I__3240 (
            .O(N__26458),
            .I(N__26448));
    InMux I__3239 (
            .O(N__26457),
            .I(N__26445));
    LocalMux I__3238 (
            .O(N__26454),
            .I(N__26442));
    Span4Mux_v I__3237 (
            .O(N__26451),
            .I(N__26437));
    Span4Mux_h I__3236 (
            .O(N__26448),
            .I(N__26437));
    LocalMux I__3235 (
            .O(N__26445),
            .I(N__26434));
    Span4Mux_h I__3234 (
            .O(N__26442),
            .I(N__26427));
    Span4Mux_v I__3233 (
            .O(N__26437),
            .I(N__26427));
    Span4Mux_h I__3232 (
            .O(N__26434),
            .I(N__26427));
    Odrv4 I__3231 (
            .O(N__26427),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_454_0 ));
    InMux I__3230 (
            .O(N__26424),
            .I(N__26421));
    LocalMux I__3229 (
            .O(N__26421),
            .I(N__26416));
    InMux I__3228 (
            .O(N__26420),
            .I(N__26413));
    InMux I__3227 (
            .O(N__26419),
            .I(N__26409));
    Span4Mux_v I__3226 (
            .O(N__26416),
            .I(N__26404));
    LocalMux I__3225 (
            .O(N__26413),
            .I(N__26404));
    InMux I__3224 (
            .O(N__26412),
            .I(N__26401));
    LocalMux I__3223 (
            .O(N__26409),
            .I(N__26398));
    Span4Mux_v I__3222 (
            .O(N__26404),
            .I(N__26393));
    LocalMux I__3221 (
            .O(N__26401),
            .I(N__26393));
    Span4Mux_v I__3220 (
            .O(N__26398),
            .I(N__26388));
    Span4Mux_v I__3219 (
            .O(N__26393),
            .I(N__26388));
    Odrv4 I__3218 (
            .O(N__26388),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_453_0 ));
    InMux I__3217 (
            .O(N__26385),
            .I(N__26381));
    InMux I__3216 (
            .O(N__26384),
            .I(N__26377));
    LocalMux I__3215 (
            .O(N__26381),
            .I(N__26373));
    InMux I__3214 (
            .O(N__26380),
            .I(N__26370));
    LocalMux I__3213 (
            .O(N__26377),
            .I(N__26367));
    InMux I__3212 (
            .O(N__26376),
            .I(N__26364));
    Span4Mux_h I__3211 (
            .O(N__26373),
            .I(N__26361));
    LocalMux I__3210 (
            .O(N__26370),
            .I(N__26358));
    Span4Mux_h I__3209 (
            .O(N__26367),
            .I(N__26355));
    LocalMux I__3208 (
            .O(N__26364),
            .I(N__26352));
    Span4Mux_v I__3207 (
            .O(N__26361),
            .I(N__26343));
    Span4Mux_h I__3206 (
            .O(N__26358),
            .I(N__26343));
    Span4Mux_v I__3205 (
            .O(N__26355),
            .I(N__26343));
    Span4Mux_h I__3204 (
            .O(N__26352),
            .I(N__26343));
    Odrv4 I__3203 (
            .O(N__26343),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_463_0 ));
    CascadeMux I__3202 (
            .O(N__26340),
            .I(N__26321));
    CascadeMux I__3201 (
            .O(N__26339),
            .I(N__26317));
    CascadeMux I__3200 (
            .O(N__26338),
            .I(N__26313));
    InMux I__3199 (
            .O(N__26337),
            .I(N__26307));
    InMux I__3198 (
            .O(N__26336),
            .I(N__26307));
    InMux I__3197 (
            .O(N__26335),
            .I(N__26302));
    InMux I__3196 (
            .O(N__26334),
            .I(N__26302));
    InMux I__3195 (
            .O(N__26333),
            .I(N__26297));
    InMux I__3194 (
            .O(N__26332),
            .I(N__26297));
    CascadeMux I__3193 (
            .O(N__26331),
            .I(N__26293));
    CascadeMux I__3192 (
            .O(N__26330),
            .I(N__26289));
    CascadeMux I__3191 (
            .O(N__26329),
            .I(N__26285));
    CascadeMux I__3190 (
            .O(N__26328),
            .I(N__26281));
    CascadeMux I__3189 (
            .O(N__26327),
            .I(N__26278));
    CascadeMux I__3188 (
            .O(N__26326),
            .I(N__26273));
    CascadeMux I__3187 (
            .O(N__26325),
            .I(N__26268));
    CascadeMux I__3186 (
            .O(N__26324),
            .I(N__26265));
    InMux I__3185 (
            .O(N__26321),
            .I(N__26258));
    InMux I__3184 (
            .O(N__26320),
            .I(N__26258));
    InMux I__3183 (
            .O(N__26317),
            .I(N__26249));
    InMux I__3182 (
            .O(N__26316),
            .I(N__26249));
    InMux I__3181 (
            .O(N__26313),
            .I(N__26249));
    InMux I__3180 (
            .O(N__26312),
            .I(N__26249));
    LocalMux I__3179 (
            .O(N__26307),
            .I(N__26246));
    LocalMux I__3178 (
            .O(N__26302),
            .I(N__26241));
    LocalMux I__3177 (
            .O(N__26297),
            .I(N__26241));
    InMux I__3176 (
            .O(N__26296),
            .I(N__26230));
    InMux I__3175 (
            .O(N__26293),
            .I(N__26230));
    InMux I__3174 (
            .O(N__26292),
            .I(N__26230));
    InMux I__3173 (
            .O(N__26289),
            .I(N__26230));
    InMux I__3172 (
            .O(N__26288),
            .I(N__26230));
    InMux I__3171 (
            .O(N__26285),
            .I(N__26213));
    InMux I__3170 (
            .O(N__26284),
            .I(N__26213));
    InMux I__3169 (
            .O(N__26281),
            .I(N__26213));
    InMux I__3168 (
            .O(N__26278),
            .I(N__26213));
    InMux I__3167 (
            .O(N__26277),
            .I(N__26213));
    InMux I__3166 (
            .O(N__26276),
            .I(N__26213));
    InMux I__3165 (
            .O(N__26273),
            .I(N__26213));
    InMux I__3164 (
            .O(N__26272),
            .I(N__26213));
    InMux I__3163 (
            .O(N__26271),
            .I(N__26202));
    InMux I__3162 (
            .O(N__26268),
            .I(N__26202));
    InMux I__3161 (
            .O(N__26265),
            .I(N__26202));
    InMux I__3160 (
            .O(N__26264),
            .I(N__26202));
    InMux I__3159 (
            .O(N__26263),
            .I(N__26202));
    LocalMux I__3158 (
            .O(N__26258),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    LocalMux I__3157 (
            .O(N__26249),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    Odrv4 I__3156 (
            .O(N__26246),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    Odrv4 I__3155 (
            .O(N__26241),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    LocalMux I__3154 (
            .O(N__26230),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    LocalMux I__3153 (
            .O(N__26213),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    LocalMux I__3152 (
            .O(N__26202),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ));
    InMux I__3151 (
            .O(N__26187),
            .I(N__26183));
    InMux I__3150 (
            .O(N__26186),
            .I(N__26179));
    LocalMux I__3149 (
            .O(N__26183),
            .I(N__26176));
    InMux I__3148 (
            .O(N__26182),
            .I(N__26173));
    LocalMux I__3147 (
            .O(N__26179),
            .I(N__26170));
    Span4Mux_h I__3146 (
            .O(N__26176),
            .I(N__26166));
    LocalMux I__3145 (
            .O(N__26173),
            .I(N__26163));
    Span4Mux_h I__3144 (
            .O(N__26170),
            .I(N__26160));
    InMux I__3143 (
            .O(N__26169),
            .I(N__26157));
    Span4Mux_v I__3142 (
            .O(N__26166),
            .I(N__26152));
    Span4Mux_h I__3141 (
            .O(N__26163),
            .I(N__26152));
    Span4Mux_v I__3140 (
            .O(N__26160),
            .I(N__26147));
    LocalMux I__3139 (
            .O(N__26157),
            .I(N__26147));
    Odrv4 I__3138 (
            .O(N__26152),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0 ));
    Odrv4 I__3137 (
            .O(N__26147),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0 ));
    InMux I__3136 (
            .O(N__26142),
            .I(N__26139));
    LocalMux I__3135 (
            .O(N__26139),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_21 ));
    InMux I__3134 (
            .O(N__26136),
            .I(N__26133));
    LocalMux I__3133 (
            .O(N__26133),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_20 ));
    InMux I__3132 (
            .O(N__26130),
            .I(N__26127));
    LocalMux I__3131 (
            .O(N__26127),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_22 ));
    InMux I__3130 (
            .O(N__26124),
            .I(N__26121));
    LocalMux I__3129 (
            .O(N__26121),
            .I(N__26118));
    Odrv12 I__3128 (
            .O(N__26118),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_op ));
    InMux I__3127 (
            .O(N__26115),
            .I(N__26111));
    InMux I__3126 (
            .O(N__26114),
            .I(N__26108));
    LocalMux I__3125 (
            .O(N__26111),
            .I(N__26105));
    LocalMux I__3124 (
            .O(N__26108),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0 ));
    Odrv4 I__3123 (
            .O(N__26105),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0 ));
    InMux I__3122 (
            .O(N__26100),
            .I(bfn_9_22_0_));
    InMux I__3121 (
            .O(N__26097),
            .I(N__26093));
    InMux I__3120 (
            .O(N__26096),
            .I(N__26090));
    LocalMux I__3119 (
            .O(N__26093),
            .I(N__26087));
    LocalMux I__3118 (
            .O(N__26090),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1 ));
    Odrv12 I__3117 (
            .O(N__26087),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1 ));
    InMux I__3116 (
            .O(N__26082),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0 ));
    InMux I__3115 (
            .O(N__26079),
            .I(N__26075));
    InMux I__3114 (
            .O(N__26078),
            .I(N__26072));
    LocalMux I__3113 (
            .O(N__26075),
            .I(N__26069));
    LocalMux I__3112 (
            .O(N__26072),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2 ));
    Odrv4 I__3111 (
            .O(N__26069),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2 ));
    InMux I__3110 (
            .O(N__26064),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1 ));
    InMux I__3109 (
            .O(N__26061),
            .I(N__26058));
    LocalMux I__3108 (
            .O(N__26058),
            .I(N__26054));
    InMux I__3107 (
            .O(N__26057),
            .I(N__26051));
    Span4Mux_h I__3106 (
            .O(N__26054),
            .I(N__26048));
    LocalMux I__3105 (
            .O(N__26051),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3 ));
    Odrv4 I__3104 (
            .O(N__26048),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3 ));
    InMux I__3103 (
            .O(N__26043),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2 ));
    InMux I__3102 (
            .O(N__26040),
            .I(N__26029));
    InMux I__3101 (
            .O(N__26039),
            .I(N__26029));
    InMux I__3100 (
            .O(N__26038),
            .I(N__26029));
    InMux I__3099 (
            .O(N__26037),
            .I(N__26024));
    InMux I__3098 (
            .O(N__26036),
            .I(N__26024));
    LocalMux I__3097 (
            .O(N__26029),
            .I(N__26019));
    LocalMux I__3096 (
            .O(N__26024),
            .I(N__26019));
    Odrv4 I__3095 (
            .O(N__26019),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_391_i ));
    InMux I__3094 (
            .O(N__26016),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_3 ));
    InMux I__3093 (
            .O(N__26013),
            .I(N__26010));
    LocalMux I__3092 (
            .O(N__26010),
            .I(N__26006));
    InMux I__3091 (
            .O(N__26009),
            .I(N__26003));
    Span4Mux_h I__3090 (
            .O(N__26006),
            .I(N__26000));
    LocalMux I__3089 (
            .O(N__26003),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4 ));
    Odrv4 I__3088 (
            .O(N__26000),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4 ));
    InMux I__3087 (
            .O(N__25995),
            .I(N__25992));
    LocalMux I__3086 (
            .O(N__25992),
            .I(N__25987));
    InMux I__3085 (
            .O(N__25991),
            .I(N__25984));
    InMux I__3084 (
            .O(N__25990),
            .I(N__25981));
    Span4Mux_h I__3083 (
            .O(N__25987),
            .I(N__25978));
    LocalMux I__3082 (
            .O(N__25984),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1 ));
    LocalMux I__3081 (
            .O(N__25981),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1 ));
    Odrv4 I__3080 (
            .O(N__25978),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1 ));
    InMux I__3079 (
            .O(N__25971),
            .I(N__25968));
    LocalMux I__3078 (
            .O(N__25968),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_CO ));
    InMux I__3077 (
            .O(N__25965),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0 ));
    InMux I__3076 (
            .O(N__25962),
            .I(N__25959));
    LocalMux I__3075 (
            .O(N__25959),
            .I(N__25954));
    InMux I__3074 (
            .O(N__25958),
            .I(N__25951));
    InMux I__3073 (
            .O(N__25957),
            .I(N__25948));
    Span4Mux_h I__3072 (
            .O(N__25954),
            .I(N__25945));
    LocalMux I__3071 (
            .O(N__25951),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2 ));
    LocalMux I__3070 (
            .O(N__25948),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2 ));
    Odrv4 I__3069 (
            .O(N__25945),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2 ));
    CascadeMux I__3068 (
            .O(N__25938),
            .I(N__25935));
    InMux I__3067 (
            .O(N__25935),
            .I(N__25932));
    LocalMux I__3066 (
            .O(N__25932),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_CO ));
    InMux I__3065 (
            .O(N__25929),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1 ));
    InMux I__3064 (
            .O(N__25926),
            .I(N__25922));
    CascadeMux I__3063 (
            .O(N__25925),
            .I(N__25919));
    LocalMux I__3062 (
            .O(N__25922),
            .I(N__25915));
    InMux I__3061 (
            .O(N__25919),
            .I(N__25912));
    InMux I__3060 (
            .O(N__25918),
            .I(N__25909));
    Span4Mux_v I__3059 (
            .O(N__25915),
            .I(N__25906));
    LocalMux I__3058 (
            .O(N__25912),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3 ));
    LocalMux I__3057 (
            .O(N__25909),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3 ));
    Odrv4 I__3056 (
            .O(N__25906),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3 ));
    InMux I__3055 (
            .O(N__25899),
            .I(N__25896));
    LocalMux I__3054 (
            .O(N__25896),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_CO ));
    InMux I__3053 (
            .O(N__25893),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2 ));
    InMux I__3052 (
            .O(N__25890),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_3 ));
    CascadeMux I__3051 (
            .O(N__25887),
            .I(N__25884));
    InMux I__3050 (
            .O(N__25884),
            .I(N__25880));
    InMux I__3049 (
            .O(N__25883),
            .I(N__25877));
    LocalMux I__3048 (
            .O(N__25880),
            .I(N__25874));
    LocalMux I__3047 (
            .O(N__25877),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4 ));
    Odrv4 I__3046 (
            .O(N__25874),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4 ));
    InMux I__3045 (
            .O(N__25869),
            .I(N__25866));
    LocalMux I__3044 (
            .O(N__25866),
            .I(N__25863));
    Span4Mux_v I__3043 (
            .O(N__25863),
            .I(N__25860));
    Odrv4 I__3042 (
            .O(N__25860),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_a2_1_0 ));
    InMux I__3041 (
            .O(N__25857),
            .I(N__25854));
    LocalMux I__3040 (
            .O(N__25854),
            .I(N__25851));
    Span4Mux_h I__3039 (
            .O(N__25851),
            .I(N__25848));
    Odrv4 I__3038 (
            .O(N__25848),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_3 ));
    CascadeMux I__3037 (
            .O(N__25845),
            .I(N__25841));
    InMux I__3036 (
            .O(N__25844),
            .I(N__25835));
    InMux I__3035 (
            .O(N__25841),
            .I(N__25832));
    InMux I__3034 (
            .O(N__25840),
            .I(N__25829));
    InMux I__3033 (
            .O(N__25839),
            .I(N__25824));
    InMux I__3032 (
            .O(N__25838),
            .I(N__25824));
    LocalMux I__3031 (
            .O(N__25835),
            .I(N__25821));
    LocalMux I__3030 (
            .O(N__25832),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14 ));
    LocalMux I__3029 (
            .O(N__25829),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14 ));
    LocalMux I__3028 (
            .O(N__25824),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14 ));
    Odrv12 I__3027 (
            .O(N__25821),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14 ));
    CascadeMux I__3026 (
            .O(N__25812),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_cascade_ ));
    InMux I__3025 (
            .O(N__25809),
            .I(N__25805));
    InMux I__3024 (
            .O(N__25808),
            .I(N__25799));
    LocalMux I__3023 (
            .O(N__25805),
            .I(N__25796));
    InMux I__3022 (
            .O(N__25804),
            .I(N__25789));
    InMux I__3021 (
            .O(N__25803),
            .I(N__25789));
    InMux I__3020 (
            .O(N__25802),
            .I(N__25789));
    LocalMux I__3019 (
            .O(N__25799),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6 ));
    Odrv4 I__3018 (
            .O(N__25796),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6 ));
    LocalMux I__3017 (
            .O(N__25789),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6 ));
    CascadeMux I__3016 (
            .O(N__25782),
            .I(N__25775));
    InMux I__3015 (
            .O(N__25781),
            .I(N__25766));
    InMux I__3014 (
            .O(N__25780),
            .I(N__25766));
    InMux I__3013 (
            .O(N__25779),
            .I(N__25766));
    InMux I__3012 (
            .O(N__25778),
            .I(N__25766));
    InMux I__3011 (
            .O(N__25775),
            .I(N__25763));
    LocalMux I__3010 (
            .O(N__25766),
            .I(N__25760));
    LocalMux I__3009 (
            .O(N__25763),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0 ));
    Odrv4 I__3008 (
            .O(N__25760),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0 ));
    InMux I__3007 (
            .O(N__25755),
            .I(N__25752));
    LocalMux I__3006 (
            .O(N__25752),
            .I(N__25748));
    CascadeMux I__3005 (
            .O(N__25751),
            .I(N__25737));
    Span4Mux_v I__3004 (
            .O(N__25748),
            .I(N__25733));
    InMux I__3003 (
            .O(N__25747),
            .I(N__25716));
    InMux I__3002 (
            .O(N__25746),
            .I(N__25716));
    InMux I__3001 (
            .O(N__25745),
            .I(N__25716));
    InMux I__3000 (
            .O(N__25744),
            .I(N__25716));
    InMux I__2999 (
            .O(N__25743),
            .I(N__25716));
    InMux I__2998 (
            .O(N__25742),
            .I(N__25716));
    InMux I__2997 (
            .O(N__25741),
            .I(N__25716));
    InMux I__2996 (
            .O(N__25740),
            .I(N__25716));
    InMux I__2995 (
            .O(N__25737),
            .I(N__25711));
    InMux I__2994 (
            .O(N__25736),
            .I(N__25711));
    Odrv4 I__2993 (
            .O(N__25733),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10 ));
    LocalMux I__2992 (
            .O(N__25716),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10 ));
    LocalMux I__2991 (
            .O(N__25711),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10 ));
    CascadeMux I__2990 (
            .O(N__25704),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.csb_u_i_a2_0_0_cascade_ ));
    CascadeMux I__2989 (
            .O(N__25701),
            .I(N__25698));
    InMux I__2988 (
            .O(N__25698),
            .I(N__25690));
    InMux I__2987 (
            .O(N__25697),
            .I(N__25690));
    CascadeMux I__2986 (
            .O(N__25696),
            .I(N__25687));
    InMux I__2985 (
            .O(N__25695),
            .I(N__25683));
    LocalMux I__2984 (
            .O(N__25690),
            .I(N__25678));
    InMux I__2983 (
            .O(N__25687),
            .I(N__25673));
    InMux I__2982 (
            .O(N__25686),
            .I(N__25673));
    LocalMux I__2981 (
            .O(N__25683),
            .I(N__25670));
    InMux I__2980 (
            .O(N__25682),
            .I(N__25665));
    InMux I__2979 (
            .O(N__25681),
            .I(N__25665));
    Span4Mux_v I__2978 (
            .O(N__25678),
            .I(N__25660));
    LocalMux I__2977 (
            .O(N__25673),
            .I(N__25660));
    Odrv4 I__2976 (
            .O(N__25670),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0 ));
    LocalMux I__2975 (
            .O(N__25665),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0 ));
    Odrv4 I__2974 (
            .O(N__25660),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0 ));
    IoInMux I__2973 (
            .O(N__25653),
            .I(N__25650));
    LocalMux I__2972 (
            .O(N__25650),
            .I(N__25647));
    Span4Mux_s0_h I__2971 (
            .O(N__25647),
            .I(N__25644));
    Sp12to4 I__2970 (
            .O(N__25644),
            .I(N__25641));
    Span12Mux_v I__2969 (
            .O(N__25641),
            .I(N__25638));
    Odrv12 I__2968 (
            .O(N__25638),
            .I(N_1822_0));
    InMux I__2967 (
            .O(N__25635),
            .I(N__25632));
    LocalMux I__2966 (
            .O(N__25632),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.csb_u_i_a2_0 ));
    InMux I__2965 (
            .O(N__25629),
            .I(N__25623));
    InMux I__2964 (
            .O(N__25628),
            .I(N__25618));
    InMux I__2963 (
            .O(N__25627),
            .I(N__25618));
    InMux I__2962 (
            .O(N__25626),
            .I(N__25613));
    LocalMux I__2961 (
            .O(N__25623),
            .I(N__25608));
    LocalMux I__2960 (
            .O(N__25618),
            .I(N__25608));
    InMux I__2959 (
            .O(N__25617),
            .I(N__25605));
    InMux I__2958 (
            .O(N__25616),
            .I(N__25602));
    LocalMux I__2957 (
            .O(N__25613),
            .I(N__25595));
    Span4Mux_v I__2956 (
            .O(N__25608),
            .I(N__25595));
    LocalMux I__2955 (
            .O(N__25605),
            .I(N__25595));
    LocalMux I__2954 (
            .O(N__25602),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0 ));
    Odrv4 I__2953 (
            .O(N__25595),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0 ));
    InMux I__2952 (
            .O(N__25590),
            .I(N__25587));
    LocalMux I__2951 (
            .O(N__25587),
            .I(N__25584));
    Span4Mux_h I__2950 (
            .O(N__25584),
            .I(N__25578));
    InMux I__2949 (
            .O(N__25583),
            .I(N__25574));
    InMux I__2948 (
            .O(N__25582),
            .I(N__25569));
    InMux I__2947 (
            .O(N__25581),
            .I(N__25569));
    Span4Mux_v I__2946 (
            .O(N__25578),
            .I(N__25566));
    InMux I__2945 (
            .O(N__25577),
            .I(N__25563));
    LocalMux I__2944 (
            .O(N__25574),
            .I(N__25560));
    LocalMux I__2943 (
            .O(N__25569),
            .I(N__25557));
    Span4Mux_v I__2942 (
            .O(N__25566),
            .I(N__25554));
    LocalMux I__2941 (
            .O(N__25563),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0 ));
    Odrv4 I__2940 (
            .O(N__25560),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0 ));
    Odrv12 I__2939 (
            .O(N__25557),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0 ));
    Odrv4 I__2938 (
            .O(N__25554),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0 ));
    InMux I__2937 (
            .O(N__25545),
            .I(N__25542));
    LocalMux I__2936 (
            .O(N__25542),
            .I(N__25539));
    Odrv4 I__2935 (
            .O(N__25539),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_CO ));
    InMux I__2934 (
            .O(N__25536),
            .I(N__25531));
    CascadeMux I__2933 (
            .O(N__25535),
            .I(N__25527));
    CascadeMux I__2932 (
            .O(N__25534),
            .I(N__25524));
    LocalMux I__2931 (
            .O(N__25531),
            .I(N__25520));
    InMux I__2930 (
            .O(N__25530),
            .I(N__25517));
    InMux I__2929 (
            .O(N__25527),
            .I(N__25514));
    InMux I__2928 (
            .O(N__25524),
            .I(N__25509));
    InMux I__2927 (
            .O(N__25523),
            .I(N__25509));
    Sp12to4 I__2926 (
            .O(N__25520),
            .I(N__25506));
    LocalMux I__2925 (
            .O(N__25517),
            .I(N__25503));
    LocalMux I__2924 (
            .O(N__25514),
            .I(N__25496));
    LocalMux I__2923 (
            .O(N__25509),
            .I(N__25496));
    Span12Mux_v I__2922 (
            .O(N__25506),
            .I(N__25496));
    Odrv4 I__2921 (
            .O(N__25503),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i ));
    Odrv12 I__2920 (
            .O(N__25496),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i ));
    CascadeMux I__2919 (
            .O(N__25491),
            .I(N__25488));
    InMux I__2918 (
            .O(N__25488),
            .I(N__25484));
    InMux I__2917 (
            .O(N__25487),
            .I(N__25480));
    LocalMux I__2916 (
            .O(N__25484),
            .I(N__25477));
    InMux I__2915 (
            .O(N__25483),
            .I(N__25474));
    LocalMux I__2914 (
            .O(N__25480),
            .I(N__25471));
    Span4Mux_h I__2913 (
            .O(N__25477),
            .I(N__25468));
    LocalMux I__2912 (
            .O(N__25474),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1 ));
    Odrv4 I__2911 (
            .O(N__25471),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1 ));
    Odrv4 I__2910 (
            .O(N__25468),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1 ));
    InMux I__2909 (
            .O(N__25461),
            .I(N__25453));
    InMux I__2908 (
            .O(N__25460),
            .I(N__25453));
    InMux I__2907 (
            .O(N__25459),
            .I(N__25448));
    InMux I__2906 (
            .O(N__25458),
            .I(N__25448));
    LocalMux I__2905 (
            .O(N__25453),
            .I(N__25444));
    LocalMux I__2904 (
            .O(N__25448),
            .I(N__25441));
    InMux I__2903 (
            .O(N__25447),
            .I(N__25437));
    Span4Mux_v I__2902 (
            .O(N__25444),
            .I(N__25432));
    Span4Mux_v I__2901 (
            .O(N__25441),
            .I(N__25432));
    InMux I__2900 (
            .O(N__25440),
            .I(N__25429));
    LocalMux I__2899 (
            .O(N__25437),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0 ));
    Odrv4 I__2898 (
            .O(N__25432),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0 ));
    LocalMux I__2897 (
            .O(N__25429),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0 ));
    IoInMux I__2896 (
            .O(N__25422),
            .I(N__25419));
    LocalMux I__2895 (
            .O(N__25419),
            .I(N__25416));
    IoSpan4Mux I__2894 (
            .O(N__25416),
            .I(N__25413));
    Span4Mux_s3_h I__2893 (
            .O(N__25413),
            .I(N__25410));
    Span4Mux_h I__2892 (
            .O(N__25410),
            .I(N__25407));
    Odrv4 I__2891 (
            .O(N__25407),
            .I(\I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_iZ0 ));
    CascadeMux I__2890 (
            .O(N__25404),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_596_cascade_ ));
    InMux I__2889 (
            .O(N__25401),
            .I(N__25398));
    LocalMux I__2888 (
            .O(N__25398),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_597 ));
    InMux I__2887 (
            .O(N__25395),
            .I(N__25392));
    LocalMux I__2886 (
            .O(N__25392),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_oZ0Z_26 ));
    CascadeMux I__2885 (
            .O(N__25389),
            .I(\cemf_module_64ch_ctrl_inst1.N_1615_cascade_ ));
    CascadeMux I__2884 (
            .O(N__25386),
            .I(N__25382));
    CascadeMux I__2883 (
            .O(N__25385),
            .I(N__25379));
    CascadeBuf I__2882 (
            .O(N__25382),
            .I(N__25376));
    CascadeBuf I__2881 (
            .O(N__25379),
            .I(N__25373));
    CascadeMux I__2880 (
            .O(N__25376),
            .I(N__25370));
    CascadeMux I__2879 (
            .O(N__25373),
            .I(N__25367));
    CascadeBuf I__2878 (
            .O(N__25370),
            .I(N__25364));
    CascadeBuf I__2877 (
            .O(N__25367),
            .I(N__25361));
    CascadeMux I__2876 (
            .O(N__25364),
            .I(N__25358));
    CascadeMux I__2875 (
            .O(N__25361),
            .I(N__25355));
    CascadeBuf I__2874 (
            .O(N__25358),
            .I(N__25352));
    CascadeBuf I__2873 (
            .O(N__25355),
            .I(N__25349));
    CascadeMux I__2872 (
            .O(N__25352),
            .I(N__25346));
    CascadeMux I__2871 (
            .O(N__25349),
            .I(N__25343));
    CascadeBuf I__2870 (
            .O(N__25346),
            .I(N__25340));
    CascadeBuf I__2869 (
            .O(N__25343),
            .I(N__25337));
    CascadeMux I__2868 (
            .O(N__25340),
            .I(N__25334));
    CascadeMux I__2867 (
            .O(N__25337),
            .I(N__25331));
    CascadeBuf I__2866 (
            .O(N__25334),
            .I(N__25328));
    CascadeBuf I__2865 (
            .O(N__25331),
            .I(N__25325));
    CascadeMux I__2864 (
            .O(N__25328),
            .I(N__25322));
    CascadeMux I__2863 (
            .O(N__25325),
            .I(N__25319));
    CascadeBuf I__2862 (
            .O(N__25322),
            .I(N__25316));
    CascadeBuf I__2861 (
            .O(N__25319),
            .I(N__25313));
    CascadeMux I__2860 (
            .O(N__25316),
            .I(N__25310));
    CascadeMux I__2859 (
            .O(N__25313),
            .I(N__25307));
    CascadeBuf I__2858 (
            .O(N__25310),
            .I(N__25304));
    CascadeBuf I__2857 (
            .O(N__25307),
            .I(N__25301));
    CascadeMux I__2856 (
            .O(N__25304),
            .I(N__25298));
    CascadeMux I__2855 (
            .O(N__25301),
            .I(N__25295));
    InMux I__2854 (
            .O(N__25298),
            .I(N__25292));
    InMux I__2853 (
            .O(N__25295),
            .I(N__25289));
    LocalMux I__2852 (
            .O(N__25292),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0 ));
    LocalMux I__2851 (
            .O(N__25289),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0 ));
    CascadeMux I__2850 (
            .O(N__25284),
            .I(N__25280));
    CascadeMux I__2849 (
            .O(N__25283),
            .I(N__25277));
    CascadeBuf I__2848 (
            .O(N__25280),
            .I(N__25274));
    CascadeBuf I__2847 (
            .O(N__25277),
            .I(N__25271));
    CascadeMux I__2846 (
            .O(N__25274),
            .I(N__25268));
    CascadeMux I__2845 (
            .O(N__25271),
            .I(N__25265));
    CascadeBuf I__2844 (
            .O(N__25268),
            .I(N__25262));
    CascadeBuf I__2843 (
            .O(N__25265),
            .I(N__25259));
    CascadeMux I__2842 (
            .O(N__25262),
            .I(N__25256));
    CascadeMux I__2841 (
            .O(N__25259),
            .I(N__25253));
    CascadeBuf I__2840 (
            .O(N__25256),
            .I(N__25250));
    CascadeBuf I__2839 (
            .O(N__25253),
            .I(N__25247));
    CascadeMux I__2838 (
            .O(N__25250),
            .I(N__25244));
    CascadeMux I__2837 (
            .O(N__25247),
            .I(N__25241));
    CascadeBuf I__2836 (
            .O(N__25244),
            .I(N__25238));
    CascadeBuf I__2835 (
            .O(N__25241),
            .I(N__25235));
    CascadeMux I__2834 (
            .O(N__25238),
            .I(N__25232));
    CascadeMux I__2833 (
            .O(N__25235),
            .I(N__25229));
    CascadeBuf I__2832 (
            .O(N__25232),
            .I(N__25226));
    CascadeBuf I__2831 (
            .O(N__25229),
            .I(N__25223));
    CascadeMux I__2830 (
            .O(N__25226),
            .I(N__25220));
    CascadeMux I__2829 (
            .O(N__25223),
            .I(N__25217));
    CascadeBuf I__2828 (
            .O(N__25220),
            .I(N__25214));
    CascadeBuf I__2827 (
            .O(N__25217),
            .I(N__25211));
    CascadeMux I__2826 (
            .O(N__25214),
            .I(N__25208));
    CascadeMux I__2825 (
            .O(N__25211),
            .I(N__25205));
    CascadeBuf I__2824 (
            .O(N__25208),
            .I(N__25202));
    CascadeBuf I__2823 (
            .O(N__25205),
            .I(N__25199));
    CascadeMux I__2822 (
            .O(N__25202),
            .I(N__25196));
    CascadeMux I__2821 (
            .O(N__25199),
            .I(N__25193));
    InMux I__2820 (
            .O(N__25196),
            .I(N__25190));
    InMux I__2819 (
            .O(N__25193),
            .I(N__25187));
    LocalMux I__2818 (
            .O(N__25190),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0 ));
    LocalMux I__2817 (
            .O(N__25187),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0 ));
    CascadeMux I__2816 (
            .O(N__25182),
            .I(N__25178));
    CascadeMux I__2815 (
            .O(N__25181),
            .I(N__25175));
    CascadeBuf I__2814 (
            .O(N__25178),
            .I(N__25172));
    CascadeBuf I__2813 (
            .O(N__25175),
            .I(N__25169));
    CascadeMux I__2812 (
            .O(N__25172),
            .I(N__25166));
    CascadeMux I__2811 (
            .O(N__25169),
            .I(N__25163));
    CascadeBuf I__2810 (
            .O(N__25166),
            .I(N__25160));
    CascadeBuf I__2809 (
            .O(N__25163),
            .I(N__25157));
    CascadeMux I__2808 (
            .O(N__25160),
            .I(N__25154));
    CascadeMux I__2807 (
            .O(N__25157),
            .I(N__25151));
    CascadeBuf I__2806 (
            .O(N__25154),
            .I(N__25148));
    CascadeBuf I__2805 (
            .O(N__25151),
            .I(N__25145));
    CascadeMux I__2804 (
            .O(N__25148),
            .I(N__25142));
    CascadeMux I__2803 (
            .O(N__25145),
            .I(N__25139));
    CascadeBuf I__2802 (
            .O(N__25142),
            .I(N__25136));
    CascadeBuf I__2801 (
            .O(N__25139),
            .I(N__25133));
    CascadeMux I__2800 (
            .O(N__25136),
            .I(N__25130));
    CascadeMux I__2799 (
            .O(N__25133),
            .I(N__25127));
    CascadeBuf I__2798 (
            .O(N__25130),
            .I(N__25124));
    CascadeBuf I__2797 (
            .O(N__25127),
            .I(N__25121));
    CascadeMux I__2796 (
            .O(N__25124),
            .I(N__25118));
    CascadeMux I__2795 (
            .O(N__25121),
            .I(N__25115));
    CascadeBuf I__2794 (
            .O(N__25118),
            .I(N__25112));
    CascadeBuf I__2793 (
            .O(N__25115),
            .I(N__25109));
    CascadeMux I__2792 (
            .O(N__25112),
            .I(N__25106));
    CascadeMux I__2791 (
            .O(N__25109),
            .I(N__25103));
    CascadeBuf I__2790 (
            .O(N__25106),
            .I(N__25100));
    CascadeBuf I__2789 (
            .O(N__25103),
            .I(N__25097));
    CascadeMux I__2788 (
            .O(N__25100),
            .I(N__25094));
    CascadeMux I__2787 (
            .O(N__25097),
            .I(N__25091));
    InMux I__2786 (
            .O(N__25094),
            .I(N__25088));
    InMux I__2785 (
            .O(N__25091),
            .I(N__25085));
    LocalMux I__2784 (
            .O(N__25088),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3 ));
    LocalMux I__2783 (
            .O(N__25085),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3 ));
    InMux I__2782 (
            .O(N__25080),
            .I(N__25077));
    LocalMux I__2781 (
            .O(N__25077),
            .I(N__25071));
    InMux I__2780 (
            .O(N__25076),
            .I(N__25064));
    InMux I__2779 (
            .O(N__25075),
            .I(N__25064));
    InMux I__2778 (
            .O(N__25074),
            .I(N__25064));
    Odrv12 I__2777 (
            .O(N__25071),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9 ));
    LocalMux I__2776 (
            .O(N__25064),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9 ));
    InMux I__2775 (
            .O(N__25059),
            .I(N__25056));
    LocalMux I__2774 (
            .O(N__25056),
            .I(N__25053));
    Odrv4 I__2773 (
            .O(N__25053),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_6));
    CascadeMux I__2772 (
            .O(N__25050),
            .I(N__25047));
    InMux I__2771 (
            .O(N__25047),
            .I(N__25044));
    LocalMux I__2770 (
            .O(N__25044),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_6 ));
    InMux I__2769 (
            .O(N__25041),
            .I(N__25038));
    LocalMux I__2768 (
            .O(N__25038),
            .I(N__25035));
    Odrv4 I__2767 (
            .O(N__25035),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_7));
    CascadeMux I__2766 (
            .O(N__25032),
            .I(N__25029));
    InMux I__2765 (
            .O(N__25029),
            .I(N__25026));
    LocalMux I__2764 (
            .O(N__25026),
            .I(N__25023));
    Span4Mux_h I__2763 (
            .O(N__25023),
            .I(N__25020));
    Span4Mux_h I__2762 (
            .O(N__25020),
            .I(N__25017));
    Odrv4 I__2761 (
            .O(N__25017),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_7 ));
    InMux I__2760 (
            .O(N__25014),
            .I(N__25011));
    LocalMux I__2759 (
            .O(N__25011),
            .I(N__25008));
    Odrv4 I__2758 (
            .O(N__25008),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_7 ));
    CascadeMux I__2757 (
            .O(N__25005),
            .I(N__25001));
    CascadeMux I__2756 (
            .O(N__25004),
            .I(N__24998));
    CascadeBuf I__2755 (
            .O(N__25001),
            .I(N__24995));
    CascadeBuf I__2754 (
            .O(N__24998),
            .I(N__24992));
    CascadeMux I__2753 (
            .O(N__24995),
            .I(N__24989));
    CascadeMux I__2752 (
            .O(N__24992),
            .I(N__24986));
    CascadeBuf I__2751 (
            .O(N__24989),
            .I(N__24983));
    CascadeBuf I__2750 (
            .O(N__24986),
            .I(N__24980));
    CascadeMux I__2749 (
            .O(N__24983),
            .I(N__24977));
    CascadeMux I__2748 (
            .O(N__24980),
            .I(N__24974));
    CascadeBuf I__2747 (
            .O(N__24977),
            .I(N__24971));
    CascadeBuf I__2746 (
            .O(N__24974),
            .I(N__24968));
    CascadeMux I__2745 (
            .O(N__24971),
            .I(N__24965));
    CascadeMux I__2744 (
            .O(N__24968),
            .I(N__24962));
    CascadeBuf I__2743 (
            .O(N__24965),
            .I(N__24959));
    CascadeBuf I__2742 (
            .O(N__24962),
            .I(N__24956));
    CascadeMux I__2741 (
            .O(N__24959),
            .I(N__24953));
    CascadeMux I__2740 (
            .O(N__24956),
            .I(N__24950));
    CascadeBuf I__2739 (
            .O(N__24953),
            .I(N__24947));
    CascadeBuf I__2738 (
            .O(N__24950),
            .I(N__24944));
    CascadeMux I__2737 (
            .O(N__24947),
            .I(N__24941));
    CascadeMux I__2736 (
            .O(N__24944),
            .I(N__24938));
    CascadeBuf I__2735 (
            .O(N__24941),
            .I(N__24935));
    CascadeBuf I__2734 (
            .O(N__24938),
            .I(N__24932));
    CascadeMux I__2733 (
            .O(N__24935),
            .I(N__24929));
    CascadeMux I__2732 (
            .O(N__24932),
            .I(N__24926));
    CascadeBuf I__2731 (
            .O(N__24929),
            .I(N__24923));
    CascadeBuf I__2730 (
            .O(N__24926),
            .I(N__24920));
    CascadeMux I__2729 (
            .O(N__24923),
            .I(N__24917));
    CascadeMux I__2728 (
            .O(N__24920),
            .I(N__24914));
    InMux I__2727 (
            .O(N__24917),
            .I(N__24911));
    InMux I__2726 (
            .O(N__24914),
            .I(N__24908));
    LocalMux I__2725 (
            .O(N__24911),
            .I(N__24905));
    LocalMux I__2724 (
            .O(N__24908),
            .I(N__24902));
    Span4Mux_h I__2723 (
            .O(N__24905),
            .I(N__24899));
    Span4Mux_h I__2722 (
            .O(N__24902),
            .I(N__24896));
    Odrv4 I__2721 (
            .O(N__24899),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4 ));
    Odrv4 I__2720 (
            .O(N__24896),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4 ));
    CEMux I__2719 (
            .O(N__24891),
            .I(N__24888));
    LocalMux I__2718 (
            .O(N__24888),
            .I(N__24884));
    CEMux I__2717 (
            .O(N__24887),
            .I(N__24881));
    Span4Mux_h I__2716 (
            .O(N__24884),
            .I(N__24876));
    LocalMux I__2715 (
            .O(N__24881),
            .I(N__24876));
    Odrv4 I__2714 (
            .O(N__24876),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1827_0 ));
    CascadeMux I__2713 (
            .O(N__24873),
            .I(N__24870));
    InMux I__2712 (
            .O(N__24870),
            .I(N__24867));
    LocalMux I__2711 (
            .O(N__24867),
            .I(N__24864));
    Span4Mux_h I__2710 (
            .O(N__24864),
            .I(N__24861));
    Span4Mux_v I__2709 (
            .O(N__24861),
            .I(N__24858));
    Odrv4 I__2708 (
            .O(N__24858),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_7));
    CascadeMux I__2707 (
            .O(N__24855),
            .I(N__24852));
    InMux I__2706 (
            .O(N__24852),
            .I(N__24849));
    LocalMux I__2705 (
            .O(N__24849),
            .I(N__24846));
    Span4Mux_h I__2704 (
            .O(N__24846),
            .I(N__24843));
    Odrv4 I__2703 (
            .O(N__24843),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.N_863 ));
    IoInMux I__2702 (
            .O(N__24840),
            .I(N__24837));
    LocalMux I__2701 (
            .O(N__24837),
            .I(N__24833));
    IoInMux I__2700 (
            .O(N__24836),
            .I(N__24830));
    IoSpan4Mux I__2699 (
            .O(N__24833),
            .I(N__24825));
    LocalMux I__2698 (
            .O(N__24830),
            .I(N__24825));
    IoSpan4Mux I__2697 (
            .O(N__24825),
            .I(N__24822));
    Span4Mux_s3_h I__2696 (
            .O(N__24822),
            .I(N__24819));
    Span4Mux_h I__2695 (
            .O(N__24819),
            .I(N__24815));
    InMux I__2694 (
            .O(N__24818),
            .I(N__24812));
    Odrv4 I__2693 (
            .O(N__24815),
            .I(s1_c));
    LocalMux I__2692 (
            .O(N__24812),
            .I(s1_c));
    CascadeMux I__2691 (
            .O(N__24807),
            .I(N__24804));
    CascadeBuf I__2690 (
            .O(N__24804),
            .I(N__24800));
    CascadeMux I__2689 (
            .O(N__24803),
            .I(N__24797));
    CascadeMux I__2688 (
            .O(N__24800),
            .I(N__24794));
    CascadeBuf I__2687 (
            .O(N__24797),
            .I(N__24791));
    CascadeBuf I__2686 (
            .O(N__24794),
            .I(N__24788));
    CascadeMux I__2685 (
            .O(N__24791),
            .I(N__24785));
    CascadeMux I__2684 (
            .O(N__24788),
            .I(N__24782));
    CascadeBuf I__2683 (
            .O(N__24785),
            .I(N__24779));
    CascadeBuf I__2682 (
            .O(N__24782),
            .I(N__24776));
    CascadeMux I__2681 (
            .O(N__24779),
            .I(N__24773));
    CascadeMux I__2680 (
            .O(N__24776),
            .I(N__24770));
    CascadeBuf I__2679 (
            .O(N__24773),
            .I(N__24767));
    CascadeBuf I__2678 (
            .O(N__24770),
            .I(N__24764));
    CascadeMux I__2677 (
            .O(N__24767),
            .I(N__24761));
    CascadeMux I__2676 (
            .O(N__24764),
            .I(N__24758));
    CascadeBuf I__2675 (
            .O(N__24761),
            .I(N__24755));
    CascadeBuf I__2674 (
            .O(N__24758),
            .I(N__24752));
    CascadeMux I__2673 (
            .O(N__24755),
            .I(N__24749));
    CascadeMux I__2672 (
            .O(N__24752),
            .I(N__24746));
    CascadeBuf I__2671 (
            .O(N__24749),
            .I(N__24743));
    CascadeBuf I__2670 (
            .O(N__24746),
            .I(N__24740));
    CascadeMux I__2669 (
            .O(N__24743),
            .I(N__24737));
    CascadeMux I__2668 (
            .O(N__24740),
            .I(N__24734));
    CascadeBuf I__2667 (
            .O(N__24737),
            .I(N__24731));
    CascadeBuf I__2666 (
            .O(N__24734),
            .I(N__24728));
    CascadeMux I__2665 (
            .O(N__24731),
            .I(N__24725));
    CascadeMux I__2664 (
            .O(N__24728),
            .I(N__24722));
    CascadeBuf I__2663 (
            .O(N__24725),
            .I(N__24719));
    InMux I__2662 (
            .O(N__24722),
            .I(N__24716));
    CascadeMux I__2661 (
            .O(N__24719),
            .I(N__24713));
    LocalMux I__2660 (
            .O(N__24716),
            .I(N__24710));
    InMux I__2659 (
            .O(N__24713),
            .I(N__24707));
    Odrv4 I__2658 (
            .O(N__24710),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5 ));
    LocalMux I__2657 (
            .O(N__24707),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5 ));
    InMux I__2656 (
            .O(N__24702),
            .I(N__24699));
    LocalMux I__2655 (
            .O(N__24699),
            .I(N__24694));
    InMux I__2654 (
            .O(N__24698),
            .I(N__24691));
    InMux I__2653 (
            .O(N__24697),
            .I(N__24688));
    Span4Mux_s3_v I__2652 (
            .O(N__24694),
            .I(N__24683));
    LocalMux I__2651 (
            .O(N__24691),
            .I(N__24683));
    LocalMux I__2650 (
            .O(N__24688),
            .I(N__24680));
    Span4Mux_v I__2649 (
            .O(N__24683),
            .I(N__24674));
    Span4Mux_v I__2648 (
            .O(N__24680),
            .I(N__24674));
    InMux I__2647 (
            .O(N__24679),
            .I(N__24671));
    Odrv4 I__2646 (
            .O(N__24674),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0 ));
    LocalMux I__2645 (
            .O(N__24671),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0 ));
    InMux I__2644 (
            .O(N__24666),
            .I(N__24662));
    InMux I__2643 (
            .O(N__24665),
            .I(N__24658));
    LocalMux I__2642 (
            .O(N__24662),
            .I(N__24654));
    InMux I__2641 (
            .O(N__24661),
            .I(N__24651));
    LocalMux I__2640 (
            .O(N__24658),
            .I(N__24648));
    InMux I__2639 (
            .O(N__24657),
            .I(N__24645));
    Span4Mux_h I__2638 (
            .O(N__24654),
            .I(N__24642));
    LocalMux I__2637 (
            .O(N__24651),
            .I(N__24639));
    Span4Mux_v I__2636 (
            .O(N__24648),
            .I(N__24634));
    LocalMux I__2635 (
            .O(N__24645),
            .I(N__24634));
    Span4Mux_v I__2634 (
            .O(N__24642),
            .I(N__24629));
    Span4Mux_h I__2633 (
            .O(N__24639),
            .I(N__24629));
    Odrv4 I__2632 (
            .O(N__24634),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0 ));
    Odrv4 I__2631 (
            .O(N__24629),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0 ));
    InMux I__2630 (
            .O(N__24624),
            .I(N__24621));
    LocalMux I__2629 (
            .O(N__24621),
            .I(N__24616));
    InMux I__2628 (
            .O(N__24620),
            .I(N__24613));
    InMux I__2627 (
            .O(N__24619),
            .I(N__24610));
    Span4Mux_s3_v I__2626 (
            .O(N__24616),
            .I(N__24605));
    LocalMux I__2625 (
            .O(N__24613),
            .I(N__24605));
    LocalMux I__2624 (
            .O(N__24610),
            .I(N__24602));
    Span4Mux_v I__2623 (
            .O(N__24605),
            .I(N__24596));
    Span4Mux_v I__2622 (
            .O(N__24602),
            .I(N__24596));
    InMux I__2621 (
            .O(N__24601),
            .I(N__24593));
    Odrv4 I__2620 (
            .O(N__24596),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0 ));
    LocalMux I__2619 (
            .O(N__24593),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0 ));
    InMux I__2618 (
            .O(N__24588),
            .I(N__24585));
    LocalMux I__2617 (
            .O(N__24585),
            .I(N__24580));
    InMux I__2616 (
            .O(N__24584),
            .I(N__24577));
    InMux I__2615 (
            .O(N__24583),
            .I(N__24574));
    Span4Mux_s2_v I__2614 (
            .O(N__24580),
            .I(N__24571));
    LocalMux I__2613 (
            .O(N__24577),
            .I(N__24568));
    LocalMux I__2612 (
            .O(N__24574),
            .I(N__24565));
    Span4Mux_v I__2611 (
            .O(N__24571),
            .I(N__24557));
    Span4Mux_v I__2610 (
            .O(N__24568),
            .I(N__24557));
    Span4Mux_h I__2609 (
            .O(N__24565),
            .I(N__24557));
    InMux I__2608 (
            .O(N__24564),
            .I(N__24554));
    Odrv4 I__2607 (
            .O(N__24557),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0 ));
    LocalMux I__2606 (
            .O(N__24554),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0 ));
    CEMux I__2605 (
            .O(N__24549),
            .I(N__24545));
    CEMux I__2604 (
            .O(N__24548),
            .I(N__24542));
    LocalMux I__2603 (
            .O(N__24545),
            .I(N__24537));
    LocalMux I__2602 (
            .O(N__24542),
            .I(N__24537));
    Odrv4 I__2601 (
            .O(N__24537),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1826_0 ));
    InMux I__2600 (
            .O(N__24534),
            .I(N__24529));
    InMux I__2599 (
            .O(N__24533),
            .I(N__24526));
    InMux I__2598 (
            .O(N__24532),
            .I(N__24523));
    LocalMux I__2597 (
            .O(N__24529),
            .I(N__24520));
    LocalMux I__2596 (
            .O(N__24526),
            .I(N__24517));
    LocalMux I__2595 (
            .O(N__24523),
            .I(N__24514));
    Span4Mux_v I__2594 (
            .O(N__24520),
            .I(N__24510));
    Span4Mux_v I__2593 (
            .O(N__24517),
            .I(N__24505));
    Span4Mux_h I__2592 (
            .O(N__24514),
            .I(N__24505));
    InMux I__2591 (
            .O(N__24513),
            .I(N__24502));
    Odrv4 I__2590 (
            .O(N__24510),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0 ));
    Odrv4 I__2589 (
            .O(N__24505),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0 ));
    LocalMux I__2588 (
            .O(N__24502),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0 ));
    InMux I__2587 (
            .O(N__24495),
            .I(N__24492));
    LocalMux I__2586 (
            .O(N__24492),
            .I(N__24488));
    InMux I__2585 (
            .O(N__24491),
            .I(N__24485));
    Span4Mux_s2_v I__2584 (
            .O(N__24488),
            .I(N__24478));
    LocalMux I__2583 (
            .O(N__24485),
            .I(N__24478));
    InMux I__2582 (
            .O(N__24484),
            .I(N__24475));
    InMux I__2581 (
            .O(N__24483),
            .I(N__24472));
    Span4Mux_v I__2580 (
            .O(N__24478),
            .I(N__24467));
    LocalMux I__2579 (
            .O(N__24475),
            .I(N__24467));
    LocalMux I__2578 (
            .O(N__24472),
            .I(N__24464));
    Odrv4 I__2577 (
            .O(N__24467),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0 ));
    Odrv4 I__2576 (
            .O(N__24464),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0 ));
    InMux I__2575 (
            .O(N__24459),
            .I(N__24456));
    LocalMux I__2574 (
            .O(N__24456),
            .I(N__24453));
    Span4Mux_s2_v I__2573 (
            .O(N__24453),
            .I(N__24449));
    InMux I__2572 (
            .O(N__24452),
            .I(N__24446));
    Span4Mux_v I__2571 (
            .O(N__24449),
            .I(N__24440));
    LocalMux I__2570 (
            .O(N__24446),
            .I(N__24440));
    InMux I__2569 (
            .O(N__24445),
            .I(N__24437));
    Span4Mux_h I__2568 (
            .O(N__24440),
            .I(N__24434));
    LocalMux I__2567 (
            .O(N__24437),
            .I(N__24431));
    Span4Mux_v I__2566 (
            .O(N__24434),
            .I(N__24425));
    Span4Mux_v I__2565 (
            .O(N__24431),
            .I(N__24425));
    InMux I__2564 (
            .O(N__24430),
            .I(N__24422));
    Odrv4 I__2563 (
            .O(N__24425),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0 ));
    LocalMux I__2562 (
            .O(N__24422),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0 ));
    InMux I__2561 (
            .O(N__24417),
            .I(N__24414));
    LocalMux I__2560 (
            .O(N__24414),
            .I(N__24411));
    Odrv4 I__2559 (
            .O(N__24411),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_5));
    CascadeMux I__2558 (
            .O(N__24408),
            .I(N__24405));
    InMux I__2557 (
            .O(N__24405),
            .I(N__24402));
    LocalMux I__2556 (
            .O(N__24402),
            .I(N__24399));
    Span4Mux_h I__2555 (
            .O(N__24399),
            .I(N__24396));
    Odrv4 I__2554 (
            .O(N__24396),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_5 ));
    InMux I__2553 (
            .O(N__24393),
            .I(N__24388));
    InMux I__2552 (
            .O(N__24392),
            .I(N__24384));
    InMux I__2551 (
            .O(N__24391),
            .I(N__24381));
    LocalMux I__2550 (
            .O(N__24388),
            .I(N__24378));
    InMux I__2549 (
            .O(N__24387),
            .I(N__24375));
    LocalMux I__2548 (
            .O(N__24384),
            .I(N__24372));
    LocalMux I__2547 (
            .O(N__24381),
            .I(N__24369));
    Span4Mux_s3_v I__2546 (
            .O(N__24378),
            .I(N__24364));
    LocalMux I__2545 (
            .O(N__24375),
            .I(N__24364));
    Span4Mux_v I__2544 (
            .O(N__24372),
            .I(N__24359));
    Span4Mux_h I__2543 (
            .O(N__24369),
            .I(N__24359));
    Odrv4 I__2542 (
            .O(N__24364),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0 ));
    Odrv4 I__2541 (
            .O(N__24359),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0 ));
    InMux I__2540 (
            .O(N__24354),
            .I(N__24350));
    InMux I__2539 (
            .O(N__24353),
            .I(N__24346));
    LocalMux I__2538 (
            .O(N__24350),
            .I(N__24342));
    InMux I__2537 (
            .O(N__24349),
            .I(N__24339));
    LocalMux I__2536 (
            .O(N__24346),
            .I(N__24336));
    InMux I__2535 (
            .O(N__24345),
            .I(N__24333));
    Span4Mux_s3_v I__2534 (
            .O(N__24342),
            .I(N__24328));
    LocalMux I__2533 (
            .O(N__24339),
            .I(N__24328));
    Span4Mux_v I__2532 (
            .O(N__24336),
            .I(N__24323));
    LocalMux I__2531 (
            .O(N__24333),
            .I(N__24323));
    Odrv4 I__2530 (
            .O(N__24328),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0 ));
    Odrv4 I__2529 (
            .O(N__24323),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0 ));
    InMux I__2528 (
            .O(N__24318),
            .I(N__24314));
    InMux I__2527 (
            .O(N__24317),
            .I(N__24311));
    LocalMux I__2526 (
            .O(N__24314),
            .I(N__24307));
    LocalMux I__2525 (
            .O(N__24311),
            .I(N__24304));
    InMux I__2524 (
            .O(N__24310),
            .I(N__24301));
    Span4Mux_h I__2523 (
            .O(N__24307),
            .I(N__24298));
    Span4Mux_v I__2522 (
            .O(N__24304),
            .I(N__24293));
    LocalMux I__2521 (
            .O(N__24301),
            .I(N__24293));
    Span4Mux_v I__2520 (
            .O(N__24298),
            .I(N__24287));
    Span4Mux_v I__2519 (
            .O(N__24293),
            .I(N__24287));
    InMux I__2518 (
            .O(N__24292),
            .I(N__24284));
    Odrv4 I__2517 (
            .O(N__24287),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0 ));
    LocalMux I__2516 (
            .O(N__24284),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0 ));
    InMux I__2515 (
            .O(N__24279),
            .I(N__24276));
    LocalMux I__2514 (
            .O(N__24276),
            .I(N__24271));
    InMux I__2513 (
            .O(N__24275),
            .I(N__24268));
    InMux I__2512 (
            .O(N__24274),
            .I(N__24265));
    Span4Mux_s0_v I__2511 (
            .O(N__24271),
            .I(N__24262));
    LocalMux I__2510 (
            .O(N__24268),
            .I(N__24259));
    LocalMux I__2509 (
            .O(N__24265),
            .I(N__24256));
    Span4Mux_v I__2508 (
            .O(N__24262),
            .I(N__24248));
    Span4Mux_v I__2507 (
            .O(N__24259),
            .I(N__24248));
    Span4Mux_h I__2506 (
            .O(N__24256),
            .I(N__24248));
    InMux I__2505 (
            .O(N__24255),
            .I(N__24245));
    Odrv4 I__2504 (
            .O(N__24248),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0 ));
    LocalMux I__2503 (
            .O(N__24245),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0 ));
    InMux I__2502 (
            .O(N__24240),
            .I(N__24236));
    InMux I__2501 (
            .O(N__24239),
            .I(N__24232));
    LocalMux I__2500 (
            .O(N__24236),
            .I(N__24228));
    InMux I__2499 (
            .O(N__24235),
            .I(N__24225));
    LocalMux I__2498 (
            .O(N__24232),
            .I(N__24222));
    InMux I__2497 (
            .O(N__24231),
            .I(N__24219));
    Span4Mux_h I__2496 (
            .O(N__24228),
            .I(N__24216));
    LocalMux I__2495 (
            .O(N__24225),
            .I(N__24213));
    Span4Mux_v I__2494 (
            .O(N__24222),
            .I(N__24208));
    LocalMux I__2493 (
            .O(N__24219),
            .I(N__24208));
    Span4Mux_v I__2492 (
            .O(N__24216),
            .I(N__24203));
    Span4Mux_h I__2491 (
            .O(N__24213),
            .I(N__24203));
    Odrv4 I__2490 (
            .O(N__24208),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0 ));
    Odrv4 I__2489 (
            .O(N__24203),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0 ));
    InMux I__2488 (
            .O(N__24198),
            .I(N__24194));
    InMux I__2487 (
            .O(N__24197),
            .I(N__24190));
    LocalMux I__2486 (
            .O(N__24194),
            .I(N__24186));
    InMux I__2485 (
            .O(N__24193),
            .I(N__24183));
    LocalMux I__2484 (
            .O(N__24190),
            .I(N__24180));
    InMux I__2483 (
            .O(N__24189),
            .I(N__24177));
    Span4Mux_v I__2482 (
            .O(N__24186),
            .I(N__24172));
    LocalMux I__2481 (
            .O(N__24183),
            .I(N__24172));
    Span4Mux_v I__2480 (
            .O(N__24180),
            .I(N__24167));
    LocalMux I__2479 (
            .O(N__24177),
            .I(N__24167));
    Span4Mux_v I__2478 (
            .O(N__24172),
            .I(N__24164));
    Odrv4 I__2477 (
            .O(N__24167),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0 ));
    Odrv4 I__2476 (
            .O(N__24164),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0 ));
    InMux I__2475 (
            .O(N__24159),
            .I(N__24155));
    InMux I__2474 (
            .O(N__24158),
            .I(N__24151));
    LocalMux I__2473 (
            .O(N__24155),
            .I(N__24147));
    InMux I__2472 (
            .O(N__24154),
            .I(N__24144));
    LocalMux I__2471 (
            .O(N__24151),
            .I(N__24141));
    InMux I__2470 (
            .O(N__24150),
            .I(N__24138));
    Span4Mux_v I__2469 (
            .O(N__24147),
            .I(N__24133));
    LocalMux I__2468 (
            .O(N__24144),
            .I(N__24133));
    Span4Mux_v I__2467 (
            .O(N__24141),
            .I(N__24128));
    LocalMux I__2466 (
            .O(N__24138),
            .I(N__24128));
    Span4Mux_v I__2465 (
            .O(N__24133),
            .I(N__24123));
    Span4Mux_v I__2464 (
            .O(N__24128),
            .I(N__24123));
    Odrv4 I__2463 (
            .O(N__24123),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_448_0 ));
    InMux I__2462 (
            .O(N__24120),
            .I(N__24114));
    InMux I__2461 (
            .O(N__24119),
            .I(N__24111));
    InMux I__2460 (
            .O(N__24118),
            .I(N__24108));
    InMux I__2459 (
            .O(N__24117),
            .I(N__24105));
    LocalMux I__2458 (
            .O(N__24114),
            .I(N__24102));
    LocalMux I__2457 (
            .O(N__24111),
            .I(N__24099));
    LocalMux I__2456 (
            .O(N__24108),
            .I(N__24096));
    LocalMux I__2455 (
            .O(N__24105),
            .I(N__24093));
    Span4Mux_v I__2454 (
            .O(N__24102),
            .I(N__24090));
    Span4Mux_v I__2453 (
            .O(N__24099),
            .I(N__24083));
    Span4Mux_h I__2452 (
            .O(N__24096),
            .I(N__24083));
    Span4Mux_h I__2451 (
            .O(N__24093),
            .I(N__24083));
    Odrv4 I__2450 (
            .O(N__24090),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0 ));
    Odrv4 I__2449 (
            .O(N__24083),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0 ));
    InMux I__2448 (
            .O(N__24078),
            .I(N__24074));
    InMux I__2447 (
            .O(N__24077),
            .I(N__24070));
    LocalMux I__2446 (
            .O(N__24074),
            .I(N__24066));
    InMux I__2445 (
            .O(N__24073),
            .I(N__24063));
    LocalMux I__2444 (
            .O(N__24070),
            .I(N__24060));
    InMux I__2443 (
            .O(N__24069),
            .I(N__24057));
    Span4Mux_v I__2442 (
            .O(N__24066),
            .I(N__24052));
    LocalMux I__2441 (
            .O(N__24063),
            .I(N__24052));
    Span4Mux_v I__2440 (
            .O(N__24060),
            .I(N__24047));
    LocalMux I__2439 (
            .O(N__24057),
            .I(N__24047));
    Odrv4 I__2438 (
            .O(N__24052),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0 ));
    Odrv4 I__2437 (
            .O(N__24047),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0 ));
    InMux I__2436 (
            .O(N__24042),
            .I(N__24038));
    InMux I__2435 (
            .O(N__24041),
            .I(N__24034));
    LocalMux I__2434 (
            .O(N__24038),
            .I(N__24030));
    InMux I__2433 (
            .O(N__24037),
            .I(N__24027));
    LocalMux I__2432 (
            .O(N__24034),
            .I(N__24024));
    InMux I__2431 (
            .O(N__24033),
            .I(N__24021));
    Span4Mux_v I__2430 (
            .O(N__24030),
            .I(N__24016));
    LocalMux I__2429 (
            .O(N__24027),
            .I(N__24016));
    Span4Mux_s2_v I__2428 (
            .O(N__24024),
            .I(N__24011));
    LocalMux I__2427 (
            .O(N__24021),
            .I(N__24011));
    Odrv4 I__2426 (
            .O(N__24016),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0 ));
    Odrv4 I__2425 (
            .O(N__24011),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0 ));
    InMux I__2424 (
            .O(N__24006),
            .I(N__24002));
    InMux I__2423 (
            .O(N__24005),
            .I(N__23999));
    LocalMux I__2422 (
            .O(N__24002),
            .I(N__23995));
    LocalMux I__2421 (
            .O(N__23999),
            .I(N__23992));
    InMux I__2420 (
            .O(N__23998),
            .I(N__23988));
    Span4Mux_s0_v I__2419 (
            .O(N__23995),
            .I(N__23985));
    Span4Mux_h I__2418 (
            .O(N__23992),
            .I(N__23982));
    InMux I__2417 (
            .O(N__23991),
            .I(N__23979));
    LocalMux I__2416 (
            .O(N__23988),
            .I(N__23976));
    Span4Mux_v I__2415 (
            .O(N__23985),
            .I(N__23967));
    Span4Mux_v I__2414 (
            .O(N__23982),
            .I(N__23967));
    LocalMux I__2413 (
            .O(N__23979),
            .I(N__23967));
    Span4Mux_h I__2412 (
            .O(N__23976),
            .I(N__23967));
    Odrv4 I__2411 (
            .O(N__23967),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_459_0 ));
    InMux I__2410 (
            .O(N__23964),
            .I(N__23958));
    InMux I__2409 (
            .O(N__23963),
            .I(N__23955));
    InMux I__2408 (
            .O(N__23962),
            .I(N__23952));
    InMux I__2407 (
            .O(N__23961),
            .I(N__23949));
    LocalMux I__2406 (
            .O(N__23958),
            .I(N__23946));
    LocalMux I__2405 (
            .O(N__23955),
            .I(N__23943));
    LocalMux I__2404 (
            .O(N__23952),
            .I(N__23940));
    LocalMux I__2403 (
            .O(N__23949),
            .I(N__23937));
    Span4Mux_s2_v I__2402 (
            .O(N__23946),
            .I(N__23934));
    Span4Mux_v I__2401 (
            .O(N__23943),
            .I(N__23927));
    Span4Mux_h I__2400 (
            .O(N__23940),
            .I(N__23927));
    Span4Mux_h I__2399 (
            .O(N__23937),
            .I(N__23927));
    Odrv4 I__2398 (
            .O(N__23934),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0 ));
    Odrv4 I__2397 (
            .O(N__23927),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0 ));
    InMux I__2396 (
            .O(N__23922),
            .I(N__23917));
    InMux I__2395 (
            .O(N__23921),
            .I(N__23914));
    InMux I__2394 (
            .O(N__23920),
            .I(N__23910));
    LocalMux I__2393 (
            .O(N__23917),
            .I(N__23907));
    LocalMux I__2392 (
            .O(N__23914),
            .I(N__23904));
    InMux I__2391 (
            .O(N__23913),
            .I(N__23901));
    LocalMux I__2390 (
            .O(N__23910),
            .I(N__23898));
    Span4Mux_s3_v I__2389 (
            .O(N__23907),
            .I(N__23895));
    Span4Mux_v I__2388 (
            .O(N__23904),
            .I(N__23888));
    LocalMux I__2387 (
            .O(N__23901),
            .I(N__23888));
    Span4Mux_h I__2386 (
            .O(N__23898),
            .I(N__23888));
    Odrv4 I__2385 (
            .O(N__23895),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0 ));
    Odrv4 I__2384 (
            .O(N__23888),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0 ));
    InMux I__2383 (
            .O(N__23883),
            .I(N__23879));
    InMux I__2382 (
            .O(N__23882),
            .I(N__23875));
    LocalMux I__2381 (
            .O(N__23879),
            .I(N__23872));
    InMux I__2380 (
            .O(N__23878),
            .I(N__23869));
    LocalMux I__2379 (
            .O(N__23875),
            .I(N__23866));
    Span4Mux_v I__2378 (
            .O(N__23872),
            .I(N__23861));
    LocalMux I__2377 (
            .O(N__23869),
            .I(N__23861));
    Span4Mux_v I__2376 (
            .O(N__23866),
            .I(N__23855));
    Span4Mux_v I__2375 (
            .O(N__23861),
            .I(N__23855));
    InMux I__2374 (
            .O(N__23860),
            .I(N__23852));
    Odrv4 I__2373 (
            .O(N__23855),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0 ));
    LocalMux I__2372 (
            .O(N__23852),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0 ));
    InMux I__2371 (
            .O(N__23847),
            .I(N__23844));
    LocalMux I__2370 (
            .O(N__23844),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_8));
    InMux I__2369 (
            .O(N__23841),
            .I(N__23837));
    InMux I__2368 (
            .O(N__23840),
            .I(N__23833));
    LocalMux I__2367 (
            .O(N__23837),
            .I(N__23830));
    InMux I__2366 (
            .O(N__23836),
            .I(N__23827));
    LocalMux I__2365 (
            .O(N__23833),
            .I(N__23824));
    Span4Mux_v I__2364 (
            .O(N__23830),
            .I(N__23819));
    LocalMux I__2363 (
            .O(N__23827),
            .I(N__23819));
    Span4Mux_h I__2362 (
            .O(N__23824),
            .I(N__23815));
    Span4Mux_v I__2361 (
            .O(N__23819),
            .I(N__23812));
    InMux I__2360 (
            .O(N__23818),
            .I(N__23809));
    Odrv4 I__2359 (
            .O(N__23815),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0 ));
    Odrv4 I__2358 (
            .O(N__23812),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0 ));
    LocalMux I__2357 (
            .O(N__23809),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0 ));
    CascadeMux I__2356 (
            .O(N__23802),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0_cascade_ ));
    InMux I__2355 (
            .O(N__23799),
            .I(N__23795));
    InMux I__2354 (
            .O(N__23798),
            .I(N__23791));
    LocalMux I__2353 (
            .O(N__23795),
            .I(N__23787));
    InMux I__2352 (
            .O(N__23794),
            .I(N__23784));
    LocalMux I__2351 (
            .O(N__23791),
            .I(N__23781));
    InMux I__2350 (
            .O(N__23790),
            .I(N__23778));
    Span4Mux_s3_v I__2349 (
            .O(N__23787),
            .I(N__23773));
    LocalMux I__2348 (
            .O(N__23784),
            .I(N__23773));
    Span4Mux_v I__2347 (
            .O(N__23781),
            .I(N__23768));
    LocalMux I__2346 (
            .O(N__23778),
            .I(N__23768));
    Span4Mux_v I__2345 (
            .O(N__23773),
            .I(N__23763));
    Span4Mux_v I__2344 (
            .O(N__23768),
            .I(N__23763));
    Odrv4 I__2343 (
            .O(N__23763),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_466_0 ));
    CascadeMux I__2342 (
            .O(N__23760),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.csb_u_i_a2_0_0_cascade_ ));
    CascadeMux I__2341 (
            .O(N__23757),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_331_cascade_ ));
    CascadeMux I__2340 (
            .O(N__23754),
            .I(N__23751));
    InMux I__2339 (
            .O(N__23751),
            .I(N__23748));
    LocalMux I__2338 (
            .O(N__23748),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_0 ));
    InMux I__2337 (
            .O(N__23745),
            .I(N__23742));
    LocalMux I__2336 (
            .O(N__23742),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.m7_0_a2_3 ));
    CEMux I__2335 (
            .O(N__23739),
            .I(N__23736));
    LocalMux I__2334 (
            .O(N__23736),
            .I(N__23733));
    Span4Mux_v I__2333 (
            .O(N__23733),
            .I(N__23729));
    CEMux I__2332 (
            .O(N__23732),
            .I(N__23726));
    Odrv4 I__2331 (
            .O(N__23729),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0 ));
    LocalMux I__2330 (
            .O(N__23726),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0 ));
    InMux I__2329 (
            .O(N__23721),
            .I(N__23717));
    InMux I__2328 (
            .O(N__23720),
            .I(N__23713));
    LocalMux I__2327 (
            .O(N__23717),
            .I(N__23710));
    InMux I__2326 (
            .O(N__23716),
            .I(N__23707));
    LocalMux I__2325 (
            .O(N__23713),
            .I(N__23704));
    Span4Mux_v I__2324 (
            .O(N__23710),
            .I(N__23699));
    LocalMux I__2323 (
            .O(N__23707),
            .I(N__23699));
    Span4Mux_v I__2322 (
            .O(N__23704),
            .I(N__23693));
    Span4Mux_v I__2321 (
            .O(N__23699),
            .I(N__23693));
    InMux I__2320 (
            .O(N__23698),
            .I(N__23690));
    Odrv4 I__2319 (
            .O(N__23693),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0 ));
    LocalMux I__2318 (
            .O(N__23690),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0 ));
    InMux I__2317 (
            .O(N__23685),
            .I(N__23681));
    InMux I__2316 (
            .O(N__23684),
            .I(N__23678));
    LocalMux I__2315 (
            .O(N__23681),
            .I(N__23674));
    LocalMux I__2314 (
            .O(N__23678),
            .I(N__23671));
    InMux I__2313 (
            .O(N__23677),
            .I(N__23668));
    Span4Mux_s1_v I__2312 (
            .O(N__23674),
            .I(N__23665));
    Span4Mux_v I__2311 (
            .O(N__23671),
            .I(N__23660));
    LocalMux I__2310 (
            .O(N__23668),
            .I(N__23660));
    Span4Mux_v I__2309 (
            .O(N__23665),
            .I(N__23654));
    Span4Mux_v I__2308 (
            .O(N__23660),
            .I(N__23654));
    InMux I__2307 (
            .O(N__23659),
            .I(N__23651));
    Odrv4 I__2306 (
            .O(N__23654),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0 ));
    LocalMux I__2305 (
            .O(N__23651),
            .I(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0 ));
    CascadeMux I__2304 (
            .O(N__23646),
            .I(N__23643));
    InMux I__2303 (
            .O(N__23643),
            .I(N__23640));
    LocalMux I__2302 (
            .O(N__23640),
            .I(N__23637));
    Span4Mux_h I__2301 (
            .O(N__23637),
            .I(N__23634));
    Span4Mux_v I__2300 (
            .O(N__23634),
            .I(N__23631));
    Span4Mux_v I__2299 (
            .O(N__23631),
            .I(N__23628));
    Odrv4 I__2298 (
            .O(N__23628),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_CO ));
    InMux I__2297 (
            .O(N__23625),
            .I(N__23622));
    LocalMux I__2296 (
            .O(N__23622),
            .I(N__23618));
    InMux I__2295 (
            .O(N__23621),
            .I(N__23615));
    Span4Mux_v I__2294 (
            .O(N__23618),
            .I(N__23610));
    LocalMux I__2293 (
            .O(N__23615),
            .I(N__23610));
    Span4Mux_h I__2292 (
            .O(N__23610),
            .I(N__23607));
    Span4Mux_v I__2291 (
            .O(N__23607),
            .I(N__23603));
    InMux I__2290 (
            .O(N__23606),
            .I(N__23600));
    Span4Mux_v I__2289 (
            .O(N__23603),
            .I(N__23597));
    LocalMux I__2288 (
            .O(N__23600),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2 ));
    Odrv4 I__2287 (
            .O(N__23597),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2 ));
    CascadeMux I__2286 (
            .O(N__23592),
            .I(N__23588));
    InMux I__2285 (
            .O(N__23591),
            .I(N__23582));
    InMux I__2284 (
            .O(N__23588),
            .I(N__23582));
    InMux I__2283 (
            .O(N__23587),
            .I(N__23579));
    LocalMux I__2282 (
            .O(N__23582),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15 ));
    LocalMux I__2281 (
            .O(N__23579),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15 ));
    InMux I__2280 (
            .O(N__23574),
            .I(N__23568));
    InMux I__2279 (
            .O(N__23573),
            .I(N__23568));
    LocalMux I__2278 (
            .O(N__23568),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_13 ));
    InMux I__2277 (
            .O(N__23565),
            .I(N__23560));
    InMux I__2276 (
            .O(N__23564),
            .I(N__23557));
    InMux I__2275 (
            .O(N__23563),
            .I(N__23554));
    LocalMux I__2274 (
            .O(N__23560),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2 ));
    LocalMux I__2273 (
            .O(N__23557),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2 ));
    LocalMux I__2272 (
            .O(N__23554),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2 ));
    InMux I__2271 (
            .O(N__23547),
            .I(N__23542));
    InMux I__2270 (
            .O(N__23546),
            .I(N__23539));
    InMux I__2269 (
            .O(N__23545),
            .I(N__23536));
    LocalMux I__2268 (
            .O(N__23542),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1 ));
    LocalMux I__2267 (
            .O(N__23539),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1 ));
    LocalMux I__2266 (
            .O(N__23536),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1 ));
    CascadeMux I__2265 (
            .O(N__23529),
            .I(N__23524));
    InMux I__2264 (
            .O(N__23528),
            .I(N__23521));
    InMux I__2263 (
            .O(N__23527),
            .I(N__23518));
    InMux I__2262 (
            .O(N__23524),
            .I(N__23515));
    LocalMux I__2261 (
            .O(N__23521),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3 ));
    LocalMux I__2260 (
            .O(N__23518),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3 ));
    LocalMux I__2259 (
            .O(N__23515),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3 ));
    InMux I__2258 (
            .O(N__23508),
            .I(N__23503));
    InMux I__2257 (
            .O(N__23507),
            .I(N__23500));
    InMux I__2256 (
            .O(N__23506),
            .I(N__23497));
    LocalMux I__2255 (
            .O(N__23503),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0 ));
    LocalMux I__2254 (
            .O(N__23500),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0 ));
    LocalMux I__2253 (
            .O(N__23497),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0 ));
    CascadeMux I__2252 (
            .O(N__23490),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383_cascade_ ));
    InMux I__2251 (
            .O(N__23487),
            .I(N__23480));
    InMux I__2250 (
            .O(N__23486),
            .I(N__23480));
    InMux I__2249 (
            .O(N__23485),
            .I(N__23477));
    LocalMux I__2248 (
            .O(N__23480),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0 ));
    LocalMux I__2247 (
            .O(N__23477),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0 ));
    CascadeMux I__2246 (
            .O(N__23472),
            .I(N__23468));
    InMux I__2245 (
            .O(N__23471),
            .I(N__23463));
    InMux I__2244 (
            .O(N__23468),
            .I(N__23463));
    LocalMux I__2243 (
            .O(N__23463),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_16 ));
    CascadeMux I__2242 (
            .O(N__23460),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_369_cascade_ ));
    InMux I__2241 (
            .O(N__23457),
            .I(N__23454));
    LocalMux I__2240 (
            .O(N__23454),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_12 ));
    CascadeMux I__2239 (
            .O(N__23451),
            .I(N__23443));
    InMux I__2238 (
            .O(N__23450),
            .I(N__23438));
    InMux I__2237 (
            .O(N__23449),
            .I(N__23433));
    InMux I__2236 (
            .O(N__23448),
            .I(N__23433));
    InMux I__2235 (
            .O(N__23447),
            .I(N__23428));
    InMux I__2234 (
            .O(N__23446),
            .I(N__23428));
    InMux I__2233 (
            .O(N__23443),
            .I(N__23425));
    InMux I__2232 (
            .O(N__23442),
            .I(N__23422));
    InMux I__2231 (
            .O(N__23441),
            .I(N__23419));
    LocalMux I__2230 (
            .O(N__23438),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ));
    LocalMux I__2229 (
            .O(N__23433),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ));
    LocalMux I__2228 (
            .O(N__23428),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ));
    LocalMux I__2227 (
            .O(N__23425),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ));
    LocalMux I__2226 (
            .O(N__23422),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ));
    LocalMux I__2225 (
            .O(N__23419),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ));
    InMux I__2224 (
            .O(N__23406),
            .I(N__23395));
    InMux I__2223 (
            .O(N__23405),
            .I(N__23395));
    InMux I__2222 (
            .O(N__23404),
            .I(N__23395));
    InMux I__2221 (
            .O(N__23403),
            .I(N__23390));
    InMux I__2220 (
            .O(N__23402),
            .I(N__23390));
    LocalMux I__2219 (
            .O(N__23395),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383 ));
    LocalMux I__2218 (
            .O(N__23390),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383 ));
    InMux I__2217 (
            .O(N__23385),
            .I(N__23378));
    InMux I__2216 (
            .O(N__23384),
            .I(N__23378));
    InMux I__2215 (
            .O(N__23383),
            .I(N__23375));
    LocalMux I__2214 (
            .O(N__23378),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7 ));
    LocalMux I__2213 (
            .O(N__23375),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7 ));
    InMux I__2212 (
            .O(N__23370),
            .I(N__23367));
    LocalMux I__2211 (
            .O(N__23367),
            .I(N__23363));
    CascadeMux I__2210 (
            .O(N__23366),
            .I(N__23360));
    Span4Mux_h I__2209 (
            .O(N__23363),
            .I(N__23357));
    InMux I__2208 (
            .O(N__23360),
            .I(N__23354));
    Odrv4 I__2207 (
            .O(N__23357),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16 ));
    LocalMux I__2206 (
            .O(N__23354),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16 ));
    InMux I__2205 (
            .O(N__23349),
            .I(N__23344));
    InMux I__2204 (
            .O(N__23348),
            .I(N__23341));
    InMux I__2203 (
            .O(N__23347),
            .I(N__23338));
    LocalMux I__2202 (
            .O(N__23344),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0 ));
    LocalMux I__2201 (
            .O(N__23341),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0 ));
    LocalMux I__2200 (
            .O(N__23338),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0 ));
    CascadeMux I__2199 (
            .O(N__23331),
            .I(N__23328));
    InMux I__2198 (
            .O(N__23328),
            .I(N__23325));
    LocalMux I__2197 (
            .O(N__23325),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_0 ));
    CascadeMux I__2196 (
            .O(N__23322),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0_cascade_ ));
    InMux I__2195 (
            .O(N__23319),
            .I(N__23316));
    LocalMux I__2194 (
            .O(N__23316),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_4 ));
    CascadeMux I__2193 (
            .O(N__23313),
            .I(N__23310));
    InMux I__2192 (
            .O(N__23310),
            .I(N__23304));
    InMux I__2191 (
            .O(N__23309),
            .I(N__23304));
    LocalMux I__2190 (
            .O(N__23304),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_5 ));
    CascadeMux I__2189 (
            .O(N__23301),
            .I(N__23298));
    InMux I__2188 (
            .O(N__23298),
            .I(N__23292));
    InMux I__2187 (
            .O(N__23297),
            .I(N__23292));
    LocalMux I__2186 (
            .O(N__23292),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_8 ));
    InMux I__2185 (
            .O(N__23289),
            .I(N__23285));
    InMux I__2184 (
            .O(N__23288),
            .I(N__23282));
    LocalMux I__2183 (
            .O(N__23285),
            .I(N__23279));
    LocalMux I__2182 (
            .O(N__23282),
            .I(N__23276));
    Span4Mux_h I__2181 (
            .O(N__23279),
            .I(N__23273));
    Odrv4 I__2180 (
            .O(N__23276),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15 ));
    Odrv4 I__2179 (
            .O(N__23273),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15 ));
    CascadeMux I__2178 (
            .O(N__23268),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1Z0Z_23_cascade_ ));
    IoInMux I__2177 (
            .O(N__23265),
            .I(N__23262));
    LocalMux I__2176 (
            .O(N__23262),
            .I(N__23259));
    IoSpan4Mux I__2175 (
            .O(N__23259),
            .I(N__23256));
    Span4Mux_s0_v I__2174 (
            .O(N__23256),
            .I(N__23253));
    Span4Mux_v I__2173 (
            .O(N__23253),
            .I(N__23250));
    Sp12to4 I__2172 (
            .O(N__23250),
            .I(N__23247));
    Odrv12 I__2171 (
            .O(N__23247),
            .I(N_29));
    InMux I__2170 (
            .O(N__23244),
            .I(N__23241));
    LocalMux I__2169 (
            .O(N__23241),
            .I(N__23238));
    Span4Mux_h I__2168 (
            .O(N__23238),
            .I(N__23235));
    Odrv4 I__2167 (
            .O(N__23235),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_read ));
    InMux I__2166 (
            .O(N__23232),
            .I(N__23229));
    LocalMux I__2165 (
            .O(N__23229),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01Z0Z_0 ));
    InMux I__2164 (
            .O(N__23226),
            .I(N__23223));
    LocalMux I__2163 (
            .O(N__23223),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_reti_0_1 ));
    InMux I__2162 (
            .O(N__23220),
            .I(N__23217));
    LocalMux I__2161 (
            .O(N__23217),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0 ));
    CascadeMux I__2160 (
            .O(N__23214),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0_cascade_ ));
    InMux I__2159 (
            .O(N__23211),
            .I(N__23208));
    LocalMux I__2158 (
            .O(N__23208),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.sclk_u_i_0 ));
    InMux I__2157 (
            .O(N__23205),
            .I(N__23202));
    LocalMux I__2156 (
            .O(N__23202),
            .I(N__23199));
    Sp12to4 I__2155 (
            .O(N__23199),
            .I(N__23196));
    Span12Mux_v I__2154 (
            .O(N__23196),
            .I(N__23193));
    Odrv12 I__2153 (
            .O(N__23193),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_7));
    CascadeMux I__2152 (
            .O(N__23190),
            .I(N__23187));
    InMux I__2151 (
            .O(N__23187),
            .I(N__23184));
    LocalMux I__2150 (
            .O(N__23184),
            .I(N__23181));
    Span4Mux_h I__2149 (
            .O(N__23181),
            .I(N__23178));
    Span4Mux_v I__2148 (
            .O(N__23178),
            .I(N__23175));
    Odrv4 I__2147 (
            .O(N__23175),
            .I(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_7));
    CascadeMux I__2146 (
            .O(N__23172),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_7_cascade_ ));
    InMux I__2145 (
            .O(N__23169),
            .I(N__23166));
    LocalMux I__2144 (
            .O(N__23166),
            .I(N__23163));
    Span4Mux_h I__2143 (
            .O(N__23163),
            .I(N__23160));
    Odrv4 I__2142 (
            .O(N__23160),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_7 ));
    CascadeMux I__2141 (
            .O(N__23157),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_7_cascade_ ));
    InMux I__2140 (
            .O(N__23154),
            .I(N__23151));
    LocalMux I__2139 (
            .O(N__23151),
            .I(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_7 ));
    InMux I__2138 (
            .O(N__23148),
            .I(N__23145));
    LocalMux I__2137 (
            .O(N__23145),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.dout_read ));
    CascadeMux I__2136 (
            .O(N__23142),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_237_cascade_ ));
    IoInMux I__2135 (
            .O(N__23139),
            .I(N__23136));
    LocalMux I__2134 (
            .O(N__23136),
            .I(N__23133));
    Span4Mux_s2_h I__2133 (
            .O(N__23133),
            .I(N__23130));
    Span4Mux_v I__2132 (
            .O(N__23130),
            .I(N__23127));
    Odrv4 I__2131 (
            .O(N__23127),
            .I(N_85_0));
    InMux I__2130 (
            .O(N__23124),
            .I(N__23121));
    LocalMux I__2129 (
            .O(N__23121),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_6 ));
    InMux I__2128 (
            .O(N__23118),
            .I(N__23115));
    LocalMux I__2127 (
            .O(N__23115),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_5 ));
    InMux I__2126 (
            .O(N__23112),
            .I(N__23109));
    LocalMux I__2125 (
            .O(N__23109),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_4 ));
    InMux I__2124 (
            .O(N__23106),
            .I(N__23103));
    LocalMux I__2123 (
            .O(N__23103),
            .I(N__23100));
    Span4Mux_v I__2122 (
            .O(N__23100),
            .I(N__23097));
    Odrv4 I__2121 (
            .O(N__23097),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_2 ));
    InMux I__2120 (
            .O(N__23094),
            .I(N__23091));
    LocalMux I__2119 (
            .O(N__23091),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_3 ));
    CEMux I__2118 (
            .O(N__23088),
            .I(N__23084));
    CEMux I__2117 (
            .O(N__23087),
            .I(N__23081));
    LocalMux I__2116 (
            .O(N__23084),
            .I(N__23078));
    LocalMux I__2115 (
            .O(N__23081),
            .I(N__23075));
    Span4Mux_v I__2114 (
            .O(N__23078),
            .I(N__23070));
    Span4Mux_h I__2113 (
            .O(N__23075),
            .I(N__23070));
    Span4Mux_s3_h I__2112 (
            .O(N__23070),
            .I(N__23067));
    Odrv4 I__2111 (
            .O(N__23067),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_370_i ));
    IoInMux I__2110 (
            .O(N__23064),
            .I(N__23061));
    LocalMux I__2109 (
            .O(N__23061),
            .I(N__23058));
    IoSpan4Mux I__2108 (
            .O(N__23058),
            .I(N__23055));
    Span4Mux_s2_v I__2107 (
            .O(N__23055),
            .I(N__23052));
    Sp12to4 I__2106 (
            .O(N__23052),
            .I(N__23049));
    Odrv12 I__2105 (
            .O(N__23049),
            .I(N_1820_0));
    InMux I__2104 (
            .O(N__23046),
            .I(N__23043));
    LocalMux I__2103 (
            .O(N__23043),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_u_i_0 ));
    InMux I__2102 (
            .O(N__23040),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2 ));
    InMux I__2101 (
            .O(N__23037),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_3 ));
    CascadeMux I__2100 (
            .O(N__23034),
            .I(N__23031));
    InMux I__2099 (
            .O(N__23031),
            .I(N__23028));
    LocalMux I__2098 (
            .O(N__23028),
            .I(N__23025));
    Odrv4 I__2097 (
            .O(N__23025),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_333 ));
    InMux I__2096 (
            .O(N__23022),
            .I(N__23019));
    LocalMux I__2095 (
            .O(N__23019),
            .I(N__23016));
    Span4Mux_h I__2094 (
            .O(N__23016),
            .I(N__23012));
    InMux I__2093 (
            .O(N__23015),
            .I(N__23009));
    Sp12to4 I__2092 (
            .O(N__23012),
            .I(N__23004));
    LocalMux I__2091 (
            .O(N__23009),
            .I(N__23004));
    Odrv12 I__2090 (
            .O(N__23004),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_376 ));
    CascadeMux I__2089 (
            .O(N__23001),
            .I(N__22998));
    InMux I__2088 (
            .O(N__22998),
            .I(N__22995));
    LocalMux I__2087 (
            .O(N__22995),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1 ));
    CascadeMux I__2086 (
            .O(N__22992),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1_cascade_ ));
    InMux I__2085 (
            .O(N__22989),
            .I(N__22978));
    InMux I__2084 (
            .O(N__22988),
            .I(N__22978));
    InMux I__2083 (
            .O(N__22987),
            .I(N__22978));
    InMux I__2082 (
            .O(N__22986),
            .I(N__22973));
    InMux I__2081 (
            .O(N__22985),
            .I(N__22973));
    LocalMux I__2080 (
            .O(N__22978),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0 ));
    LocalMux I__2079 (
            .O(N__22973),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0 ));
    InMux I__2078 (
            .O(N__22968),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0 ));
    InMux I__2077 (
            .O(N__22965),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1 ));
    InMux I__2076 (
            .O(N__22962),
            .I(N__22958));
    InMux I__2075 (
            .O(N__22961),
            .I(N__22954));
    LocalMux I__2074 (
            .O(N__22958),
            .I(N__22951));
    InMux I__2073 (
            .O(N__22957),
            .I(N__22948));
    LocalMux I__2072 (
            .O(N__22954),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3 ));
    Odrv4 I__2071 (
            .O(N__22951),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3 ));
    LocalMux I__2070 (
            .O(N__22948),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3 ));
    CascadeMux I__2069 (
            .O(N__22941),
            .I(N__22938));
    InMux I__2068 (
            .O(N__22938),
            .I(N__22935));
    LocalMux I__2067 (
            .O(N__22935),
            .I(N__22932));
    Odrv4 I__2066 (
            .O(N__22932),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_CO ));
    InMux I__2065 (
            .O(N__22929),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2 ));
    InMux I__2064 (
            .O(N__22926),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_3 ));
    InMux I__2063 (
            .O(N__22923),
            .I(N__22919));
    InMux I__2062 (
            .O(N__22922),
            .I(N__22916));
    LocalMux I__2061 (
            .O(N__22919),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4 ));
    LocalMux I__2060 (
            .O(N__22916),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4 ));
    InMux I__2059 (
            .O(N__22911),
            .I(bfn_6_19_0_));
    InMux I__2058 (
            .O(N__22908),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0 ));
    InMux I__2057 (
            .O(N__22905),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1 ));
    CascadeMux I__2056 (
            .O(N__22902),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93Z0Z_0_cascade_ ));
    IoInMux I__2055 (
            .O(N__22899),
            .I(N__22896));
    LocalMux I__2054 (
            .O(N__22896),
            .I(N__22893));
    Odrv12 I__2053 (
            .O(N__22893),
            .I(sclk1_c));
    InMux I__2052 (
            .O(N__22890),
            .I(N__22887));
    LocalMux I__2051 (
            .O(N__22887),
            .I(N__22884));
    Span4Mux_v I__2050 (
            .O(N__22884),
            .I(N__22879));
    InMux I__2049 (
            .O(N__22883),
            .I(N__22876));
    InMux I__2048 (
            .O(N__22882),
            .I(N__22873));
    Odrv4 I__2047 (
            .O(N__22879),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458 ));
    LocalMux I__2046 (
            .O(N__22876),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458 ));
    LocalMux I__2045 (
            .O(N__22873),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458 ));
    InMux I__2044 (
            .O(N__22866),
            .I(N__22863));
    LocalMux I__2043 (
            .O(N__22863),
            .I(N__22860));
    Span4Mux_v I__2042 (
            .O(N__22860),
            .I(N__22852));
    InMux I__2041 (
            .O(N__22859),
            .I(N__22847));
    InMux I__2040 (
            .O(N__22858),
            .I(N__22847));
    InMux I__2039 (
            .O(N__22857),
            .I(N__22840));
    InMux I__2038 (
            .O(N__22856),
            .I(N__22840));
    InMux I__2037 (
            .O(N__22855),
            .I(N__22840));
    Odrv4 I__2036 (
            .O(N__22852),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i ));
    LocalMux I__2035 (
            .O(N__22847),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i ));
    LocalMux I__2034 (
            .O(N__22840),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i ));
    InMux I__2033 (
            .O(N__22833),
            .I(N__22830));
    LocalMux I__2032 (
            .O(N__22830),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32Z0Z_0 ));
    CascadeMux I__2031 (
            .O(N__22827),
            .I(N__22822));
    InMux I__2030 (
            .O(N__22826),
            .I(N__22819));
    InMux I__2029 (
            .O(N__22825),
            .I(N__22816));
    InMux I__2028 (
            .O(N__22822),
            .I(N__22813));
    LocalMux I__2027 (
            .O(N__22819),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3 ));
    LocalMux I__2026 (
            .O(N__22816),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3 ));
    LocalMux I__2025 (
            .O(N__22813),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3 ));
    InMux I__2024 (
            .O(N__22806),
            .I(N__22801));
    InMux I__2023 (
            .O(N__22805),
            .I(N__22798));
    InMux I__2022 (
            .O(N__22804),
            .I(N__22795));
    LocalMux I__2021 (
            .O(N__22801),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2 ));
    LocalMux I__2020 (
            .O(N__22798),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2 ));
    LocalMux I__2019 (
            .O(N__22795),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2 ));
    InMux I__2018 (
            .O(N__22788),
            .I(N__22783));
    InMux I__2017 (
            .O(N__22787),
            .I(N__22780));
    InMux I__2016 (
            .O(N__22786),
            .I(N__22777));
    LocalMux I__2015 (
            .O(N__22783),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1 ));
    LocalMux I__2014 (
            .O(N__22780),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1 ));
    LocalMux I__2013 (
            .O(N__22777),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1 ));
    InMux I__2012 (
            .O(N__22770),
            .I(N__22767));
    LocalMux I__2011 (
            .O(N__22767),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.un2_count_bits_1_0_a2_2 ));
    CascadeMux I__2010 (
            .O(N__22764),
            .I(N__22759));
    CascadeMux I__2009 (
            .O(N__22763),
            .I(N__22756));
    CascadeMux I__2008 (
            .O(N__22762),
            .I(N__22752));
    InMux I__2007 (
            .O(N__22759),
            .I(N__22746));
    InMux I__2006 (
            .O(N__22756),
            .I(N__22746));
    InMux I__2005 (
            .O(N__22755),
            .I(N__22740));
    InMux I__2004 (
            .O(N__22752),
            .I(N__22737));
    InMux I__2003 (
            .O(N__22751),
            .I(N__22734));
    LocalMux I__2002 (
            .O(N__22746),
            .I(N__22731));
    InMux I__2001 (
            .O(N__22745),
            .I(N__22724));
    InMux I__2000 (
            .O(N__22744),
            .I(N__22724));
    InMux I__1999 (
            .O(N__22743),
            .I(N__22724));
    LocalMux I__1998 (
            .O(N__22740),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ));
    LocalMux I__1997 (
            .O(N__22737),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ));
    LocalMux I__1996 (
            .O(N__22734),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ));
    Odrv4 I__1995 (
            .O(N__22731),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ));
    LocalMux I__1994 (
            .O(N__22724),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ));
    InMux I__1993 (
            .O(N__22713),
            .I(N__22707));
    InMux I__1992 (
            .O(N__22712),
            .I(N__22707));
    LocalMux I__1991 (
            .O(N__22707),
            .I(N__22700));
    InMux I__1990 (
            .O(N__22706),
            .I(N__22697));
    InMux I__1989 (
            .O(N__22705),
            .I(N__22690));
    InMux I__1988 (
            .O(N__22704),
            .I(N__22690));
    InMux I__1987 (
            .O(N__22703),
            .I(N__22690));
    Odrv4 I__1986 (
            .O(N__22700),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383 ));
    LocalMux I__1985 (
            .O(N__22697),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383 ));
    LocalMux I__1984 (
            .O(N__22690),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383 ));
    InMux I__1983 (
            .O(N__22683),
            .I(N__22678));
    InMux I__1982 (
            .O(N__22682),
            .I(N__22673));
    InMux I__1981 (
            .O(N__22681),
            .I(N__22673));
    LocalMux I__1980 (
            .O(N__22678),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6 ));
    LocalMux I__1979 (
            .O(N__22673),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6 ));
    CascadeMux I__1978 (
            .O(N__22668),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0_cascade_ ));
    InMux I__1977 (
            .O(N__22665),
            .I(N__22662));
    LocalMux I__1976 (
            .O(N__22662),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_4 ));
    InMux I__1975 (
            .O(N__22659),
            .I(N__22653));
    InMux I__1974 (
            .O(N__22658),
            .I(N__22653));
    LocalMux I__1973 (
            .O(N__22653),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_5 ));
    InMux I__1972 (
            .O(N__22650),
            .I(N__22646));
    InMux I__1971 (
            .O(N__22649),
            .I(N__22643));
    LocalMux I__1970 (
            .O(N__22646),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7 ));
    LocalMux I__1969 (
            .O(N__22643),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7 ));
    InMux I__1968 (
            .O(N__22638),
            .I(N__22632));
    InMux I__1967 (
            .O(N__22637),
            .I(N__22632));
    LocalMux I__1966 (
            .O(N__22632),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_8 ));
    InMux I__1965 (
            .O(N__22629),
            .I(N__22626));
    LocalMux I__1964 (
            .O(N__22626),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_4 ));
    InMux I__1963 (
            .O(N__22623),
            .I(N__22620));
    LocalMux I__1962 (
            .O(N__22620),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_5 ));
    InMux I__1961 (
            .O(N__22617),
            .I(N__22614));
    LocalMux I__1960 (
            .O(N__22614),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_6 ));
    InMux I__1959 (
            .O(N__22611),
            .I(N__22608));
    LocalMux I__1958 (
            .O(N__22608),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_0 ));
    CEMux I__1957 (
            .O(N__22605),
            .I(N__22602));
    LocalMux I__1956 (
            .O(N__22602),
            .I(N__22599));
    Span4Mux_v I__1955 (
            .O(N__22599),
            .I(N__22596));
    Odrv4 I__1954 (
            .O(N__22596),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_i ));
    IoInMux I__1953 (
            .O(N__22593),
            .I(N__22590));
    LocalMux I__1952 (
            .O(N__22590),
            .I(N__22587));
    Span4Mux_s2_v I__1951 (
            .O(N__22587),
            .I(N__22584));
    Span4Mux_v I__1950 (
            .O(N__22584),
            .I(N__22581));
    Span4Mux_v I__1949 (
            .O(N__22581),
            .I(N__22578));
    Odrv4 I__1948 (
            .O(N__22578),
            .I(N_1821_0));
    CascadeMux I__1947 (
            .O(N__22575),
            .I(N__22572));
    InMux I__1946 (
            .O(N__22572),
            .I(N__22569));
    LocalMux I__1945 (
            .O(N__22569),
            .I(N__22566));
    Span12Mux_s8_h I__1944 (
            .O(N__22566),
            .I(N__22563));
    Span12Mux_v I__1943 (
            .O(N__22563),
            .I(N__22560));
    Span12Mux_h I__1942 (
            .O(N__22560),
            .I(N__22557));
    Odrv12 I__1941 (
            .O(N__22557),
            .I(sdin1_c));
    InMux I__1940 (
            .O(N__22554),
            .I(N__22551));
    LocalMux I__1939 (
            .O(N__22551),
            .I(N__22548));
    Span12Mux_h I__1938 (
            .O(N__22548),
            .I(N__22545));
    Span12Mux_v I__1937 (
            .O(N__22545),
            .I(N__22542));
    Span12Mux_h I__1936 (
            .O(N__22542),
            .I(N__22539));
    Odrv12 I__1935 (
            .O(N__22539),
            .I(sdin0_c));
    IoInMux I__1934 (
            .O(N__22536),
            .I(N__22533));
    LocalMux I__1933 (
            .O(N__22533),
            .I(N__22530));
    Span4Mux_s1_h I__1932 (
            .O(N__22530),
            .I(N__22527));
    Sp12to4 I__1931 (
            .O(N__22527),
            .I(N__22524));
    Span12Mux_v I__1930 (
            .O(N__22524),
            .I(N__22521));
    Odrv12 I__1929 (
            .O(N__22521),
            .I(mcu_data_c));
    InMux I__1928 (
            .O(N__22518),
            .I(N__22513));
    InMux I__1927 (
            .O(N__22517),
            .I(N__22510));
    InMux I__1926 (
            .O(N__22516),
            .I(N__22507));
    LocalMux I__1925 (
            .O(N__22513),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0 ));
    LocalMux I__1924 (
            .O(N__22510),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0 ));
    LocalMux I__1923 (
            .O(N__22507),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0 ));
    InMux I__1922 (
            .O(N__22500),
            .I(N__22496));
    InMux I__1921 (
            .O(N__22499),
            .I(N__22493));
    LocalMux I__1920 (
            .O(N__22496),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0 ));
    LocalMux I__1919 (
            .O(N__22493),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0 ));
    InMux I__1918 (
            .O(N__22488),
            .I(N__22482));
    InMux I__1917 (
            .O(N__22487),
            .I(N__22482));
    LocalMux I__1916 (
            .O(N__22482),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370 ));
    CascadeMux I__1915 (
            .O(N__22479),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_cascade_ ));
    InMux I__1914 (
            .O(N__22476),
            .I(N__22471));
    InMux I__1913 (
            .O(N__22475),
            .I(N__22466));
    InMux I__1912 (
            .O(N__22474),
            .I(N__22466));
    LocalMux I__1911 (
            .O(N__22471),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14 ));
    LocalMux I__1910 (
            .O(N__22466),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14 ));
    InMux I__1909 (
            .O(N__22461),
            .I(N__22458));
    LocalMux I__1908 (
            .O(N__22458),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_1 ));
    InMux I__1907 (
            .O(N__22455),
            .I(N__22452));
    LocalMux I__1906 (
            .O(N__22452),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_2 ));
    InMux I__1905 (
            .O(N__22449),
            .I(N__22446));
    LocalMux I__1904 (
            .O(N__22446),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_3 ));
    CascadeMux I__1903 (
            .O(N__22443),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_17_0_cascade_ ));
    InMux I__1902 (
            .O(N__22440),
            .I(N__22437));
    LocalMux I__1901 (
            .O(N__22437),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_12 ));
    CascadeMux I__1900 (
            .O(N__22434),
            .I(N__22430));
    CascadeMux I__1899 (
            .O(N__22433),
            .I(N__22427));
    InMux I__1898 (
            .O(N__22430),
            .I(N__22424));
    InMux I__1897 (
            .O(N__22427),
            .I(N__22421));
    LocalMux I__1896 (
            .O(N__22424),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13 ));
    LocalMux I__1895 (
            .O(N__22421),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13 ));
    InMux I__1894 (
            .O(N__22416),
            .I(N__22405));
    InMux I__1893 (
            .O(N__22415),
            .I(N__22405));
    InMux I__1892 (
            .O(N__22414),
            .I(N__22405));
    InMux I__1891 (
            .O(N__22413),
            .I(N__22400));
    InMux I__1890 (
            .O(N__22412),
            .I(N__22400));
    LocalMux I__1889 (
            .O(N__22405),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0 ));
    LocalMux I__1888 (
            .O(N__22400),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0 ));
    CascadeMux I__1887 (
            .O(N__22395),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0_cascade_ ));
    InMux I__1886 (
            .O(N__22392),
            .I(N__22389));
    LocalMux I__1885 (
            .O(N__22389),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_375 ));
    InMux I__1884 (
            .O(N__22386),
            .I(N__22383));
    LocalMux I__1883 (
            .O(N__22383),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_1 ));
    InMux I__1882 (
            .O(N__22380),
            .I(N__22377));
    LocalMux I__1881 (
            .O(N__22377),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_0 ));
    InMux I__1880 (
            .O(N__22374),
            .I(bfn_5_16_0_));
    InMux I__1879 (
            .O(N__22371),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0 ));
    InMux I__1878 (
            .O(N__22368),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1 ));
    InMux I__1877 (
            .O(N__22365),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2 ));
    InMux I__1876 (
            .O(N__22362),
            .I(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_3 ));
    IoInMux I__1875 (
            .O(N__22359),
            .I(N__22356));
    LocalMux I__1874 (
            .O(N__22356),
            .I(N__22353));
    Span4Mux_s3_h I__1873 (
            .O(N__22353),
            .I(N__22350));
    Span4Mux_v I__1872 (
            .O(N__22350),
            .I(N__22347));
    Odrv4 I__1871 (
            .O(N__22347),
            .I(mcu_sclk_c));
    IoInMux I__1870 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__1869 (
            .O(N__22341),
            .I(N__22338));
    Span12Mux_s5_v I__1868 (
            .O(N__22338),
            .I(N__22335));
    Span12Mux_h I__1867 (
            .O(N__22335),
            .I(N__22332));
    Span12Mux_v I__1866 (
            .O(N__22332),
            .I(N__22329));
    Span12Mux_v I__1865 (
            .O(N__22329),
            .I(N__22326));
    Odrv12 I__1864 (
            .O(N__22326),
            .I(clock_ibuf_gb_io_gb_input));
    INV \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C  (
            .O(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .I(N__47994));
    INV \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C  (
            .O(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .I(N__47993));
    INV \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C  (
            .O(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .I(N__47991));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net ),
            .I(N__65638));
    INV \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C  (
            .O(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ),
            .I(N__47985));
    INV \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C  (
            .O(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net ),
            .I(N__47979));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net ),
            .I(N__65637));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net ),
            .I(N__65612));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net ),
            .I(N__65592));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net ),
            .I(N__65650));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net ),
            .I(N__65636));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net ),
            .I(N__65624));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net ),
            .I(N__65603));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net ),
            .I(N__65635));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net ),
            .I(N__65590));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net ),
            .I(N__65579));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net ),
            .I(N__65621));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net ),
            .I(N__65600));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net ),
            .I(N__65578));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net ),
            .I(N__65543));
    INV \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C  (
            .O(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C_net ),
            .I(N__47981));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net ),
            .I(N__65542));
    INV \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C  (
            .O(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .I(N__47982));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net ),
            .I(N__65563));
    INV \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C  (
            .O(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net ),
            .I(N__47989));
    INV \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C  (
            .O(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net ),
            .I(N__47987));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net ),
            .I(N__65526));
    INV \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C  (
            .O(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net ),
            .I(N__47988));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net ),
            .I(N__65607));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net ),
            .I(N__65540));
    INV \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C  (
            .O(\INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ),
            .I(N__47995));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net ),
            .I(N__65647));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .I(N__65630));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net ),
            .I(N__65620));
    INV \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C  (
            .O(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net ),
            .I(N__47986));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net ),
            .I(N__65574));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net ),
            .I(N__65561));
    INV \INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC  (
            .O(\INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC_net ),
            .I(N__32744));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net ),
            .I(N__65671));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C_net ),
            .I(N__65656));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .I(N__65646));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ),
            .I(N__65629));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net ),
            .I(N__65619));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net ),
            .I(N__65596));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ),
            .I(N__65645));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net ),
            .I(N__65628));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net ),
            .I(N__65655));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .I(N__65644));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net ),
            .I(N__65627));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .I(N__65713));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ),
            .I(N__65693));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .I(N__65654));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .I(N__65643));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ),
            .I(N__65617));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net ),
            .I(N__65735));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net ),
            .I(N__65752));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .I(N__65743));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net ),
            .I(N__65734));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net ),
            .I(N__65723));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net ),
            .I(N__65705));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C_net ),
            .I(N__65664));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ),
            .I(N__65753));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net ),
            .I(N__65751));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ),
            .I(N__65722));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .I(N__65750));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net ),
            .I(N__65741));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net ),
            .I(N__65732));
    INV \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C  (
            .O(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net ),
            .I(N__65749));
    defparam IN_MUX_bfv_18_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_18_0_));
    defparam IN_MUX_bfv_6_18_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_18_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_18_0_));
    defparam IN_MUX_bfv_9_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_19_0_));
    defparam IN_MUX_bfv_20_17_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_17_0_ (
            .carryinitin(),
            .carryinitout(bfn_20_17_0_));
    defparam IN_MUX_bfv_20_18_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_20_18_0_ (
            .carryinitin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7 ),
            .carryinitout(bfn_20_18_0_));
    defparam IN_MUX_bfv_21_27_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_21_27_0_ (
            .carryinitin(),
            .carryinitout(bfn_21_27_0_));
    defparam IN_MUX_bfv_5_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_16_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_19_0_));
    defparam IN_MUX_bfv_6_19_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_19_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_19_0_));
    defparam IN_MUX_bfv_9_22_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_22_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_22_0_));
    defparam IN_MUX_bfv_12_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_20_0_));
    defparam IN_MUX_bfv_18_20_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_20_0_ (
            .carryinitin(),
            .carryinitout(bfn_18_20_0_));
    defparam IN_MUX_bfv_18_21_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_18_21_0_ (
            .carryinitin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_7 ),
            .carryinitout(bfn_18_21_0_));
    defparam IN_MUX_bfv_13_23_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_13_23_0_ (
            .carryinitin(),
            .carryinitout(bfn_13_23_0_));
    ICE_GB clock_ibuf_gb_io_gb (
            .USERSIGNALTOGLOBALBUFFER(N__22344),
            .GLOBALBUFFEROUTPUT(clock_c_g));
    ICE_GB scl_ibuf_RNI7T7F (
            .USERSIGNALTOGLOBALBUFFER(N__51207),
            .GLOBALBUFFEROUTPUT(scl_c_g));
    ICE_GB \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_0_14  (
            .USERSIGNALTOGLOBALBUFFER(N__43296),
            .GLOBALBUFFEROUTPUT(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_g ));
    ICE_GB \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__32250),
            .GLOBALBUFFEROUTPUT(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g ));
    ICE_GB rst_n_ibuf_RNIBNDC_0 (
            .USERSIGNALTOGLOBALBUFFER(N__34806),
            .GLOBALBUFFEROUTPUT(rst_n_c_i_g));
    ICE_GB \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__34818),
            .GLOBALBUFFEROUTPUT(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g ));
    ICE_GB \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__25422),
            .GLOBALBUFFEROUTPUT(\I2C_top_level_inst1.c_state4_0_i_g ));
    ICE_GB IO_PIN_INST_RNIR662 (
            .USERSIGNALTOGLOBALBUFFER(N__57699),
            .GLOBALBUFFEROUTPUT(s_sda_i_g));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIK8VR2_15_LC_4_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIK8VR2_15_LC_4_14_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIK8VR2_15_LC_4_14_7 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIK8VR2_15_LC_4_14_7  (
            .in0(N__23022),
            .in1(N__65767),
            .in2(_gnd_net_),
            .in3(N__22890),
            .lcout(mcu_sclk_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1_LC_4_18_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1_LC_4_18_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1_LC_4_18_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1_LC_4_18_0  (
            .in0(_gnd_net_),
            .in1(N__22380),
            .in2(_gnd_net_),
            .in3(N__30475),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net ),
            .ce(N__23088),
            .sr(N__62944));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_2_LC_4_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_2_LC_4_18_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_2_LC_4_18_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_2_LC_4_18_1  (
            .in0(N__30476),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22386),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net ),
            .ce(N__23088),
            .sr(N__62944));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_0_LC_4_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_0_LC_4_18_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_0_LC_4_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_0_LC_4_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30477),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net ),
            .ce(N__23088),
            .sr(N__62944));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_0_LC_5_16_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_0_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_0_LC_5_16_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_0_LC_5_16_0  (
            .in0(N__22414),
            .in1(N__22518),
            .in2(_gnd_net_),
            .in3(N__22374),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_16_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0 ),
            .clk(N__65721),
            .ce(),
            .sr(N__62950));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_1_LC_5_16_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_1_LC_5_16_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_1_LC_5_16_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_1_LC_5_16_1  (
            .in0(N__22412),
            .in1(N__22788),
            .in2(_gnd_net_),
            .in3(N__22371),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1 ),
            .clk(N__65721),
            .ce(),
            .sr(N__62950));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_2_LC_5_16_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_2_LC_5_16_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_2_LC_5_16_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_2_LC_5_16_2  (
            .in0(N__22415),
            .in1(N__22806),
            .in2(_gnd_net_),
            .in3(N__22368),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2 ),
            .clk(N__65721),
            .ce(),
            .sr(N__62950));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_3_LC_5_16_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_3_LC_5_16_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_3_LC_5_16_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_3_LC_5_16_3  (
            .in0(N__22413),
            .in1(N__22826),
            .in2(_gnd_net_),
            .in3(N__22365),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_3 ),
            .clk(N__65721),
            .ce(),
            .sr(N__62950));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_4_LC_5_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_4_LC_5_16_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_4_LC_5_16_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_4_LC_5_16_4  (
            .in0(N__22416),
            .in1(N__22755),
            .in2(_gnd_net_),
            .in3(N__22362),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65721),
            .ce(),
            .sr(N__62950));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_3_LC_5_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_3_LC_5_16_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_3_LC_5_16_6 .LUT_INIT=16'b1100110000010100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_3_LC_5_16_6  (
            .in0(N__25530),
            .in1(N__22961),
            .in2(N__22941),
            .in3(N__25583),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65721),
            .ce(),
            .sr(N__62950));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13_LC_5_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13_LC_5_17_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13_LC_5_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13_LC_5_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22440),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net ),
            .ce(),
            .sr(N__62945));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m16_LC_5_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m16_LC_5_17_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m16_LC_5_17_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m16_LC_5_17_1  (
            .in0(N__22859),
            .in1(N__22703),
            .in2(_gnd_net_),
            .in3(N__22744),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_17_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_12_LC_5_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_12_LC_5_17_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_12_LC_5_17_2 .LUT_INIT=16'b1111100011111010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_12_LC_5_17_2  (
            .in0(N__23370),
            .in1(N__25629),
            .in2(N__22443),
            .in3(N__23349),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net ),
            .ce(),
            .sr(N__62945));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_14_LC_5_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_14_LC_5_17_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_14_LC_5_17_3 .LUT_INIT=16'b1111001011111010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_14_LC_5_17_3  (
            .in0(N__22475),
            .in1(N__22704),
            .in2(N__22434),
            .in3(N__22745),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net ),
            .ce(),
            .sr(N__62945));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI5JQ51_13_LC_5_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI5JQ51_13_LC_5_17_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI5JQ51_13_LC_5_17_4 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI5JQ51_13_LC_5_17_4  (
            .in0(N__22658),
            .in1(N__22858),
            .in2(N__22433),
            .in3(N__22499),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_6_LC_5_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_6_LC_5_17_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_6_LC_5_17_5 .LUT_INIT=16'b1111111100101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_6_LC_5_17_5  (
            .in0(N__22682),
            .in1(N__22705),
            .in2(N__22762),
            .in3(N__22659),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net ),
            .ce(),
            .sr(N__62945));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI1LAH_14_LC_5_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI1LAH_14_LC_5_17_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI1LAH_14_LC_5_17_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI1LAH_14_LC_5_17_6  (
            .in0(_gnd_net_),
            .in1(N__22474),
            .in2(_gnd_net_),
            .in3(N__22681),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNITF8T1_0_LC_5_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNITF8T1_0_LC_5_17_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNITF8T1_0_LC_5_17_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNITF8T1_0_LC_5_17_7  (
            .in0(N__22517),
            .in1(N__22770),
            .in2(N__22395),
            .in3(N__22743),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_375 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNILFTV2_9_LC_5_18_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNILFTV2_9_LC_5_18_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNILFTV2_9_LC_5_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNILFTV2_9_LC_5_18_0  (
            .in0(N__25075),
            .in1(N__22487),
            .in2(N__25696),
            .in3(N__22392),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10_LC_5_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10_LC_5_18_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10_LC_5_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10_LC_5_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25076),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net ),
            .ce(),
            .sr(N__62939));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_11_LC_5_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_11_LC_5_18_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_11_LC_5_18_2 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_11_LC_5_18_2  (
            .in0(N__22713),
            .in1(N__22857),
            .in2(N__22763),
            .in3(N__22488),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net ),
            .ce(),
            .sr(N__62939));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_en_count_data_i_LC_5_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_en_count_data_i_LC_5_18_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_en_count_data_i_LC_5_18_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_en_count_data_i_LC_5_18_3  (
            .in0(N__22856),
            .in1(N__25686),
            .in2(N__25751),
            .in3(N__25074),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_11_LC_5_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_11_LC_5_18_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_11_LC_5_18_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_11_LC_5_18_4  (
            .in0(_gnd_net_),
            .in1(N__25736),
            .in2(_gnd_net_),
            .in3(N__22855),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_0_11_LC_5_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_0_11_LC_5_18_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_0_11_LC_5_18_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_0_11_LC_5_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22479),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_15_LC_5_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_15_LC_5_18_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_15_LC_5_18_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_15_LC_5_18_6  (
            .in0(N__22712),
            .in1(_gnd_net_),
            .in2(N__22764),
            .in3(N__22476),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net ),
            .ce(),
            .sr(N__62939));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1_LC_5_19_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1_LC_5_19_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1_LC_5_19_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1_LC_5_19_0  (
            .in0(_gnd_net_),
            .in1(N__25740),
            .in2(_gnd_net_),
            .in3(N__22611),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_2_LC_5_19_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_2_LC_5_19_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_2_LC_5_19_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_2_LC_5_19_1  (
            .in0(N__25741),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22461),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_3_LC_5_19_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_3_LC_5_19_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_3_LC_5_19_2 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_3_LC_5_19_2  (
            .in0(_gnd_net_),
            .in1(N__25742),
            .in2(_gnd_net_),
            .in3(N__22455),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_4_LC_5_19_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_4_LC_5_19_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_4_LC_5_19_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_4_LC_5_19_3  (
            .in0(N__25743),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22449),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_5_LC_5_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_5_LC_5_19_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_5_LC_5_19_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_5_LC_5_19_4  (
            .in0(_gnd_net_),
            .in1(N__25744),
            .in2(_gnd_net_),
            .in3(N__22629),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_6_LC_5_19_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_6_LC_5_19_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_6_LC_5_19_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_6_LC_5_19_5  (
            .in0(N__25745),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22623),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_7_LC_5_19_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_7_LC_5_19_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_7_LC_5_19_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_7_LC_5_19_6  (
            .in0(_gnd_net_),
            .in1(N__25746),
            .in2(_gnd_net_),
            .in3(N__22617),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_read ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_0_LC_5_19_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_0_LC_5_19_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_0_LC_5_19_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_0_LC_5_19_7  (
            .in0(N__25747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net ),
            .ce(N__22605),
            .sr(N__62929));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNI8PPB5_0_LC_5_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNI8PPB5_0_LC_5_22_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNI8PPB5_0_LC_5_22_2 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNI8PPB5_0_LC_5_22_2  (
            .in0(N__65769),
            .in1(N__23211),
            .in2(N__23034),
            .in3(N__27210),
            .lcout(N_1821_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIBD7Q2_15_LC_6_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIBD7Q2_15_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIBD7Q2_15_LC_6_15_0 .LUT_INIT=16'b0110001001000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIBD7Q2_15_LC_6_15_0  (
            .in0(N__22883),
            .in1(N__23015),
            .in2(N__22575),
            .in3(N__22554),
            .lcout(mcu_data_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNIEJ431_0_LC_6_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNIEJ431_0_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNIEJ431_0_LC_6_16_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNIEJ431_0_LC_6_16_0  (
            .in0(N__22804),
            .in1(N__22786),
            .in2(N__22827),
            .in3(N__22516),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m33_e_LC_6_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m33_e_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m33_e_LC_6_16_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m33_e_LC_6_16_2  (
            .in0(N__23288),
            .in1(N__22650),
            .in2(_gnd_net_),
            .in3(N__22500),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93_0_LC_6_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93_0_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93_0_LC_6_16_3 .LUT_INIT=16'b1011111110110101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93_0_LC_6_16_3  (
            .in0(N__27568),
            .in1(N__27678),
            .in2(N__29970),
            .in3(N__28863),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIA8O66_0_LC_6_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIA8O66_0_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIA8O66_0_LC_6_16_4 .LUT_INIT=16'b0000100001001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIA8O66_0_LC_6_16_4  (
            .in0(N__25695),
            .in1(N__65768),
            .in2(N__22902),
            .in3(N__22833),
            .lcout(sclk1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32_0_LC_6_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32_0_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32_0_LC_6_16_5 .LUT_INIT=16'b0101111111011111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32_0_LC_6_16_5  (
            .in0(N__27567),
            .in1(N__22882),
            .in2(N__29969),
            .in3(N__22866),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNI4GBQ_1_LC_6_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNI4GBQ_1_LC_6_17_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNI4GBQ_1_LC_6_17_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNI4GBQ_1_LC_6_17_1  (
            .in0(N__22825),
            .in1(N__22805),
            .in2(_gnd_net_),
            .in3(N__22787),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.un2_count_bits_1_0_a2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7_LC_6_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7_LC_6_17_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7_LC_6_17_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7_LC_6_17_2  (
            .in0(N__22751),
            .in1(N__22706),
            .in2(_gnd_net_),
            .in3(N__22683),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ),
            .ce(),
            .sr(N__62940));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_4_LC_6_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_4_LC_6_17_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_4_LC_6_17_3 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_4_LC_6_17_3  (
            .in0(N__22637),
            .in1(N__25627),
            .in2(_gnd_net_),
            .in3(N__23347),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ),
            .ce(),
            .sr(N__62940));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_RNIICQD1_4_LC_6_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_RNIICQD1_4_LC_6_17_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_RNIICQD1_4_LC_6_17_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_RNIICQD1_4_LC_6_17_4  (
            .in0(N__22957),
            .in1(N__23621),
            .in2(N__25491),
            .in3(N__22922),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_9_LC_6_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_9_LC_6_17_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_9_LC_6_17_5 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_9_LC_6_17_5  (
            .in0(N__22638),
            .in1(_gnd_net_),
            .in2(N__22668),
            .in3(N__25628),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ),
            .ce(),
            .sr(N__62940));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_5_LC_6_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_5_LC_6_17_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_5_LC_6_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_5_LC_6_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22665),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ),
            .ce(),
            .sr(N__62940));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_8_LC_6_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_8_LC_6_17_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_8_LC_6_17_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_8_LC_6_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22649),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net ),
            .ce(),
            .sr(N__62940));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_c_0_LC_6_18_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_c_0_LC_6_18_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_c_0_LC_6_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_c_0_LC_6_18_0  (
            .in0(_gnd_net_),
            .in1(N__25617),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_18_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_6_18_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_6_18_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_6_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_6_18_1  (
            .in0(_gnd_net_),
            .in1(N__25487),
            .in2(_gnd_net_),
            .in3(N__22968),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_6_18_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_6_18_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_6_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_6_18_2  (
            .in0(_gnd_net_),
            .in1(N__23625),
            .in2(_gnd_net_),
            .in3(N__22965),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_6_18_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_6_18_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_6_18_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_6_18_3  (
            .in0(_gnd_net_),
            .in1(N__22962),
            .in2(_gnd_net_),
            .in3(N__22929),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_4_LC_6_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_4_LC_6_18_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_4_LC_6_18_4 .LUT_INIT=16'b1000100110001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_4_LC_6_18_4  (
            .in0(N__25577),
            .in1(N__22923),
            .in2(N__25535),
            .in3(N__22926),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65733),
            .ce(),
            .sr(N__62930));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_0_LC_6_19_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_0_LC_6_19_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_0_LC_6_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_0_LC_6_19_0  (
            .in0(N__22987),
            .in1(N__23508),
            .in2(_gnd_net_),
            .in3(N__22911),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_6_19_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0 ),
            .clk(N__65742),
            .ce(),
            .sr(N__62920));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_1_LC_6_19_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_1_LC_6_19_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_1_LC_6_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_1_LC_6_19_1  (
            .in0(N__22985),
            .in1(N__23547),
            .in2(_gnd_net_),
            .in3(N__22908),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1 ),
            .clk(N__65742),
            .ce(),
            .sr(N__62920));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_2_LC_6_19_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_2_LC_6_19_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_2_LC_6_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_2_LC_6_19_2  (
            .in0(N__22988),
            .in1(N__23565),
            .in2(_gnd_net_),
            .in3(N__22905),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2 ),
            .clk(N__65742),
            .ce(),
            .sr(N__62920));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_3_LC_6_19_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_3_LC_6_19_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_3_LC_6_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_3_LC_6_19_3  (
            .in0(N__22986),
            .in1(N__23528),
            .in2(_gnd_net_),
            .in3(N__23040),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_3 ),
            .clk(N__65742),
            .ce(),
            .sr(N__62920));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_4_LC_6_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_4_LC_6_19_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_4_LC_6_19_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_4_LC_6_19_4  (
            .in0(N__22989),
            .in1(N__23450),
            .in2(_gnd_net_),
            .in3(N__23037),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65742),
            .ce(),
            .sr(N__62920));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIMOE52_15_LC_6_20_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIMOE52_15_LC_6_20_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIMOE52_15_LC_6_20_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIMOE52_15_LC_6_20_1  (
            .in0(N__23385),
            .in1(N__23591),
            .in2(N__23001),
            .in3(N__26994),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_333 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI02AE1_15_LC_6_20_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI02AE1_15_LC_6_20_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI02AE1_15_LC_6_20_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI02AE1_15_LC_6_20_2  (
            .in0(N__25804),
            .in1(N__23384),
            .in2(N__23592),
            .in3(N__25839),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_376 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_sck_m8_i_a2_1_LC_6_20_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_sck_m8_i_a2_1_LC_6_20_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_sck_m8_i_a2_1_LC_6_20_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_sck_m8_i_a2_1_LC_6_20_3  (
            .in0(N__25838),
            .in1(N__26923),
            .in2(_gnd_net_),
            .in3(N__25802),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI0EFP1_13_LC_6_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI0EFP1_13_LC_6_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI0EFP1_13_LC_6_20_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI0EFP1_13_LC_6_20_4  (
            .in0(_gnd_net_),
            .in1(N__23573),
            .in2(N__22992),
            .in3(N__23309),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6_LC_6_20_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6_LC_6_20_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6_LC_6_20_5 .LUT_INIT=16'b1111011111110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6_LC_6_20_5  (
            .in0(N__23405),
            .in1(N__23449),
            .in2(N__23313),
            .in3(N__25803),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net ),
            .ce(),
            .sr(N__62912));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_14_LC_6_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_14_LC_6_20_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_14_LC_6_20_6 .LUT_INIT=16'b1111111101110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_14_LC_6_20_6  (
            .in0(N__23448),
            .in1(N__23404),
            .in2(N__25845),
            .in3(N__23574),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net ),
            .ce(),
            .sr(N__62912));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_11_LC_6_20_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_11_LC_6_20_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_11_LC_6_20_7 .LUT_INIT=16'b1111010111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_11_LC_6_20_7  (
            .in0(N__23406),
            .in1(N__30472),
            .in2(N__23451),
            .in3(N__26924),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net ),
            .ce(),
            .sr(N__62912));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7_LC_6_21_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7_LC_6_21_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7_LC_6_21_0 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7_LC_6_21_0  (
            .in0(_gnd_net_),
            .in1(N__23124),
            .in2(_gnd_net_),
            .in3(N__30463),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.dout_read ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ),
            .ce(N__23087),
            .sr(N__62901));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_RNINM921_23_LC_6_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_RNINM921_23_LC_6_21_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_RNINM921_23_LC_6_21_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_RNINM921_23_LC_6_21_1  (
            .in0(N__32633),
            .in1(N__26124),
            .in2(_gnd_net_),
            .in3(N__49560),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_237_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_RNIU7DV3_7_LC_6_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_RNIU7DV3_7_LC_6_21_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_RNIU7DV3_7_LC_6_21_2 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_RNIU7DV3_7_LC_6_21_2  (
            .in0(N__26982),
            .in1(N__23148),
            .in2(N__23142),
            .in3(N__23046),
            .lcout(N_85_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_6_LC_6_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_6_LC_6_21_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_6_LC_6_21_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_6_LC_6_21_3  (
            .in0(N__30462),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23118),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ),
            .ce(N__23087),
            .sr(N__62901));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_5_LC_6_21_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_5_LC_6_21_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_5_LC_6_21_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_5_LC_6_21_4  (
            .in0(_gnd_net_),
            .in1(N__23112),
            .in2(_gnd_net_),
            .in3(N__30461),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ),
            .ce(N__23087),
            .sr(N__62901));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_4_LC_6_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_4_LC_6_21_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_4_LC_6_21_5 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_4_LC_6_21_5  (
            .in0(N__30460),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23094),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ),
            .ce(N__23087),
            .sr(N__62901));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI7VAM_11_LC_6_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI7VAM_11_LC_6_21_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI7VAM_11_LC_6_21_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI7VAM_11_LC_6_21_6  (
            .in0(_gnd_net_),
            .in1(N__30458),
            .in2(_gnd_net_),
            .in3(N__26932),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_370_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_3_LC_6_21_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_3_LC_6_21_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_3_LC_6_21_7 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_3_LC_6_21_7  (
            .in0(N__30459),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23106),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net ),
            .ce(N__23087),
            .sr(N__62901));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNISO0C4_0_LC_6_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNISO0C4_0_LC_6_22_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNISO0C4_0_LC_6_22_1 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNISO0C4_0_LC_6_22_1  (
            .in0(N__25869),
            .in1(N__32635),
            .in2(N__23754),
            .in3(N__26997),
            .lcout(N_1820_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIS2262_0_LC_6_22_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIS2262_0_LC_6_22_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIS2262_0_LC_6_22_5 .LUT_INIT=16'b1100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIS2262_0_LC_6_22_5  (
            .in0(N__27195),
            .in1(N__23220),
            .in2(N__32640),
            .in3(N__26999),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_u_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIPJA61_0_LC_6_22_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIPJA61_0_LC_6_22_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIPJA61_0_LC_6_22_6 .LUT_INIT=16'b1010110100001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIPJA61_0_LC_6_22_6  (
            .in0(N__26998),
            .in1(N__27194),
            .in2(N__27150),
            .in3(N__32636),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNID2OK2_0_LC_6_22_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNID2OK2_0_LC_6_22_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNID2OK2_0_LC_6_22_7 .LUT_INIT=16'b1100000011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNID2OK2_0_LC_6_22_7  (
            .in0(_gnd_net_),
            .in1(N__32634),
            .in2(N__23214),
            .in3(N__31098),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.sclk_u_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_7_LC_7_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_7_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_7_LC_7_12_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_7_LC_7_12_0  (
            .in0(N__53314),
            .in1(N__40529),
            .in2(N__38319),
            .in3(N__41058),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_7_LC_7_12_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_7_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_7_LC_7_12_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_7_LC_7_12_1  (
            .in0(N__23205),
            .in1(N__52781),
            .in2(N__23190),
            .in3(N__52522),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_7_LC_7_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_7_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_7_LC_7_12_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_7_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__52236),
            .in2(N__23172),
            .in3(N__40551),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_7_LC_7_12_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_7_LC_7_12_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_7_LC_7_12_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_7_LC_7_12_3  (
            .in0(N__23169),
            .in1(N__33456),
            .in2(N__23157),
            .in3(N__23154),
            .lcout(I2C_top_level_inst1_s_data_oreg_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65639),
            .ce(N__54525),
            .sr(N__64964));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_7_LC_7_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_7_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_7_LC_7_12_4 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_7_LC_7_12_4  (
            .in0(N__51927),
            .in1(N__25014),
            .in2(N__24855),
            .in3(N__48759),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4_LC_7_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4_LC_7_14_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4_LC_7_14_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__28999),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C_net ),
            .ce(),
            .sr(N__62951));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_5_LC_7_15_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_5_LC_7_15_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_5_LC_7_15_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_5_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41806),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65679),
            .ce(N__44092),
            .sr(N__64963));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_7_LC_7_15_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_7_LC_7_15_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_7_LC_7_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_7_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41689),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65679),
            .ce(N__44092),
            .sr(N__64963));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16_LC_7_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16_LC_7_17_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16_LC_7_17_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16_LC_7_17_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23289),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62931));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_LC_7_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_LC_7_17_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_LC_7_17_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_LC_7_17_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23226),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62931));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18_LC_7_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18_LC_7_18_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18_LC_7_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18_LC_7_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29049),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net ),
            .ce(),
            .sr(N__62921));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1_23_LC_7_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1_23_LC_7_18_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1_23_LC_7_18_2 .LUT_INIT=16'b0000101011000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1_23_LC_7_18_2  (
            .in0(N__36129),
            .in1(N__26802),
            .in2(N__29968),
            .in3(N__27579),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1Z0Z_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNIUP1S2_23_LC_7_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNIUP1S2_23_LC_7_18_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNIUP1S2_23_LC_7_18_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNIUP1S2_23_LC_7_18_3  (
            .in0(N__23232),
            .in1(_gnd_net_),
            .in2(N__23268),
            .in3(N__25682),
            .lcout(N_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01_0_LC_7_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01_0_LC_7_18_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01_0_LC_7_18_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01_0_LC_7_18_4  (
            .in0(N__29958),
            .in1(N__27578),
            .in2(_gnd_net_),
            .in3(N__23244),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHF2R_0_LC_7_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHF2R_0_LC_7_18_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHF2R_0_LC_7_18_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHF2R_0_LC_7_18_5  (
            .in0(_gnd_net_),
            .in1(N__29957),
            .in2(_gnd_net_),
            .in3(N__35860),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_reti_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_1_LC_7_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_1_LC_7_18_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_1_LC_7_18_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_1_LC_7_18_6  (
            .in0(N__35861),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37173),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1867_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_0_LC_7_18_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_0_LC_7_18_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_0_LC_7_18_7 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_0_LC_7_18_7  (
            .in0(N__25626),
            .in1(N__25681),
            .in2(N__23366),
            .in3(N__23348),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net ),
            .ce(),
            .sr(N__62921));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIN9BU_0_LC_7_19_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIN9BU_0_LC_7_19_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIN9BU_0_LC_7_19_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIN9BU_0_LC_7_19_0  (
            .in0(N__23442),
            .in1(N__23546),
            .in2(N__23331),
            .in3(N__23507),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNINH4C_2_LC_7_19_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNINH4C_2_LC_7_19_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNINH4C_2_LC_7_19_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNINH4C_2_LC_7_19_1  (
            .in0(_gnd_net_),
            .in1(N__23527),
            .in2(_gnd_net_),
            .in3(N__23564),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_RNIEOU21_4_LC_7_19_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_RNIEOU21_4_LC_7_19_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_RNIEOU21_4_LC_7_19_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_RNIEOU21_4_LC_7_19_2  (
            .in0(N__25926),
            .in1(N__25962),
            .in2(N__25887),
            .in3(N__25995),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4_LC_7_19_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4_LC_7_19_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4_LC_7_19_3 .LUT_INIT=16'b0000110011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4_LC_7_19_3  (
            .in0(_gnd_net_),
            .in1(N__23297),
            .in2(N__23322),
            .in3(N__25458),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net ),
            .ce(),
            .sr(N__62913));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_9_LC_7_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_9_LC_7_19_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_9_LC_7_19_4 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_9_LC_7_19_4  (
            .in0(N__25459),
            .in1(_gnd_net_),
            .in2(N__23301),
            .in3(N__23485),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net ),
            .ce(),
            .sr(N__62913));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_5_LC_7_19_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_5_LC_7_19_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_5_LC_7_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_5_LC_7_19_5  (
            .in0(N__23319),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net ),
            .ce(),
            .sr(N__62913));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_8_LC_7_19_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_8_LC_7_19_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_8_LC_7_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_8_LC_7_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23383),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net ),
            .ce(),
            .sr(N__62913));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16_LC_7_20_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16_LC_7_20_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16_LC_7_20_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16_LC_7_20_0  (
            .in0(_gnd_net_),
            .in1(N__23587),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62902));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_15_LC_7_20_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_15_LC_7_20_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_15_LC_7_20_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_15_LC_7_20_1  (
            .in0(N__23446),
            .in1(N__23402),
            .in2(_gnd_net_),
            .in3(N__25840),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62902));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_13_LC_7_20_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_13_LC_7_20_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_13_LC_7_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_13_LC_7_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23457),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62902));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_0_LC_7_20_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_0_LC_7_20_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_0_LC_7_20_3 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_0_LC_7_20_3  (
            .in0(N__25460),
            .in1(N__23486),
            .in2(N__23472),
            .in3(N__26976),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62902));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIAV8O_0_LC_7_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIAV8O_0_LC_7_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIAV8O_0_LC_7_20_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIAV8O_0_LC_7_20_4  (
            .in0(N__23563),
            .in1(N__23545),
            .in2(N__23529),
            .in3(N__23506),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNO_0_12_LC_7_20_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNO_0_12_LC_7_20_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNO_0_12_LC_7_20_5 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNO_0_12_LC_7_20_5  (
            .in0(_gnd_net_),
            .in1(N__23441),
            .in2(N__23490),
            .in3(N__26931),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_369_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_12_LC_7_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_12_LC_7_20_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_12_LC_7_20_6 .LUT_INIT=16'b1111110011110100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_12_LC_7_20_6  (
            .in0(N__23487),
            .in1(N__23471),
            .in2(N__23460),
            .in3(N__25461),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62902));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_7_LC_7_20_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_7_LC_7_20_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_7_LC_7_20_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_7_LC_7_20_7  (
            .in0(N__23447),
            .in1(N__23403),
            .in2(_gnd_net_),
            .in3(N__25808),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net ),
            .ce(),
            .sr(N__62902));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0_LC_7_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0_LC_7_21_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0_LC_7_21_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0_LC_7_21_1  (
            .in0(N__26013),
            .in1(N__26061),
            .in2(_gnd_net_),
            .in3(N__23745),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net ),
            .ce(),
            .sr(N__62889));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_1_LC_7_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_1_LC_7_21_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_1_LC_7_21_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_1_LC_7_21_6  (
            .in0(_gnd_net_),
            .in1(N__27193),
            .in2(_gnd_net_),
            .in3(N__27107),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net ),
            .ce(),
            .sr(N__62889));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI9R351_9_LC_7_22_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI9R351_9_LC_7_22_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI9R351_9_LC_7_22_0 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI9R351_9_LC_7_22_0  (
            .in0(N__30514),
            .in1(N__32632),
            .in2(_gnd_net_),
            .in3(N__26996),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.csb_u_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNINIFT1_0_LC_7_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNINIFT1_0_LC_7_22_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNINIFT1_0_LC_7_22_1 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNINIFT1_0_LC_7_22_1  (
            .in0(N__30473),
            .in1(N__27183),
            .in2(N__23760),
            .in3(N__27069),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_331_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIG6Q33_0_LC_7_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIG6Q33_0_LC_7_22_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIG6Q33_0_LC_7_22_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIG6Q33_0_LC_7_22_2  (
            .in0(N__27035),
            .in1(N__32631),
            .in2(N__23757),
            .in3(N__26995),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_LC_7_22_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_LC_7_22_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_LC_7_22_3 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_LC_7_22_3  (
            .in0(_gnd_net_),
            .in1(N__27182),
            .in2(_gnd_net_),
            .in3(N__27068),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_391_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_ns_1_0__m7_0_a2_3_LC_7_22_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_ns_1_0__m7_0_a2_3_LC_7_22_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_ns_1_0__m7_0_a2_3_LC_7_22_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_ns_1_0__m7_0_a2_3_LC_7_22_6  (
            .in0(N__26079),
            .in1(N__26097),
            .in2(N__27036),
            .in3(N__26115),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.m7_0_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec0_0_a2_i_LC_9_2_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec0_0_a2_i_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec0_0_a2_i_LC_9_2_3 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec0_0_a2_i_LC_9_2_3  (
            .in0(N__38919),
            .in1(N__38823),
            .in2(_gnd_net_),
            .in3(N__26673),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_0_LC_9_6_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_0_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_0_LC_9_6_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_0_LC_9_6_4  (
            .in0(N__61964),
            .in1(N__26336),
            .in2(_gnd_net_),
            .in3(N__50387),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_1_LC_9_6_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_1_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_1_LC_9_6_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_1_LC_9_6_6  (
            .in0(N__61820),
            .in1(N__26337),
            .in2(_gnd_net_),
            .in3(N__50388),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_2_LC_9_7_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_2_LC_9_7_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_2_LC_9_7_0 .LUT_INIT=16'b1100110000010100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_2_LC_9_7_0  (
            .in0(N__25536),
            .in1(N__23606),
            .in2(N__23646),
            .in3(N__25590),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65555),
            .ce(),
            .sr(N__62961));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_12_LC_9_7_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_12_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_12_LC_9_7_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_12_LC_9_7_3  (
            .in0(N__58561),
            .in1(N__26288),
            .in2(_gnd_net_),
            .in3(N__50405),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_13_LC_9_7_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_13_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_13_LC_9_7_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_13_LC_9_7_4  (
            .in0(N__50403),
            .in1(_gnd_net_),
            .in2(N__26330),
            .in3(N__58332),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_459_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_14_LC_9_7_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_14_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_14_LC_9_7_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_14_LC_9_7_5  (
            .in0(N__58455),
            .in1(N__26292),
            .in2(_gnd_net_),
            .in3(N__50406),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_15_LC_9_7_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_15_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_15_LC_9_7_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_15_LC_9_7_6  (
            .in0(N__50404),
            .in1(_gnd_net_),
            .in2(N__26331),
            .in3(N__57509),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_16_LC_9_7_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_16_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_16_LC_9_7_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_16_LC_9_7_7  (
            .in0(N__57636),
            .in1(N__26296),
            .in2(_gnd_net_),
            .in3(N__50402),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_8_LC_9_8_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_8_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_8_LC_9_8_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_8_LC_9_8_0  (
            .in0(N__61963),
            .in1(N__23847),
            .in2(N__44665),
            .in3(N__38372),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_20_LC_9_8_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_20_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_20_LC_9_8_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_20_LC_9_8_1  (
            .in0(N__61545),
            .in1(N__26264),
            .in2(_gnd_net_),
            .in3(N__50390),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_o3_0_LC_9_8_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_o3_0_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_o3_0_LC_9_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_o3_0_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__59554),
            .in2(_gnd_net_),
            .in3(N__50456),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_3_LC_9_8_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_3_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_3_LC_9_8_3 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_3_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__63909),
            .in2(N__23802),
            .in3(N__50391),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_466_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_4_LC_9_8_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_4_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_4_LC_9_8_4 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_4_LC_9_8_4  (
            .in0(N__50393),
            .in1(_gnd_net_),
            .in2(N__26325),
            .in3(N__63799),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_5_LC_9_8_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_5_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_5_LC_9_8_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_5_LC_9_8_5  (
            .in0(N__63661),
            .in1(N__26271),
            .in2(_gnd_net_),
            .in3(N__50394),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_22_LC_9_8_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_22_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_22_LC_9_8_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_22_LC_9_8_6  (
            .in0(N__50389),
            .in1(_gnd_net_),
            .in2(N__26324),
            .in3(N__61310),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_9_LC_9_8_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_9_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_9_LC_9_8_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_9_LC_9_8_7  (
            .in0(N__46501),
            .in1(N__26263),
            .in2(_gnd_net_),
            .in3(N__50392),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_25_LC_9_9_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_25_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_25_LC_9_9_0 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_25_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__50348),
            .in2(N__26326),
            .in3(N__61014),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_23_LC_9_9_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_23_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_23_LC_9_9_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_23_LC_9_9_1  (
            .in0(N__61246),
            .in1(N__26277),
            .in2(_gnd_net_),
            .in3(N__50352),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_26_LC_9_9_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_26_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_26_LC_9_9_2 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_26_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__50347),
            .in2(N__26327),
            .in3(N__60912),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_448_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_21_LC_9_9_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_21_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_21_LC_9_9_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_21_LC_9_9_3  (
            .in0(N__50351),
            .in1(N__26276),
            .in2(_gnd_net_),
            .in3(N__61449),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_29_LC_9_9_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_29_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_29_LC_9_9_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_29_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__50350),
            .in2(N__26328),
            .in3(N__62265),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_10_LC_9_9_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_10_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_10_LC_9_9_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_10_LC_9_9_5  (
            .in0(N__58749),
            .in1(N__26272),
            .in2(_gnd_net_),
            .in3(N__50353),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_30_LC_9_9_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_30_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_30_LC_9_9_6 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_30_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__50349),
            .in2(N__26329),
            .in3(N__62132),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_2_LC_9_9_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_2_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_2_LC_9_9_7 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_2_LC_9_9_7  (
            .in0(N__61730),
            .in1(N__26284),
            .in2(_gnd_net_),
            .in3(N__50354),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_24_LC_9_10_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_24_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_24_LC_9_10_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_24_LC_9_10_0  (
            .in0(N__61126),
            .in1(N__50407),
            .in2(_gnd_net_),
            .in3(N__26332),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_LC_9_10_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_LC_9_10_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_LC_9_10_1  (
            .in0(N__38912),
            .in1(N__38806),
            .in2(_gnd_net_),
            .in3(N__26665),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1826_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_27_LC_9_10_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_27_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_27_LC_9_10_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_27_LC_9_10_2  (
            .in0(N__60805),
            .in1(N__50408),
            .in2(_gnd_net_),
            .in3(N__26333),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_11_LC_9_11_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_11_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_11_LC_9_11_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_11_LC_9_11_4  (
            .in0(N__58666),
            .in1(N__26334),
            .in2(_gnd_net_),
            .in3(N__50380),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_28_LC_9_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_28_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_28_LC_9_11_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_28_LC_9_11_6  (
            .in0(N__62337),
            .in1(N__26335),
            .in2(_gnd_net_),
            .in3(N__50379),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_5_LC_9_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_5_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_5_LC_9_12_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_5_LC_9_12_0  (
            .in0(N__24417),
            .in1(N__44616),
            .in2(N__24408),
            .in3(N__44372),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_6_LC_9_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_6_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_6_LC_9_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_6_LC_9_12_2  (
            .in0(N__25059),
            .in1(N__44614),
            .in2(N__25050),
            .in3(N__44370),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_6_LC_9_12_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_6_LC_9_12_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_6_LC_9_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_6_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41757),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65616),
            .ce(N__44106),
            .sr(N__64966));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_7_LC_9_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_7_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_7_LC_9_12_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_7_LC_9_12_4  (
            .in0(N__25041),
            .in1(N__44615),
            .in2(N__25032),
            .in3(N__44371),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNI7VNRE_LC_9_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNI7VNRE_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNI7VNRE_LC_9_14_0 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNI7VNRE_LC_9_14_0  (
            .in0(N__64259),
            .in1(N__38994),
            .in2(_gnd_net_),
            .in3(N__39015),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec3_0_a2_i_LC_9_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec3_0_a2_i_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec3_0_a2_i_LC_9_14_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec3_0_a2_i_LC_9_14_5  (
            .in0(N__38905),
            .in1(N__38822),
            .in2(_gnd_net_),
            .in3(N__26672),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1827_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_7_LC_9_14_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_7_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_7_LC_9_14_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_7_LC_9_14_7  (
            .in0(N__43570),
            .in1(N__37873),
            .in2(N__24873),
            .in3(N__64260),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_863 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.electr_config_test_1_LC_9_15_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.electr_config_test_1_LC_9_15_1 .SEQ_MODE=4'b1000;
    defparam \serializer_mod_inst.electr_config_test_1_LC_9_15_1 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \serializer_mod_inst.electr_config_test_1_LC_9_15_1  (
            .in0(N__24818),
            .in1(N__45486),
            .in2(N__35487),
            .in3(N__45087),
            .lcout(s1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65652),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_c_RNIA3PRE_LC_9_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_c_RNIA3PRE_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_c_RNIA3PRE_LC_9_15_3 .LUT_INIT=16'b1000100000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_c_RNIA3PRE_LC_9_15_3  (
            .in0(N__64261),
            .in1(N__38949),
            .in2(_gnd_net_),
            .in3(N__38973),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNO_LC_9_15_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNO_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNO_LC_9_15_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNO_LC_9_15_5  (
            .in0(N__35482),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50746),
            .lcout(\I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_LC_9_15_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_LC_9_15_6 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_LC_9_15_6  (
            .in0(N__50747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35483),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_1_LC_9_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_1_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_1_LC_9_16_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_1_LC_9_16_0  (
            .in0(N__40602),
            .in1(N__33654),
            .in2(_gnd_net_),
            .in3(N__36235),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_597 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_LC_9_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_LC_9_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_LC_9_16_1  (
            .in0(N__36236),
            .in1(N__25395),
            .in2(_gnd_net_),
            .in3(N__30969),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_596_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_0_LC_9_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_0_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_0_LC_9_16_2 .LUT_INIT=16'b1110110010101000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_0_LC_9_16_2  (
            .in0(N__35973),
            .in1(N__29855),
            .in2(N__25404),
            .in3(N__25401),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_id_prdata_1_4_u_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_26_LC_9_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_26_LC_9_16_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_26_LC_9_16_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_26_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__60901),
            .in2(_gnd_net_),
            .in3(N__59381),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_oZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65667),
            .ce(N__54119),
            .sr(N__62922));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIRLAS1_2_LC_9_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIRLAS1_2_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIRLAS1_2_LC_9_16_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIRLAS1_2_LC_9_16_4  (
            .in0(N__39621),
            .in1(N__46911),
            .in2(_gnd_net_),
            .in3(N__39141),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_1615 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_1615_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_2_LC_9_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_2_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_2_LC_9_16_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_2_LC_9_16_5  (
            .in0(N__64229),
            .in1(_gnd_net_),
            .in2(N__25389),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_0_LC_9_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_0_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_0_LC_9_16_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_0_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__64228),
            .in2(_gnd_net_),
            .in3(N__36237),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_3_LC_9_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_3_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_3_LC_9_16_7 .LUT_INIT=16'b0010011100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_3_LC_9_16_7  (
            .in0(N__39142),
            .in1(N__39576),
            .in2(N__54351),
            .in3(N__64230),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIP15Q1_9_LC_9_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIP15Q1_9_LC_9_17_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIP15Q1_9_LC_9_17_3 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIP15Q1_9_LC_9_17_3  (
            .in0(N__29951),
            .in1(N__27572),
            .in2(N__25701),
            .in3(N__25080),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.csb_u_i_a2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIGVSD3_0_LC_9_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIGVSD3_0_LC_9_17_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIGVSD3_0_LC_9_17_4 .LUT_INIT=16'b0010001110101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIGVSD3_0_LC_9_17_4  (
            .in0(N__25755),
            .in1(N__25635),
            .in2(N__25704),
            .in3(N__25697),
            .lcout(N_1822_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_RNI0JD21_LC_9_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_RNI0JD21_LC_9_17_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_RNI0JD21_LC_9_17_6 .LUT_INIT=16'b0011000000000010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_RNI0JD21_LC_9_17_6  (
            .in0(N__30243),
            .in1(N__27831),
            .in2(N__27798),
            .in3(N__29950),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.csb_u_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_1_LC_9_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_1_LC_9_18_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_1_LC_9_18_2 .LUT_INIT=16'b1010101100000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_1_LC_9_18_2  (
            .in0(N__25778),
            .in1(N__25971),
            .in2(N__26895),
            .in3(N__25991),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65691),
            .ce(),
            .sr(N__62903));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_2_LC_9_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_2_LC_9_18_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_2_LC_9_18_3 .LUT_INIT=16'b1100110000010100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_2_LC_9_18_3  (
            .in0(N__26893),
            .in1(N__25958),
            .in2(N__25938),
            .in3(N__25781),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65691),
            .ce(),
            .sr(N__62903));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_3_LC_9_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_3_LC_9_18_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_3_LC_9_18_4 .LUT_INIT=16'b1010000110110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_3_LC_9_18_4  (
            .in0(N__25779),
            .in1(N__26894),
            .in2(N__25925),
            .in3(N__25899),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65691),
            .ce(),
            .sr(N__62903));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_0_LC_9_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_0_LC_9_18_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_0_LC_9_18_5 .LUT_INIT=16'b1010101000010010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_0_LC_9_18_5  (
            .in0(N__25447),
            .in1(N__26889),
            .in2(N__39345),
            .in3(N__25780),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65691),
            .ce(),
            .sr(N__62903));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_0_LC_9_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_0_LC_9_18_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_0_LC_9_18_6 .LUT_INIT=16'b1010101000010010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_0_LC_9_18_6  (
            .in0(N__25616),
            .in1(N__25523),
            .in2(N__39346),
            .in3(N__25582),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65691),
            .ce(),
            .sr(N__62903));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_1_LC_9_18_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_1_LC_9_18_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_1_LC_9_18_7 .LUT_INIT=16'b1010101100000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_1_LC_9_18_7  (
            .in0(N__25581),
            .in1(N__25545),
            .in2(N__25534),
            .in3(N__25483),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65691),
            .ce(),
            .sr(N__62903));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_c_0_LC_9_19_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_c_0_LC_9_19_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_c_0_LC_9_19_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_c_0_LC_9_19_0  (
            .in0(_gnd_net_),
            .in1(N__25440),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_19_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_9_19_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_9_19_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_9_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_9_19_1  (
            .in0(_gnd_net_),
            .in1(N__25990),
            .in2(_gnd_net_),
            .in3(N__25965),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_9_19_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_9_19_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_9_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_9_19_2  (
            .in0(_gnd_net_),
            .in1(N__25957),
            .in2(_gnd_net_),
            .in3(N__25929),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_9_19_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_9_19_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_9_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_9_19_3  (
            .in0(_gnd_net_),
            .in1(N__25918),
            .in2(_gnd_net_),
            .in3(N__25893),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_4_LC_9_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_4_LC_9_19_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_4_LC_9_19_4 .LUT_INIT=16'b1100000111000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_4_LC_9_19_4  (
            .in0(N__26888),
            .in1(N__25883),
            .in2(N__25782),
            .in3(N__25890),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65706),
            .ce(),
            .sr(N__62890));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_RNIU62F_LC_9_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_RNIU62F_LC_9_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_RNIU62F_LC_9_20_4 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_RNIU62F_LC_9_20_4  (
            .in0(N__27209),
            .in1(N__27149),
            .in2(_gnd_net_),
            .in3(N__31344),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_a2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_m8_0_a2_LC_9_20_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_m8_0_a2_LC_9_20_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_m8_0_a2_LC_9_20_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_m8_0_a2_LC_9_20_5  (
            .in0(N__30515),
            .in1(N__26990),
            .in2(N__30474),
            .in3(N__26933),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIAVP33_14_LC_9_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIAVP33_14_LC_9_20_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIAVP33_14_LC_9_20_6 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIAVP33_14_LC_9_20_6  (
            .in0(N__25857),
            .in1(N__25844),
            .in2(N__25812),
            .in3(N__25809),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_0_LC_9_20_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_0_LC_9_20_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_0_LC_9_20_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_0_LC_9_20_7  (
            .in0(_gnd_net_),
            .in1(N__27208),
            .in2(_gnd_net_),
            .in3(N__27143),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22_LC_9_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22_LC_9_21_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22_LC_9_21_2 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22_LC_9_21_2  (
            .in0(N__27141),
            .in1(N__26142),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net ),
            .ce(N__27236),
            .sr(N__62872));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_21_LC_9_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_21_LC_9_21_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_21_LC_9_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_21_LC_9_21_5  (
            .in0(_gnd_net_),
            .in1(N__27138),
            .in2(_gnd_net_),
            .in3(N__26136),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net ),
            .ce(N__27236),
            .sr(N__62872));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_20_LC_9_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_20_LC_9_21_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_20_LC_9_21_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_20_LC_9_21_6  (
            .in0(N__27140),
            .in1(N__27279),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net ),
            .ce(N__27236),
            .sr(N__62872));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_23_LC_9_21_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_23_LC_9_21_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_23_LC_9_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_23_LC_9_21_7  (
            .in0(_gnd_net_),
            .in1(N__27139),
            .in2(_gnd_net_),
            .in3(N__26130),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_op ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net ),
            .ce(N__27236),
            .sr(N__62872));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_0_LC_9_22_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_0_LC_9_22_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_0_LC_9_22_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_0_LC_9_22_0  (
            .in0(N__26038),
            .in1(N__26114),
            .in2(_gnd_net_),
            .in3(N__26100),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_22_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0 ),
            .clk(N__65744),
            .ce(),
            .sr(N__62864));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_1_LC_9_22_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_1_LC_9_22_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_1_LC_9_22_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_1_LC_9_22_1  (
            .in0(N__26036),
            .in1(N__26096),
            .in2(_gnd_net_),
            .in3(N__26082),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1 ),
            .clk(N__65744),
            .ce(),
            .sr(N__62864));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_2_LC_9_22_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_2_LC_9_22_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_2_LC_9_22_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_2_LC_9_22_2  (
            .in0(N__26039),
            .in1(N__26078),
            .in2(_gnd_net_),
            .in3(N__26064),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2 ),
            .clk(N__65744),
            .ce(),
            .sr(N__62864));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_3_LC_9_22_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_3_LC_9_22_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_3_LC_9_22_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_3_LC_9_22_3  (
            .in0(N__26037),
            .in1(N__26057),
            .in2(_gnd_net_),
            .in3(N__26043),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_3 ),
            .clk(N__65744),
            .ce(),
            .sr(N__62864));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_4_LC_9_22_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_4_LC_9_22_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_4_LC_9_22_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_4_LC_9_22_4  (
            .in0(N__26040),
            .in1(N__26009),
            .in2(_gnd_net_),
            .in3(N__26016),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65744),
            .ce(),
            .sr(N__62864));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_31_LC_10_7_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_31_LC_10_7_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_31_LC_10_7_0 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_31_LC_10_7_0  (
            .in0(N__59555),
            .in1(N__28174),
            .in2(N__62060),
            .in3(N__33951),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65537),
            .ce(N__32516),
            .sr(N__62960));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_31_LC_10_7_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_31_LC_10_7_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_31_LC_10_7_1 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_31_LC_10_7_1  (
            .in0(_gnd_net_),
            .in1(N__50401),
            .in2(N__26339),
            .in3(N__62044),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_17_LC_10_7_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_17_LC_10_7_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_17_LC_10_7_2 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_17_LC_10_7_2  (
            .in0(_gnd_net_),
            .in1(N__26312),
            .in2(N__50409),
            .in3(N__57393),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_455_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_18_LC_10_7_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_18_LC_10_7_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_18_LC_10_7_3 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_18_LC_10_7_3  (
            .in0(_gnd_net_),
            .in1(N__50397),
            .in2(N__26338),
            .in3(N__59834),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_454_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_19_LC_10_7_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_19_LC_10_7_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_19_LC_10_7_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_19_LC_10_7_4  (
            .in0(N__50396),
            .in1(N__26316),
            .in2(_gnd_net_),
            .in3(N__61613),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_453_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_o2_LC_10_8_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_o2_LC_10_8_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_o2_LC_10_8_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_o2_LC_10_8_0  (
            .in0(N__38736),
            .in1(N__38675),
            .in2(N__64317),
            .in3(N__64268),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_6_LC_10_9_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_6_LC_10_9_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_6_LC_10_9_1 .LUT_INIT=16'b0000100000001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_6_LC_10_9_1  (
            .in0(N__63582),
            .in1(N__26320),
            .in2(N__50395),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_463_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_8_LC_10_9_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_8_LC_10_9_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_8_LC_10_9_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_8_LC_10_9_2  (
            .in0(N__63102),
            .in1(_gnd_net_),
            .in2(N__26340),
            .in3(N__50355),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_5_LC_10_9_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_5_LC_10_9_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_5_LC_10_9_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_5_LC_10_9_3  (
            .in0(N__63657),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59558),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65557),
            .ce(N__48722),
            .sr(N__62954));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_6_LC_10_9_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_6_LC_10_9_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_6_LC_10_9_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_6_LC_10_9_4  (
            .in0(N__59557),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63583),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65557),
            .ce(N__48722),
            .sr(N__62954));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_8_LC_10_9_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_8_LC_10_9_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_8_LC_10_9_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_8_LC_10_9_5  (
            .in0(_gnd_net_),
            .in1(N__59556),
            .in2(_gnd_net_),
            .in3(N__63103),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65557),
            .ce(N__48722),
            .sr(N__62954));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec1_0_a2_i_LC_10_9_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec1_0_a2_i_LC_10_9_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec1_0_a2_i_LC_10_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec1_0_a2_i_LC_10_9_6  (
            .in0(N__38891),
            .in1(N__38802),
            .in2(_gnd_net_),
            .in3(N__26655),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_1_LC_10_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_1_LC_10_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_1_LC_10_10_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_1_LC_10_10_0  (
            .in0(N__26613),
            .in1(N__52737),
            .in2(N__26601),
            .in3(N__52524),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_1_LC_10_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_1_LC_10_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_1_LC_10_10_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_1_LC_10_10_1  (
            .in0(_gnd_net_),
            .in1(N__52222),
            .in2(N__26586),
            .in3(N__54603),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_1_LC_10_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_1_LC_10_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_1_LC_10_10_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_1_LC_10_10_2  (
            .in0(N__26583),
            .in1(N__44617),
            .in2(N__44127),
            .in3(N__38382),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_1_LC_10_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_1_LC_10_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_1_LC_10_10_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_1_LC_10_10_3  (
            .in0(N__28422),
            .in1(N__53331),
            .in2(N__26571),
            .in3(N__57800),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_1_LC_10_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_1_LC_10_10_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_1_LC_10_10_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_1_LC_10_10_4  (
            .in0(N__27384),
            .in1(N__33540),
            .in2(N__26568),
            .in3(N__26565),
            .lcout(I2C_top_level_inst1_s_data_oreg_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65571),
            .ce(N__54522),
            .sr(N__64971));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_5_LC_10_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_5_LC_10_12_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_5_LC_10_12_0 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_5_LC_10_12_0  (
            .in0(N__51924),
            .in1(N__26559),
            .in2(N__28392),
            .in3(N__32197),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_5_LC_10_12_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_5_LC_10_12_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_5_LC_10_12_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_5_LC_10_12_1  (
            .in0(N__27495),
            .in1(N__26745),
            .in2(N__26748),
            .in3(N__26703),
            .lcout(I2C_top_level_inst1_s_data_oreg_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65595),
            .ce(N__54516),
            .sr(N__64967));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_5_LC_10_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_5_LC_10_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_5_LC_10_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_5_LC_10_12_2  (
            .in0(N__53012),
            .in1(N__32171),
            .in2(N__53315),
            .in3(N__42216),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_5_LC_10_12_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_5_LC_10_12_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_5_LC_10_12_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_5_LC_10_12_3  (
            .in0(N__26739),
            .in1(N__52772),
            .in2(N__26724),
            .in3(N__52521),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_5_LC_10_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_5_LC_10_12_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_5_LC_10_12_4 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_5_LC_10_12_4  (
            .in0(_gnd_net_),
            .in1(N__52227),
            .in2(N__26706),
            .in3(N__32127),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_6_LC_10_13_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_6_LC_10_13_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_6_LC_10_13_7 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_6_LC_10_13_7  (
            .in0(N__51860),
            .in1(N__26697),
            .in2(N__28359),
            .in3(N__33779),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_LC_10_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_LC_10_14_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_LC_10_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_LC_10_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29146),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ),
            .ce(),
            .sr(N__62923));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m12_LC_10_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m12_LC_10_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m12_LC_10_14_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m12_LC_10_14_2  (
            .in0(_gnd_net_),
            .in1(N__26691),
            .in2(_gnd_net_),
            .in3(N__28874),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQK6I1_LC_10_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQK6I1_LC_10_14_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQK6I1_LC_10_14_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQK6I1_LC_10_14_3  (
            .in0(N__26682),
            .in1(N__29145),
            .in2(N__26676),
            .in3(N__32992),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_7_LC_10_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_7_LC_10_14_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_7_LC_10_14_4 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_7_LC_10_14_4  (
            .in0(N__29235),
            .in1(N__26778),
            .in2(_gnd_net_),
            .in3(N__30137),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ),
            .ce(),
            .sr(N__62923));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_6_LC_10_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_6_LC_10_14_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_6_LC_10_14_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_6_LC_10_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28995),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ),
            .ce(),
            .sr(N__62923));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_5_LC_10_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_5_LC_10_14_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_5_LC_10_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_5_LC_10_14_6  (
            .in0(N__29147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ),
            .ce(),
            .sr(N__62923));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_4_LC_10_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_4_LC_10_14_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_4_LC_10_14_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_4_LC_10_14_7  (
            .in0(_gnd_net_),
            .in1(N__28917),
            .in2(_gnd_net_),
            .in3(N__29234),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net ),
            .ce(),
            .sr(N__62923));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17_LC_10_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17_LC_10_16_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17_LC_10_16_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17_LC_10_16_0  (
            .in0(N__27778),
            .in1(N__26766),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_18_LC_10_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_18_LC_10_16_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_18_LC_10_16_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_18_LC_10_16_1  (
            .in0(_gnd_net_),
            .in1(N__27774),
            .in2(_gnd_net_),
            .in3(N__26772),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_13_LC_10_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_13_LC_10_16_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_13_LC_10_16_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_13_LC_10_16_2  (
            .in0(N__27776),
            .in1(N__27006),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_16_LC_10_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_16_LC_10_16_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_16_LC_10_16_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_16_LC_10_16_3  (
            .in0(_gnd_net_),
            .in1(N__27773),
            .in2(_gnd_net_),
            .in3(N__26760),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_22_LC_10_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_22_LC_10_16_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_22_LC_10_16_4 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_22_LC_10_16_4  (
            .in0(N__27779),
            .in1(N__26838),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_15_LC_10_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_15_LC_10_16_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_15_LC_10_16_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_15_LC_10_16_5  (
            .in0(_gnd_net_),
            .in1(N__27772),
            .in2(_gnd_net_),
            .in3(N__26844),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_14_LC_10_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_14_LC_10_16_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_14_LC_10_16_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_14_LC_10_16_6  (
            .in0(N__27777),
            .in1(N__26754),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_21_LC_10_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_21_LC_10_16_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_21_LC_10_16_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_21_LC_10_16_7  (
            .in0(_gnd_net_),
            .in1(N__27775),
            .in2(_gnd_net_),
            .in3(N__26832),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net ),
            .ce(N__27707),
            .sr(N__62904));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10_LC_10_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10_LC_10_17_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10_LC_10_17_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10_LC_10_17_0  (
            .in0(_gnd_net_),
            .in1(N__27784),
            .in2(_gnd_net_),
            .in3(N__26826),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_20_LC_10_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_20_LC_10_17_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_20_LC_10_17_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_20_LC_10_17_1  (
            .in0(N__27781),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26784),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_9_LC_10_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_9_LC_10_17_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_9_LC_10_17_2 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_9_LC_10_17_2  (
            .in0(_gnd_net_),
            .in1(N__27787),
            .in2(_gnd_net_),
            .in3(N__26820),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_8_LC_10_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_8_LC_10_17_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_8_LC_10_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_8_LC_10_17_3  (
            .in0(N__27783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_11_LC_10_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_11_LC_10_17_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_11_LC_10_17_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_11_LC_10_17_4  (
            .in0(_gnd_net_),
            .in1(N__27785),
            .in2(_gnd_net_),
            .in3(N__26814),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_23_LC_10_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_23_LC_10_17_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_23_LC_10_17_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_23_LC_10_17_5  (
            .in0(N__27782),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26808),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.dout_op ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_19_LC_10_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_19_LC_10_17_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_19_LC_10_17_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_19_LC_10_17_6  (
            .in0(N__26790),
            .in1(N__27786),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_12_LC_10_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_12_LC_10_17_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_12_LC_10_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_12_LC_10_17_7  (
            .in0(N__27780),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27012),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net ),
            .ce(N__27708),
            .sr(N__62891));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_LC_10_18_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_LC_10_18_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_LC_10_18_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_LC_10_18_4  (
            .in0(N__51190),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.s_stop ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__32743),
            .ce(),
            .sr(N__31005));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_en_count_data_i_LC_10_19_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_en_count_data_i_LC_10_19_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_en_count_data_i_LC_10_19_5 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_en_count_data_i_LC_10_19_5  (
            .in0(N__30513),
            .in1(N__27000),
            .in2(N__30471),
            .in3(N__26937),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12_LC_10_20_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12_LC_10_20_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12_LC_10_20_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12_LC_10_20_0  (
            .in0(N__27145),
            .in1(N__27261),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ),
            .ce(N__27235),
            .sr(N__62866));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_15_LC_10_20_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_15_LC_10_20_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_15_LC_10_20_2 .LUT_INIT=16'b1101110111011101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_15_LC_10_20_2  (
            .in0(N__27147),
            .in1(N__26856),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ),
            .ce(N__27235),
            .sr(N__62866));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_13_LC_10_20_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_13_LC_10_20_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_13_LC_10_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_13_LC_10_20_3  (
            .in0(_gnd_net_),
            .in1(N__27144),
            .in2(_gnd_net_),
            .in3(N__26868),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ),
            .ce(N__27235),
            .sr(N__62866));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_14_LC_10_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_14_LC_10_20_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_14_LC_10_20_4 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_14_LC_10_20_4  (
            .in0(N__27146),
            .in1(N__26862),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ),
            .ce(N__27235),
            .sr(N__62866));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_16_LC_10_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_16_LC_10_20_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_16_LC_10_20_6 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_16_LC_10_20_6  (
            .in0(N__27148),
            .in1(N__26850),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net ),
            .ce(N__27235),
            .sr(N__62866));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18_LC_10_21_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18_LC_10_21_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18_LC_10_21_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18_LC_10_21_0  (
            .in0(N__27132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27267),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_19_LC_10_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_19_LC_10_21_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_19_LC_10_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_19_LC_10_21_1  (
            .in0(_gnd_net_),
            .in1(N__27285),
            .in2(_gnd_net_),
            .in3(N__27136),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_8_LC_10_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_8_LC_10_21_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_8_LC_10_21_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_8_LC_10_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27137),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_17_LC_10_21_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_17_LC_10_21_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_17_LC_10_21_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_17_LC_10_21_4  (
            .in0(N__27131),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27273),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_11_LC_10_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_11_LC_10_21_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_11_LC_10_21_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_11_LC_10_21_5  (
            .in0(_gnd_net_),
            .in1(N__27243),
            .in2(_gnd_net_),
            .in3(N__27135),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_9_LC_10_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_9_LC_10_21_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_9_LC_10_21_6 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_9_LC_10_21_6  (
            .in0(N__27133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27255),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_10_LC_10_21_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_10_LC_10_21_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_10_LC_10_21_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_10_LC_10_21_7  (
            .in0(_gnd_net_),
            .in1(N__27249),
            .in2(_gnd_net_),
            .in3(N__27134),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net ),
            .ce(N__27237),
            .sr(N__62860));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_1_0_LC_10_22_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_1_0_LC_10_22_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_1_0_LC_10_22_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_1_0_LC_10_22_0  (
            .in0(_gnd_net_),
            .in1(N__27207),
            .in2(_gnd_net_),
            .in3(N__27142),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_391 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIT2U5_16_LC_10_22_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIT2U5_16_LC_10_22_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIT2U5_16_LC_10_22_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIT2U5_16_LC_10_22_4  (
            .in0(N__28181),
            .in1(N__29367),
            .in2(_gnd_net_),
            .in3(N__27966),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_8_LC_11_8_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_8_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_8_LC_11_8_5 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_8_LC_11_8_5  (
            .in0(N__32382),
            .in1(N__27021),
            .in2(N__53329),
            .in3(N__40698),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_1_LC_11_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_1_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_1_LC_11_9_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_1_LC_11_9_4  (
            .in0(N__38315),
            .in1(N__57834),
            .in2(N__51946),
            .in3(N__54639),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_10_LC_11_9_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_10_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_10_LC_11_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_10_LC_11_9_7  (
            .in0(N__37881),
            .in1(N__43577),
            .in2(N__27372),
            .in3(N__64267),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_830 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_3_LC_11_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_3_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_3_LC_11_10_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_3_LC_11_10_0  (
            .in0(N__53016),
            .in1(N__49676),
            .in2(N__53330),
            .in3(N__49641),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_3_LC_11_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_3_LC_11_10_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_3_LC_11_10_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_3_LC_11_10_1  (
            .in0(N__35553),
            .in1(N__27357),
            .in2(N__27360),
            .in3(N__27318),
            .lcout(I2C_top_level_inst1_s_data_oreg_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65558),
            .ce(N__54520),
            .sr(N__64974));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_3_LC_11_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_3_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_3_LC_11_10_2 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_3_LC_11_10_2  (
            .in0(N__51892),
            .in1(N__27519),
            .in2(N__28500),
            .in3(N__49719),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_3_LC_11_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_3_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_3_LC_11_10_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_3_LC_11_10_3  (
            .in0(N__27351),
            .in1(N__52736),
            .in2(N__27336),
            .in3(N__52523),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_3_LC_11_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_3_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_3_LC_11_10_4 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_3_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__52221),
            .in2(N__27321),
            .in3(N__33741),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_31_LC_11_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_31_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_31_LC_11_11_0 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_31_LC_11_11_0  (
            .in0(N__28449),
            .in1(N__51936),
            .in2(N__38505),
            .in3(N__27390),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_31_LC_11_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_31_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_31_LC_11_11_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_31_LC_11_11_1  (
            .in0(N__52439),
            .in1(N__27312),
            .in2(N__27300),
            .in3(N__52779),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_31_LC_11_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_31_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_31_LC_11_11_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_31_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__46134),
            .in2(N__27468),
            .in3(N__52232),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_31_LC_11_11_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_31_LC_11_11_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_31_LC_11_11_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_31_LC_11_11_3  (
            .in0(N__27465),
            .in1(N__27456),
            .in2(N__27459),
            .in3(N__28152),
            .lcout(I2C_top_level_inst1_s_data_oreg_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65572),
            .ce(N__54517),
            .sr(N__64972));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_31_LC_11_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_31_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_31_LC_11_11_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_31_LC_11_11_4  (
            .in0(N__53445),
            .in1(N__53257),
            .in2(N__46227),
            .in3(N__52987),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_27_LC_11_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_27_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_27_LC_11_12_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_27_LC_11_12_0  (
            .in0(N__27450),
            .in1(N__44533),
            .in2(N__61632),
            .in3(N__44326),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_28_LC_11_12_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_28_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_28_LC_11_12_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_28_LC_11_12_1  (
            .in0(N__44327),
            .in1(N__61544),
            .in2(N__44591),
            .in3(N__27438),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_29_LC_11_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_29_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_29_LC_11_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_29_LC_11_12_2  (
            .in0(N__27426),
            .in1(N__44534),
            .in2(N__61448),
            .in3(N__44328),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_3_LC_11_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_3_LC_11_12_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_3_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_3_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48057),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65583),
            .ce(N__44105),
            .sr(N__64968));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_30_LC_11_12_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_30_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_30_LC_11_12_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_30_LC_11_12_5  (
            .in0(N__44329),
            .in1(N__61318),
            .in2(N__44592),
            .in3(N__27414),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_31_LC_11_12_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_31_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_31_LC_11_12_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_31_LC_11_12_6  (
            .in0(N__27402),
            .in1(N__44541),
            .in2(N__61252),
            .in3(N__44330),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_3_LC_11_13_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_3_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_3_LC_11_13_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_3_LC_11_13_0  (
            .in0(N__44508),
            .in1(N__27540),
            .in2(N__27534),
            .in3(N__44333),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_4_LC_11_13_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_4_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_4_LC_11_13_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_4_LC_11_13_1  (
            .in0(N__44334),
            .in1(N__27510),
            .in2(N__33081),
            .in3(N__44509),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_4_LC_11_13_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_4_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_4_LC_11_13_2 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_4_LC_11_13_2  (
            .in0(N__30174),
            .in1(N__51866),
            .in2(N__27498),
            .in3(N__42486),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_5_LC_11_13_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_5_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_5_LC_11_13_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_5_LC_11_13_3  (
            .in0(N__38302),
            .in1(N__37705),
            .in2(N__32229),
            .in3(N__41127),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_4_LC_11_14_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_4_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_4_LC_11_14_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_4_LC_11_14_0  (
            .in0(N__53015),
            .in1(N__42252),
            .in2(N__53319),
            .in3(N__29697),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_4_LC_11_14_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_4_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_4_LC_11_14_2 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_4_LC_11_14_2  (
            .in0(N__28602),
            .in1(N__52234),
            .in2(_gnd_net_),
            .in3(N__33703),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_4_LC_11_14_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_4_LC_11_14_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_4_LC_11_14_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_4_LC_11_14_3  (
            .in0(N__28137),
            .in1(N__27489),
            .in2(N__27483),
            .in3(N__27480),
            .lcout(I2C_top_level_inst1_s_data_oreg_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65605),
            .ce(N__54507),
            .sr(N__64965));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_0_LC_11_15_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_0_LC_11_15_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_0_LC_11_15_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_0_LC_11_15_0  (
            .in0(N__27599),
            .in1(N__27612),
            .in2(_gnd_net_),
            .in3(N__27474),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_15_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0 ),
            .clk(N__65618),
            .ce(),
            .sr(N__62905));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_1_LC_11_15_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_1_LC_11_15_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_1_LC_11_15_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_1_LC_11_15_1  (
            .in0(N__27596),
            .in1(N__27639),
            .in2(_gnd_net_),
            .in3(N__27471),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1 ),
            .clk(N__65618),
            .ce(),
            .sr(N__62905));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_2_LC_11_15_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_2_LC_11_15_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_2_LC_11_15_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_2_LC_11_15_2  (
            .in0(N__27600),
            .in1(N__27654),
            .in2(_gnd_net_),
            .in3(N__27687),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2 ),
            .clk(N__65618),
            .ce(),
            .sr(N__62905));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_3_LC_11_15_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_3_LC_11_15_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_3_LC_11_15_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_3_LC_11_15_3  (
            .in0(N__27597),
            .in1(N__27627),
            .in2(_gnd_net_),
            .in3(N__27684),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_3 ),
            .clk(N__65618),
            .ce(),
            .sr(N__62905));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_4_LC_11_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_4_LC_11_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_4_LC_11_15_4 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_4_LC_11_15_4  (
            .in0(N__27666),
            .in1(N__27598),
            .in2(_gnd_net_),
            .in3(N__27681),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65618),
            .ce(),
            .sr(N__62905));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1_LC_11_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1_LC_11_16_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1_LC_11_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1_LC_11_16_1  (
            .in0(_gnd_net_),
            .in1(N__27822),
            .in2(_gnd_net_),
            .in3(N__27771),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net ),
            .ce(),
            .sr(N__62892));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_0_LC_11_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_0_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_0_LC_11_16_2 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_0_LC_11_16_2  (
            .in0(N__27770),
            .in1(_gnd_net_),
            .in2(N__27827),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_3_LC_11_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_3_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_3_LC_11_16_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_3_LC_11_16_3  (
            .in0(N__27665),
            .in1(N__27653),
            .in2(N__27642),
            .in3(N__27638),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m7_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_0_LC_11_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_0_LC_11_16_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_0_LC_11_16_4 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_0_LC_11_16_4  (
            .in0(_gnd_net_),
            .in1(N__27626),
            .in2(N__27615),
            .in3(N__27611),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net ),
            .ce(),
            .sr(N__62892));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_LC_11_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_LC_11_16_5 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_LC_11_16_5  (
            .in0(_gnd_net_),
            .in1(N__27817),
            .in2(_gnd_net_),
            .in3(N__27768),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_1_0_LC_11_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_1_0_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_1_0_LC_11_16_6 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_1_0_LC_11_16_6  (
            .in0(N__27823),
            .in1(N__27788),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_0_LC_11_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_0_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_0_LC_11_16_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_0_LC_11_16_7  (
            .in0(_gnd_net_),
            .in1(N__27821),
            .in2(_gnd_net_),
            .in3(N__27769),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIQO531_LC_11_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIQO531_LC_11_17_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIQO531_LC_11_17_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIQO531_LC_11_17_0  (
            .in0(N__28956),
            .in1(N__29074),
            .in2(N__30122),
            .in3(N__30081),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9_LC_11_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9_LC_11_17_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9_LC_11_17_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9_LC_11_17_1  (
            .in0(N__29075),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62882));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_LC_11_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_LC_11_17_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_LC_11_17_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_LC_11_17_2  (
            .in0(N__28957),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62882));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_8_LC_11_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_8_LC_11_17_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_8_LC_11_17_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_8_LC_11_17_3  (
            .in0(_gnd_net_),
            .in1(N__29222),
            .in2(_gnd_net_),
            .in3(N__28887),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62882));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_16_LC_11_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_16_LC_11_17_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_16_LC_11_17_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_16_LC_11_17_5  (
            .in0(_gnd_net_),
            .in1(N__30034),
            .in2(_gnd_net_),
            .in3(N__29221),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62882));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_17_LC_11_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_17_LC_11_17_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_17_LC_11_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_17_LC_11_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29099),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62882));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_3_LC_11_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_3_LC_11_17_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_3_LC_11_17_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_3_LC_11_17_7  (
            .in0(N__29061),
            .in1(N__29037),
            .in2(N__29006),
            .in3(N__28958),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62882));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIE8O3_0_LC_11_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIE8O3_0_LC_11_18_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIE8O3_0_LC_11_18_1 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIE8O3_0_LC_11_18_1  (
            .in0(N__27869),
            .in1(N__27884),
            .in2(N__27855),
            .in3(N__29106),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3_LC_11_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3_LC_11_18_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3_LC_11_18_2 .LUT_INIT=16'b0000101011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3_LC_11_18_2  (
            .in0(N__28909),
            .in1(_gnd_net_),
            .in2(N__27690),
            .in3(N__27912),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net ),
            .ce(),
            .sr(N__62874));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_1_LC_11_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_1_LC_11_18_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_1_LC_11_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_1_LC_11_18_3  (
            .in0(N__29942),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35853),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net ),
            .ce(),
            .sr(N__62874));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_LC_11_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_LC_11_18_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_LC_11_18_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_LC_11_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29190),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net ),
            .ce(),
            .sr(N__62874));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_RNIFTTJ_LC_11_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_RNIFTTJ_LC_11_18_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_RNIFTTJ_LC_11_18_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_RNIFTTJ_LC_11_18_5  (
            .in0(_gnd_net_),
            .in1(N__27911),
            .in2(_gnd_net_),
            .in3(N__28908),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1OR71_LC_11_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1OR71_LC_11_18_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1OR71_LC_11_18_6 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1OR71_LC_11_18_6  (
            .in0(_gnd_net_),
            .in1(N__27900),
            .in2(N__27888),
            .in3(N__29941),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_0_LC_11_19_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_0_LC_11_19_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_0_LC_11_19_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_0_LC_11_19_0  (
            .in0(N__28861),
            .in1(N__27885),
            .in2(_gnd_net_),
            .in3(N__27873),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_11_19_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0 ),
            .clk(N__65669),
            .ce(),
            .sr(N__62867));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_1_LC_11_19_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_1_LC_11_19_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_1_LC_11_19_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_1_LC_11_19_1  (
            .in0(N__28847),
            .in1(N__27870),
            .in2(_gnd_net_),
            .in3(N__27858),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1 ),
            .clk(N__65669),
            .ce(),
            .sr(N__62867));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_2_LC_11_19_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_2_LC_11_19_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_2_LC_11_19_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_2_LC_11_19_2  (
            .in0(N__28862),
            .in1(N__27854),
            .in2(_gnd_net_),
            .in3(N__27840),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2 ),
            .clk(N__65669),
            .ce(),
            .sr(N__62867));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_3_LC_11_19_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_3_LC_11_19_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_3_LC_11_19_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_3_LC_11_19_3  (
            .in0(N__28848),
            .in1(N__29118),
            .in2(_gnd_net_),
            .in3(N__27837),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_3 ),
            .clk(N__65669),
            .ce(),
            .sr(N__62867));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_4_LC_11_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_4_LC_11_19_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_4_LC_11_19_4 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_4_LC_11_19_4  (
            .in0(N__29130),
            .in1(N__28849),
            .in2(_gnd_net_),
            .in3(N__27834),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65669),
            .ce(),
            .sr(N__62867));
    defparam \cemf_module_64ch_ctrl_inst1.ch_cnt_0_LC_11_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.ch_cnt_0_LC_11_21_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.ch_cnt_0_LC_11_21_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.ch_cnt_0_LC_11_21_2  (
            .in0(N__29256),
            .in1(N__36873),
            .in2(_gnd_net_),
            .in3(N__27978),
            .lcout(\cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65694),
            .ce(),
            .sr(N__62854));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_0_LC_11_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_0_LC_11_22_2 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_0_LC_11_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_0_LC_11_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27996),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65714),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNI07M9_LC_11_22_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNI07M9_LC_11_22_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNI07M9_LC_11_22_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNI07M9_LC_11_22_5  (
            .in0(N__27977),
            .in1(N__29405),
            .in2(_gnd_net_),
            .in3(N__27965),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_410_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_410_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m56_i_LC_11_22_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m56_i_LC_11_22_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m56_i_LC_11_22_6 .LUT_INIT=16'b0101111100010011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m56_i_LC_11_22_6  (
            .in0(N__30596),
            .in1(N__31456),
            .in2(N__27954),
            .in3(N__31479),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_68_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_68_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_i_i_0_o2_i_o2_0_4_LC_11_22_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_i_i_0_o2_i_o2_0_4_LC_11_22_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_i_i_0_o2_i_o2_0_4_LC_11_22_7 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_i_i_0_o2_i_o2_0_4_LC_11_22_7  (
            .in0(N__29389),
            .in1(N__35762),
            .in2(N__27951),
            .in3(N__29363),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_reti_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_8_LC_12_7_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_8_LC_12_7_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_8_LC_12_7_1 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_8_LC_12_7_1  (
            .in0(N__37707),
            .in1(N__53011),
            .in2(N__28803),
            .in3(N__40731),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_8_LC_12_8_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_8_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_8_LC_12_8_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_8_LC_12_8_1  (
            .in0(N__38316),
            .in1(N__40759),
            .in2(N__51951),
            .in3(N__41025),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_8_LC_12_8_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_8_LC_12_8_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_8_LC_12_8_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_8_LC_12_8_2  (
            .in0(N__27948),
            .in1(N__52744),
            .in2(N__27933),
            .in3(N__52527),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_8_LC_12_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_8_LC_12_8_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_8_LC_12_8_3 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_8_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(N__52203),
            .in2(N__27915),
            .in3(N__40833),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_8_LC_12_8_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_8_LC_12_8_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_8_LC_12_8_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_8_LC_12_8_4  (
            .in0(N__28125),
            .in1(N__28119),
            .in2(N__28113),
            .in3(N__28110),
            .lcout(I2C_top_level_inst1_s_data_oreg_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65527),
            .ce(N__54523),
            .sr(N__64985));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_14_LC_12_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_14_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_14_LC_12_9_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_14_LC_12_9_0  (
            .in0(N__28104),
            .in1(N__52761),
            .in2(N__28089),
            .in3(N__52520),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_14_LC_12_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_14_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_14_LC_12_9_1 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_14_LC_12_9_1  (
            .in0(N__52206),
            .in1(_gnd_net_),
            .in2(N__28071),
            .in3(N__32097),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_14_LC_12_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_14_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_14_LC_12_9_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_14_LC_12_9_2  (
            .in0(N__44368),
            .in1(N__63568),
            .in2(N__44662),
            .in3(N__28068),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_14_LC_12_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_14_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_14_LC_12_9_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_14_LC_12_9_3  (
            .in0(N__28698),
            .in1(N__51950),
            .in2(N__28053),
            .in3(N__38487),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_14_LC_12_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_14_LC_12_9_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_14_LC_12_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_14_LC_12_9_4  (
            .in0(N__34968),
            .in1(N__30771),
            .in2(N__28050),
            .in3(N__28047),
            .lcout(I2C_top_level_inst1_s_data_oreg_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65538),
            .ce(N__54521),
            .sr(N__64982));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_22_LC_12_9_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_22_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_22_LC_12_9_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_22_LC_12_9_5  (
            .in0(N__28041),
            .in1(N__44635),
            .in2(N__58440),
            .in3(N__44367),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_30_LC_12_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_30_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_30_LC_12_10_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_30_LC_12_10_0  (
            .in0(N__38550),
            .in1(N__53271),
            .in2(N__46293),
            .in3(N__53004),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_30_LC_12_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_30_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_30_LC_12_10_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_30_LC_12_10_1  (
            .in0(N__28026),
            .in1(N__52780),
            .in2(N__28011),
            .in3(N__52445),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_30_LC_12_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_30_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_30_LC_12_10_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_30_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__34026),
            .in2(N__28227),
            .in3(N__52233),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_30_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_30_LC_12_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_30_LC_12_10_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_30_LC_12_10_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_30_LC_12_10_3  (
            .in0(N__28200),
            .in1(N__28224),
            .in2(N__28218),
            .in3(N__28206),
            .lcout(I2C_top_level_inst1_s_data_oreg_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65547),
            .ce(N__54518),
            .sr(N__64978));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_30_LC_12_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_30_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_30_LC_12_10_4 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_30_LC_12_10_4  (
            .in0(N__51925),
            .in1(N__28470),
            .in2(N__38097),
            .in3(N__28215),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_30_LC_12_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_30_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_30_LC_12_11_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_30_LC_12_11_0  (
            .in0(N__28584),
            .in1(N__38276),
            .in2(N__28194),
            .in3(N__37689),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_30_LC_12_11_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_30_LC_12_11_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_30_LC_12_11_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_30_LC_12_11_1  (
            .in0(N__62125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59441),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65559),
            .ce(N__45572),
            .sr(N__62932));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_31_LC_12_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_31_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_31_LC_12_11_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_31_LC_12_11_2  (
            .in0(N__28182),
            .in1(N__38277),
            .in2(N__28146),
            .in3(N__37690),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_31_LC_12_11_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_31_LC_12_11_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_31_LC_12_11_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_31_LC_12_11_3  (
            .in0(N__62024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59442),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65559),
            .ce(N__45572),
            .sr(N__62932));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_4_LC_12_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_4_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_4_LC_12_11_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_4_LC_12_11_4  (
            .in0(N__38268),
            .in1(N__37688),
            .in2(N__28566),
            .in3(N__28325),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_4_LC_12_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_4_LC_12_11_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_4_LC_12_11_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_4_LC_12_11_5  (
            .in0(_gnd_net_),
            .in1(N__63775),
            .in2(_gnd_net_),
            .in3(N__59443),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65559),
            .ce(N__45572),
            .sr(N__62932));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMAFN1_LC_12_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMAFN1_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMAFN1_LC_12_11_6 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMAFN1_LC_12_11_6  (
            .in0(N__55198),
            .in1(N__55438),
            .in2(N__33714),
            .in3(N__28321),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9GQL2_LC_12_11_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9GQL2_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9GQL2_LC_12_11_7 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9GQL2_LC_12_11_7  (
            .in0(N__33710),
            .in1(N__54954),
            .in2(N__28326),
            .in3(N__54757),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_26_LC_12_12_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_26_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_26_LC_12_12_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_26_LC_12_12_1  (
            .in0(N__28311),
            .in1(N__37844),
            .in2(_gnd_net_),
            .in3(N__66815),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_26_LC_12_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_26_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_26_LC_12_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_26_LC_12_12_2  (
            .in0(N__28299),
            .in1(N__32362),
            .in2(N__28281),
            .in3(N__34050),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_1_26_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_26_LC_12_12_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_26_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_26_LC_12_12_3 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_26_LC_12_12_3  (
            .in0(N__33432),
            .in1(N__28263),
            .in2(N__28257),
            .in3(N__28254),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_3_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_26_LC_12_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_26_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_26_LC_12_12_4 .LUT_INIT=16'b0101010100000101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_26_LC_12_12_4  (
            .in0(N__57249),
            .in1(_gnd_net_),
            .in2(N__66819),
            .in3(N__59851),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_LC_12_12_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_LC_12_12_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_LC_12_12_5  (
            .in0(_gnd_net_),
            .in1(N__66814),
            .in2(_gnd_net_),
            .in3(N__57248),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_21_LC_12_12_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_21_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_21_LC_12_12_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_21_LC_12_12_6  (
            .in0(N__64252),
            .in1(N__32363),
            .in2(N__43576),
            .in3(N__28242),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNITSQ5D_0_LC_12_12_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNITSQ5D_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNITSQ5D_0_LC_12_12_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNITSQ5D_0_LC_12_12_7  (
            .in0(N__32361),
            .in1(N__43533),
            .in2(_gnd_net_),
            .in3(N__64251),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1318 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_9_LC_12_13_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_9_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_9_LC_12_13_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_9_LC_12_13_0  (
            .in0(N__64208),
            .in1(N__28542),
            .in2(N__43562),
            .in3(N__37869),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_841 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_29_LC_12_13_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_29_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_29_LC_12_13_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_29_LC_12_13_1  (
            .in0(N__37863),
            .in1(N__28527),
            .in2(N__43575),
            .in3(N__64202),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_632 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_3_LC_12_13_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_3_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_3_LC_12_13_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_3_LC_12_13_2  (
            .in0(N__64204),
            .in1(N__28512),
            .in2(N__43560),
            .in3(N__37866),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_907 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_30_LC_12_13_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_30_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_30_LC_12_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_30_LC_12_13_3  (
            .in0(N__37864),
            .in1(N__43491),
            .in2(N__28488),
            .in3(N__64205),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_621 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_31_LC_12_13_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_31_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_31_LC_12_13_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_31_LC_12_13_4  (
            .in0(N__64201),
            .in1(N__28461),
            .in2(N__43559),
            .in3(N__37865),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_610 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_1_LC_12_13_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_1_LC_12_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_1_LC_12_13_5  (
            .in0(N__32360),
            .in1(N__43492),
            .in2(N__28437),
            .in3(N__64207),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_5_LC_12_13_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_5_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_5_LC_12_13_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_5_LC_12_13_6  (
            .in0(N__64206),
            .in1(N__28410),
            .in2(N__43561),
            .in3(N__37868),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_885 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_6_LC_12_13_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_6_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_6_LC_12_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_6_LC_12_13_7  (
            .in0(N__37867),
            .in1(N__43487),
            .in2(N__28377),
            .in3(N__64203),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_874 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_9_LC_12_14_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_9_LC_12_14_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_9_LC_12_14_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_9_LC_12_14_0  (
            .in0(N__52739),
            .in1(N__28347),
            .in2(N__28656),
            .in3(N__52370),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_4_LC_12_14_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_4_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_4_LC_12_14_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_4_LC_12_14_1  (
            .in0(N__52371),
            .in1(N__28635),
            .in2(N__28620),
            .in3(N__52740),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_9_LC_12_14_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_9_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_9_LC_12_14_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_9_LC_12_14_6  (
            .in0(N__44590),
            .in1(N__28596),
            .in2(N__61862),
            .in3(N__44369),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_0_LC_12_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_0_LC_12_15_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_0_LC_12_15_0 .LUT_INIT=16'b0000110010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_0_LC_12_15_0  (
            .in0(N__40060),
            .in1(N__61971),
            .in2(N__59445),
            .in3(N__33932),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_0_6_LC_12_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_0_6_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_0_6_LC_12_15_1 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_0_6_LC_12_15_1  (
            .in0(N__40000),
            .in1(N__40059),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_349 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_28_LC_12_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_28_LC_12_15_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_28_LC_12_15_2 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_28_LC_12_15_2  (
            .in0(N__35651),
            .in1(N__59275),
            .in2(N__62376),
            .in3(N__33933),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_29_LC_12_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_29_LC_12_15_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_29_LC_12_15_3 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_29_LC_12_15_3  (
            .in0(N__33929),
            .in1(N__62259),
            .in2(N__59446),
            .in3(N__35603),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_3_LC_12_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_3_LC_12_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_3_LC_12_15_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_3_LC_12_15_4  (
            .in0(N__63914),
            .in1(N__59276),
            .in2(N__35573),
            .in3(N__33934),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_30_LC_12_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_30_LC_12_15_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_30_LC_12_15_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_30_LC_12_15_5  (
            .in0(N__33930),
            .in1(N__62147),
            .in2(N__59447),
            .in3(N__28583),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_4_LC_12_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_4_LC_12_15_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_4_LC_12_15_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_4_LC_12_15_6  (
            .in0(N__63822),
            .in1(N__59277),
            .in2(N__28562),
            .in3(N__33935),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_8_LC_12_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_8_LC_12_15_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_8_LC_12_15_7 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_8_LC_12_15_7  (
            .in0(N__33931),
            .in1(N__28796),
            .in2(N__59448),
            .in3(N__63144),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65606),
            .ce(N__32517),
            .sr(N__62893));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_0_LC_12_16_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_0_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_0_LC_12_16_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_0_LC_12_16_0  (
            .in0(N__37805),
            .in1(N__43540),
            .in2(N__28782),
            .in3(N__64213),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_940 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_11_LC_12_16_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_11_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_11_LC_12_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_11_LC_12_16_2  (
            .in0(N__37806),
            .in1(N__43545),
            .in2(N__28764),
            .in3(N__64217),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_819 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_12_LC_12_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_12_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_12_LC_12_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_12_LC_12_16_3  (
            .in0(N__64215),
            .in1(N__28749),
            .in2(N__43579),
            .in3(N__37807),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_808 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_13_LC_12_16_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_13_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_13_LC_12_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_13_LC_12_16_4  (
            .in0(N__37808),
            .in1(N__43541),
            .in2(N__28731),
            .in3(N__64216),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_797 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_14_LC_12_16_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_14_LC_12_16_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_14_LC_12_16_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_14_LC_12_16_5  (
            .in0(N__64218),
            .in1(N__28713),
            .in2(N__43580),
            .in3(N__37809),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_786 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_15_LC_12_16_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_15_LC_12_16_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_15_LC_12_16_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_15_LC_12_16_6  (
            .in0(N__37810),
            .in1(N__43549),
            .in2(N__28686),
            .in3(N__64219),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_775 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_20_LC_12_16_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_20_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_20_LC_12_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_20_LC_12_16_7  (
            .in0(N__64214),
            .in1(N__28665),
            .in2(N__43578),
            .in3(N__32364),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_283 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIT5I21_16_LC_12_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIT5I21_16_LC_12_17_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIT5I21_16_LC_12_17_0 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIT5I21_16_LC_12_17_0  (
            .in0(N__29095),
            .in1(N__32973),
            .in2(N__29041),
            .in3(N__29999),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_LC_12_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_LC_12_17_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_LC_12_17_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_LC_12_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29033),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62875));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m10_LC_12_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m10_LC_12_17_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m10_LC_12_17_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m10_LC_12_17_2  (
            .in0(_gnd_net_),
            .in1(N__28941),
            .in2(_gnd_net_),
            .in3(N__28819),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_19_LC_12_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_19_LC_12_17_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_19_LC_12_17_3 .LUT_INIT=16'b1100110000001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_19_LC_12_17_3  (
            .in0(_gnd_net_),
            .in1(N__28935),
            .in2(N__28920),
            .in3(N__29224),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62875));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_11_LC_12_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_11_LC_12_17_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_11_LC_12_17_4 .LUT_INIT=16'b0101000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_11_LC_12_17_4  (
            .in0(N__29223),
            .in1(_gnd_net_),
            .in2(N__30084),
            .in3(N__30121),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62875));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_0_LC_12_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_0_LC_12_17_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_0_LC_12_17_5 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_0_LC_12_17_5  (
            .in0(N__28820),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30077),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_LC_12_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_LC_12_17_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_LC_12_17_6 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_LC_12_17_6  (
            .in0(N__28910),
            .in1(N__30036),
            .in2(N__28890),
            .in3(N__28886),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_20_LC_12_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_20_LC_12_17_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_20_LC_12_17_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_20_LC_12_17_7  (
            .in0(N__28821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29225),
            .lcout(\cemf_module_64ch_ctrl_inst1.end_conf_b ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62875));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_RNI63PT_LC_12_18_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_RNI63PT_LC_12_18_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_RNI63PT_LC_12_18_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_RNI63PT_LC_12_18_0  (
            .in0(N__28809),
            .in1(N__30026),
            .in2(N__30054),
            .in3(N__29166),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_LC_12_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_LC_12_18_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_LC_12_18_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_LC_12_18_1  (
            .in0(N__29168),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ),
            .ce(),
            .sr(N__62868));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_12_LC_12_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_12_LC_12_18_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_12_LC_12_18_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_12_LC_12_18_2  (
            .in0(_gnd_net_),
            .in1(N__29219),
            .in2(_gnd_net_),
            .in3(N__30083),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ),
            .ce(),
            .sr(N__62868));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_15_LC_12_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_15_LC_12_18_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_15_LC_12_18_3 .LUT_INIT=16'b0101000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_15_LC_12_18_3  (
            .in0(N__29220),
            .in1(_gnd_net_),
            .in2(N__30035),
            .in3(N__30052),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ),
            .ce(),
            .sr(N__62868));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_13_LC_12_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_13_LC_12_18_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_13_LC_12_18_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_13_LC_12_18_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29169),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ),
            .ce(),
            .sr(N__62868));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_LC_12_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_LC_12_18_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_LC_12_18_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_LC_12_18_5  (
            .in0(N__29178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net ),
            .ce(),
            .sr(N__62868));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_1_LC_12_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_1_LC_12_18_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_1_LC_12_18_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_1_LC_12_18_6  (
            .in0(N__29189),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29177),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHNKP_12_LC_12_18_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHNKP_12_LC_12_18_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHNKP_12_LC_12_18_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHNKP_12_LC_12_18_7  (
            .in0(N__29167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29154),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIF6G1_4_LC_12_19_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIF6G1_4_LC_12_19_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIF6G1_4_LC_12_19_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIF6G1_4_LC_12_19_3  (
            .in0(_gnd_net_),
            .in1(N__29129),
            .in2(_gnd_net_),
            .in3(N__29117),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_i_a2_1_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIPVKP_16_LC_12_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIPVKP_16_LC_12_19_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIPVKP_16_LC_12_19_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIPVKP_16_LC_12_19_4  (
            .in0(_gnd_net_),
            .in1(N__29100),
            .in2(_gnd_net_),
            .in3(N__29079),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_LC_12_19_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_LC_12_19_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_LC_12_19_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_LC_12_19_7  (
            .in0(N__29060),
            .in1(N__29048),
            .in2(N__29007),
            .in3(N__28965),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_276i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_0_LC_12_20_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_0_LC_12_20_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_0_LC_12_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_0_LC_12_20_0  (
            .in0(N__31090),
            .in1(N__30285),
            .in2(_gnd_net_),
            .in3(N__29271),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0 ),
            .ltout(),
            .carryin(bfn_12_20_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0 ),
            .clk(N__65670),
            .ce(),
            .sr(N__62855));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_1_LC_12_20_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_1_LC_12_20_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_1_LC_12_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_1_LC_12_20_1  (
            .in0(N__31087),
            .in1(N__30300),
            .in2(_gnd_net_),
            .in3(N__29268),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1 ),
            .clk(N__65670),
            .ce(),
            .sr(N__62855));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_2_LC_12_20_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_2_LC_12_20_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_2_LC_12_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_2_LC_12_20_2  (
            .in0(N__31091),
            .in1(N__30312),
            .in2(_gnd_net_),
            .in3(N__29265),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2 ),
            .clk(N__65670),
            .ce(),
            .sr(N__62855));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_3_LC_12_20_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_3_LC_12_20_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_3_LC_12_20_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_3_LC_12_20_3  (
            .in0(N__31088),
            .in1(N__30324),
            .in2(_gnd_net_),
            .in3(N__29262),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_3 ),
            .clk(N__65670),
            .ce(),
            .sr(N__62855));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_4_LC_12_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_4_LC_12_20_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_4_LC_12_20_4 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_4_LC_12_20_4  (
            .in0(N__30336),
            .in1(N__31089),
            .in2(_gnd_net_),
            .in3(N__29259),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65670),
            .ce(),
            .sr(N__62855));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIFUVN_LC_12_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIFUVN_LC_12_21_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIFUVN_LC_12_21_2 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIFUVN_LC_12_21_2  (
            .in0(N__29390),
            .in1(N__40037),
            .in2(_gnd_net_),
            .in3(N__32825),
            .lcout(\cemf_module_64ch_ctrl_inst1.en_ch_cnt_0_a2_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_0_LC_12_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_0_LC_12_21_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_0_LC_12_21_3 .LUT_INIT=16'b1111010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_0_LC_12_21_3  (
            .in0(N__29250),
            .in1(N__29391),
            .in2(N__31455),
            .in3(N__36839),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un40_0_a2_4_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_m3_i_0_a2_LC_12_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_m3_i_0_a2_LC_12_21_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_m3_i_0_a2_LC_12_21_6 .LUT_INIT=16'b0010101000101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_m3_i_0_a2_LC_12_21_6  (
            .in0(N__32770),
            .in1(N__36869),
            .in2(N__36843),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1945 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_LC_12_22_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_LC_12_22_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_LC_12_22_0 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_LC_12_22_0  (
            .in0(N__30350),
            .in1(N__29366),
            .in2(N__35763),
            .in3(N__29394),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65695),
            .ce(),
            .sr(N__62844));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_LC_12_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_LC_12_22_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_LC_12_22_1 .LUT_INIT=16'b0111011100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_LC_12_22_1  (
            .in0(N__29412),
            .in1(N__31314),
            .in2(_gnd_net_),
            .in3(N__29406),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65695),
            .ce(),
            .sr(N__62844));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_LC_12_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_LC_12_22_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_LC_12_22_2 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_LC_12_22_2  (
            .in0(N__30349),
            .in1(N__29393),
            .in2(_gnd_net_),
            .in3(N__29365),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1844 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65695),
            .ce(),
            .sr(N__62844));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_17_LC_12_22_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_17_LC_12_22_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_17_LC_12_22_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_17_LC_12_22_4  (
            .in0(_gnd_net_),
            .in1(N__29392),
            .in2(_gnd_net_),
            .in3(N__29364),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65695),
            .ce(),
            .sr(N__62844));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_16_LC_12_22_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_16_LC_12_22_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_16_LC_12_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_16_LC_12_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35757),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65695),
            .ce(),
            .sr(N__62844));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIANE51_11_LC_12_23_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIANE51_11_LC_12_23_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIANE51_11_LC_12_23_2 .LUT_INIT=16'b0101011101010101;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIANE51_11_LC_12_23_2  (
            .in0(N__36552),
            .in1(N__63281),
            .in2(N__41529),
            .in3(N__50994),
            .lcout(sda_o),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_22_LC_13_7_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_22_LC_13_7_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_22_LC_13_7_0 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_22_LC_13_7_0  (
            .in0(N__52223),
            .in1(N__29277),
            .in2(_gnd_net_),
            .in3(N__38607),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_22_LC_13_7_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_22_LC_13_7_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_22_LC_13_7_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_22_LC_13_7_1  (
            .in0(N__30744),
            .in1(N__29316),
            .in2(N__29319),
            .in3(N__29532),
            .lcout(I2C_top_level_inst1_s_data_oreg_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65518),
            .ce(N__54524),
            .sr(N__64996));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_22_LC_13_7_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_22_LC_13_7_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_22_LC_13_7_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_22_LC_13_7_2  (
            .in0(N__42279),
            .in1(N__53010),
            .in2(N__53328),
            .in3(N__38532),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_22_LC_13_7_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_22_LC_13_7_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_22_LC_13_7_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_22_LC_13_7_3  (
            .in0(N__29310),
            .in1(N__52743),
            .in2(N__29295),
            .in3(N__52438),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_22_LC_13_8_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_22_LC_13_8_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_22_LC_13_8_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_22_LC_13_8_5  (
            .in0(N__51903),
            .in1(N__29538),
            .in2(N__33324),
            .in3(N__38436),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_28_LC_13_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_28_LC_13_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_28_LC_13_9_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_28_LC_13_9_0  (
            .in0(N__54177),
            .in1(N__53270),
            .in2(N__40623),
            .in3(N__52994),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_28_LC_13_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_28_LC_13_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_28_LC_13_9_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_28_LC_13_9_1  (
            .in0(N__29526),
            .in1(N__52768),
            .in2(N__29514),
            .in3(N__52486),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_28_LC_13_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_28_LC_13_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_28_LC_13_9_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_28_LC_13_9_2  (
            .in0(_gnd_net_),
            .in1(N__49128),
            .in2(N__29496),
            .in3(N__52213),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_28_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_28_LC_13_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_28_LC_13_9_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_28_LC_13_9_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_28_LC_13_9_3  (
            .in0(N__35631),
            .in1(N__29493),
            .in2(N__29487),
            .in3(N__29472),
            .lcout(I2C_top_level_inst1_s_data_oreg_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65528),
            .ce(N__54519),
            .sr(N__64986));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_28_LC_13_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_28_LC_13_9_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_28_LC_13_9_4 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_28_LC_13_9_4  (
            .in0(N__29823),
            .in1(N__51904),
            .in2(N__48795),
            .in3(N__29484),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_15_LC_13_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_15_LC_13_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_15_LC_13_10_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_15_LC_13_10_0  (
            .in0(N__29466),
            .in1(N__52700),
            .in2(N__29448),
            .in3(N__52488),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_15_LC_13_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_15_LC_13_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_15_LC_13_10_1 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_15_LC_13_10_1  (
            .in0(N__52182),
            .in1(_gnd_net_),
            .in2(N__29430),
            .in3(N__46605),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_15_LC_13_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_15_LC_13_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_15_LC_13_10_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_15_LC_13_10_2  (
            .in0(N__44407),
            .in1(N__63481),
            .in2(N__44659),
            .in3(N__29427),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_15_LC_13_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_15_LC_13_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_15_LC_13_10_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_15_LC_13_10_3  (
            .in0(N__29661),
            .in1(N__51859),
            .in2(N__29649),
            .in3(N__48581),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_15_LC_13_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_15_LC_13_10_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_15_LC_13_10_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_15_LC_13_10_4  (
            .in0(N__34923),
            .in1(N__30759),
            .in2(N__29646),
            .in3(N__29643),
            .lcout(I2C_top_level_inst1_s_data_oreg_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65539),
            .ce(N__54513),
            .sr(N__64983));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_23_LC_13_10_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_23_LC_13_10_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_23_LC_13_10_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_23_LC_13_10_5  (
            .in0(N__29637),
            .in1(N__44624),
            .in2(N__57475),
            .in3(N__44406),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_17_LC_13_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_17_LC_13_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_17_LC_13_11_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_17_LC_13_11_0  (
            .in0(N__52742),
            .in1(N__29622),
            .in2(N__29604),
            .in3(N__52487),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_17_LC_13_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_17_LC_13_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_17_LC_13_11_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_17_LC_13_11_1  (
            .in0(_gnd_net_),
            .in1(N__52215),
            .in2(N__29586),
            .in3(N__46563),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_17_LC_13_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_17_LC_13_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_17_LC_13_11_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_17_LC_13_11_2  (
            .in0(N__44332),
            .in1(N__29583),
            .in2(N__46507),
            .in3(N__44548),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_17_LC_13_11_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_17_LC_13_11_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_17_LC_13_11_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_17_LC_13_11_3  (
            .in0(N__33135),
            .in1(N__51919),
            .in2(N__29568),
            .in3(N__51624),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_17_LC_13_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_17_LC_13_11_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_17_LC_13_11_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_17_LC_13_11_4  (
            .in0(N__35316),
            .in1(N__30804),
            .in2(N__29565),
            .in3(N__29562),
            .lcout(I2C_top_level_inst1_s_data_oreg_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65548),
            .ce(N__54510),
            .sr(N__64979));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_25_LC_13_11_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_25_LC_13_11_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_25_LC_13_11_5 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_25_LC_13_11_5  (
            .in0(N__44547),
            .in1(N__29556),
            .in2(N__57374),
            .in3(N__44331),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIUMB92_17_LC_13_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIUMB92_17_LC_13_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIUMB92_17_LC_13_12_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIUMB92_17_LC_13_12_0  (
            .in0(N__57978),
            .in1(N__58156),
            .in2(N__42481),
            .in3(N__29689),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3Q5_LC_13_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3Q5_LC_13_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3Q5_LC_13_12_1 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3Q5_LC_13_12_1  (
            .in0(N__60474),
            .in1(N__42247),
            .in2(N__29715),
            .in3(N__29712),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3QZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_4_LC_13_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_4_LC_13_12_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_4_LC_13_12_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_4_LC_13_12_2  (
            .in0(_gnd_net_),
            .in1(N__63785),
            .in2(_gnd_net_),
            .in3(N__59444),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65560),
            .ce(N__54113),
            .sr(N__62914));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0FK93_LC_13_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0FK93_LC_13_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0FK93_LC_13_12_3 .LUT_INIT=16'b1111010100110001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0FK93_LC_13_12_3  (
            .in0(N__42482),
            .in1(N__42248),
            .in2(N__46041),
            .in3(N__45867),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRL7_LC_13_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRL7_LC_13_12_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRL7_LC_13_12_4 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRL7_LC_13_12_4  (
            .in0(N__53959),
            .in1(N__29706),
            .in2(N__29700),
            .in3(N__29690),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7LCO7_LC_13_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7LCO7_LC_13_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7LCO7_LC_13_12_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7LCO7_LC_13_12_5  (
            .in0(N__53672),
            .in1(_gnd_net_),
            .in2(N__29676),
            .in3(N__30905),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0RV43_LC_13_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0RV43_LC_13_12_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0RV43_LC_13_12_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0RV43_LC_13_12_6  (
            .in0(N__45866),
            .in1(N__45992),
            .in2(N__38077),
            .in3(N__46270),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_6_LC_13_13_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_6_LC_13_13_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_6_LC_13_13_0 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_6_LC_13_13_0  (
            .in0(N__52220),
            .in1(N__29760),
            .in2(_gnd_net_),
            .in3(N__33678),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_6_LC_13_13_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_6_LC_13_13_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_6_LC_13_13_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_6_LC_13_13_1  (
            .in0(N__32049),
            .in1(N__29808),
            .in2(N__29673),
            .in3(N__29670),
            .lcout(I2C_top_level_inst1_s_data_oreg_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65573),
            .ce(N__54503),
            .sr(N__64973));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_6_LC_13_13_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_6_LC_13_13_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_6_LC_13_13_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_6_LC_13_13_2  (
            .in0(N__31985),
            .in1(N__53281),
            .in2(N__53013),
            .in3(N__42175),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_6_LC_13_13_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_6_LC_13_13_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_6_LC_13_13_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_6_LC_13_13_3  (
            .in0(N__52741),
            .in1(N__29802),
            .in2(N__29781),
            .in3(N__52437),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_9_LC_13_14_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_9_LC_13_14_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_9_LC_13_14_0 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_9_LC_13_14_0  (
            .in0(N__51906),
            .in1(N__29754),
            .in2(N__29748),
            .in3(N__49386),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_9_LC_13_14_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_9_LC_13_14_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_9_LC_13_14_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_9_LC_13_14_1  (
            .in0(N__30885),
            .in1(N__29724),
            .in2(N__29739),
            .in3(N__29730),
            .lcout(I2C_top_level_inst1_s_data_oreg_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65584),
            .ce(N__54502),
            .sr(N__64969));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_9_LC_13_14_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_9_LC_13_14_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_9_LC_13_14_2 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_9_LC_13_14_2  (
            .in0(N__29736),
            .in1(N__52216),
            .in2(_gnd_net_),
            .in3(N__46641),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_9_LC_13_14_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_9_LC_13_14_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_9_LC_13_14_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_9_LC_13_14_4  (
            .in0(N__52990),
            .in1(N__49842),
            .in2(N__53316),
            .in3(N__49423),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI0PB92_17_LC_13_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI0PB92_17_LC_13_15_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI0PB92_17_LC_13_15_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI0PB92_17_LC_13_15_0  (
            .in0(N__58112),
            .in1(N__57941),
            .in2(N__32172),
            .in3(N__32207),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3Q5_LC_13_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3Q5_LC_13_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3Q5_LC_13_15_1 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3Q5_LC_13_15_1  (
            .in0(N__60472),
            .in1(N__42208),
            .in2(N__29718),
            .in3(N__29814),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3QZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6_LC_13_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6_LC_13_15_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6_LC_13_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6_LC_13_15_2  (
            .in0(N__60149),
            .in1(N__29862),
            .in2(_gnd_net_),
            .in3(N__29888),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net ),
            .ce(N__59940),
            .sr(N__62883));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI2RB92_17_LC_13_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI2RB92_17_LC_13_15_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI2RB92_17_LC_13_15_3 .LUT_INIT=16'b1011101100001011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI2RB92_17_LC_13_15_3  (
            .in0(N__57942),
            .in1(N__31989),
            .in2(N__33786),
            .in3(N__58113),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3Q5_LC_13_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3Q5_LC_13_15_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3Q5_LC_13_15_4 .LUT_INIT=16'b0011111110111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3Q5_LC_13_15_4  (
            .in0(N__42177),
            .in1(N__32001),
            .in2(N__29895),
            .in3(N__60473),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNII2U76_LC_13_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNII2U76_LC_13_15_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNII2U76_LC_13_15_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNII2U76_LC_13_15_5  (
            .in0(N__60355),
            .in1(_gnd_net_),
            .in2(N__29892),
            .in3(N__29889),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIDTT76_LC_13_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIDTT76_LC_13_15_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIDTT76_LC_13_15_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIDTT76_LC_13_15_6  (
            .in0(N__29877),
            .in1(N__60354),
            .in2(_gnd_net_),
            .in3(N__29871),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_5_LC_13_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_5_LC_13_15_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_5_LC_13_15_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_5_LC_13_15_7  (
            .in0(N__30822),
            .in1(_gnd_net_),
            .in2(N__29865),
            .in3(N__60148),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net ),
            .ce(N__59940),
            .sr(N__62883));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIPJAS1_1_LC_13_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIPJAS1_1_LC_13_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIPJAS1_1_LC_13_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIPJAS1_1_LC_13_16_0  (
            .in0(N__39653),
            .in1(N__46817),
            .in2(_gnd_net_),
            .in3(N__39140),
            .lcout(N_1614),
            .ltout(N_1614_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_a2_LC_13_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_a2_LC_13_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_a2_LC_13_16_1 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_a2_LC_13_16_1  (
            .in0(_gnd_net_),
            .in1(N__29856),
            .in2(N__29841),
            .in3(N__36201),
            .lcout(N_979),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_28_LC_13_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_28_LC_13_16_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_28_LC_13_16_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_28_LC_13_16_3  (
            .in0(N__43512),
            .in1(N__29838),
            .in2(N__37823),
            .in3(N__64153),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_643 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOCFN1_LC_13_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOCFN1_LC_13_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOCFN1_LC_13_16_5 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOCFN1_LC_13_16_5  (
            .in0(N__55351),
            .in1(N__55113),
            .in2(N__41125),
            .in3(N__32123),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_4_LC_13_16_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_4_LC_13_16_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_4_LC_13_16_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_4_LC_13_16_7  (
            .in0(N__43511),
            .in1(N__30186),
            .in2(N__37824),
            .in3(N__64152),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_896 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIR6CE2_0_LC_13_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIR6CE2_0_LC_13_17_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIR6CE2_0_LC_13_17_0 .LUT_INIT=16'b0010000010100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIR6CE2_0_LC_13_17_0  (
            .in0(N__30259),
            .in1(N__29920),
            .in2(N__29988),
            .in3(N__35854),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_291_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_LC_13_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_LC_13_17_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_LC_13_17_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_LC_13_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30162),
            .in3(N__30159),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_retZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net ),
            .ce(),
            .sr(N__62869));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_RNIB3H2_LC_13_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_RNIB3H2_LC_13_17_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_RNIB3H2_LC_13_17_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_RNIB3H2_LC_13_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30150),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNO_0_0_LC_13_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNO_0_0_LC_13_17_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNO_0_0_LC_13_17_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNO_0_0_LC_13_17_3  (
            .in0(N__30242),
            .in1(N__29986),
            .in2(N__30264),
            .in3(N__30989),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_LC_13_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_LC_13_17_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_LC_13_17_4 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_LC_13_17_4  (
            .in0(N__30238),
            .in1(N__32982),
            .in2(N__30144),
            .in3(N__35856),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net ),
            .ce(),
            .sr(N__62869));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5EOM1_LC_13_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5EOM1_LC_13_17_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5EOM1_LC_13_17_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5EOM1_LC_13_17_5  (
            .in0(N__30141),
            .in1(N__30123),
            .in2(N__30099),
            .in3(N__30082),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_LC_13_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_LC_13_17_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_LC_13_17_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_LC_13_17_6  (
            .in0(N__30053),
            .in1(N__30033),
            .in2(N__30003),
            .in3(N__30000),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_LC_13_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_LC_13_17_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_LC_13_17_7 .LUT_INIT=16'b0100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_LC_13_17_7  (
            .in0(N__35855),
            .in1(N__29987),
            .in2(N__29940),
            .in3(N__30260),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net ),
            .ce(),
            .sr(N__62869));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_LC_13_18_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_LC_13_18_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_LC_13_18_0 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_LC_13_18_0  (
            .in0(_gnd_net_),
            .in1(N__30555),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ),
            .ce(),
            .sr(N__62861));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_RNIJA1F_LC_13_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_RNIJA1F_LC_13_18_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_RNIJA1F_LC_13_18_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_RNIJA1F_LC_13_18_1  (
            .in0(_gnd_net_),
            .in1(N__30219),
            .in2(_gnd_net_),
            .in3(N__31123),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_o3_i_a2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI0RBC1_LC_13_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI0RBC1_LC_13_18_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI0RBC1_LC_13_18_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI0RBC1_LC_13_18_2  (
            .in0(N__30210),
            .in1(N__30554),
            .in2(N__30213),
            .in3(N__32884),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_LC_13_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_LC_13_18_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_LC_13_18_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_LC_13_18_3  (
            .in0(N__30203),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ),
            .ce(),
            .sr(N__62861));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_5_LC_13_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_5_LC_13_18_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_5_LC_13_18_4 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_5_LC_13_18_4  (
            .in0(_gnd_net_),
            .in1(N__30556),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ),
            .ce(),
            .sr(N__62861));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_6_LC_13_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_6_LC_13_18_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_6_LC_13_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_6_LC_13_18_5  (
            .in0(N__30204),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ),
            .ce(),
            .sr(N__62861));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI496Q_5_LC_13_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI496Q_5_LC_13_18_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI496Q_5_LC_13_18_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI496Q_5_LC_13_18_6  (
            .in0(_gnd_net_),
            .in1(N__30380),
            .in2(_gnd_net_),
            .in3(N__30202),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m20_0_a2_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_10_LC_13_18_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_10_LC_13_18_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_10_LC_13_18_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_10_LC_13_18_7  (
            .in0(N__30381),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net ),
            .ce(),
            .sr(N__62861));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11_LC_13_19_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11_LC_13_19_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11_LC_13_19_0 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11_LC_13_19_0  (
            .in0(N__30192),
            .in1(N__31029),
            .in2(_gnd_net_),
            .in3(N__31255),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .ce(),
            .sr(N__62856));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_4_LC_13_19_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_4_LC_13_19_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_4_LC_13_19_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_4_LC_13_19_1  (
            .in0(N__31256),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31385),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .ce(),
            .sr(N__62856));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNIDC2S_4_LC_13_19_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNIDC2S_4_LC_13_19_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNIDC2S_4_LC_13_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNIDC2S_4_LC_13_19_2  (
            .in0(_gnd_net_),
            .in1(N__30335),
            .in2(_gnd_net_),
            .in3(N__30323),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ns_i_a2_1_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNI9N562_0_LC_13_19_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNI9N562_0_LC_13_19_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNI9N562_0_LC_13_19_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNI9N562_0_LC_13_19_3  (
            .in0(N__30311),
            .in1(N__30299),
            .in2(N__30288),
            .in3(N__30284),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_3_LC_13_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_3_LC_13_19_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_3_LC_13_19_4 .LUT_INIT=16'b1100101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_3_LC_13_19_4  (
            .in0(N__31386),
            .in1(N__30270),
            .in2(N__30273),
            .in3(N__31364),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .ce(),
            .sr(N__62856));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_8_LC_13_19_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_8_LC_13_19_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_8_LC_13_19_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_8_LC_13_19_5  (
            .in0(N__31257),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31124),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .ce(),
            .sr(N__62856));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_2_LC_13_19_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_2_LC_13_19_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_2_LC_13_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_2_LC_13_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32568),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .ce(),
            .sr(N__62856));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_10_LC_13_19_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_10_LC_13_19_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_10_LC_13_19_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_10_LC_13_19_7  (
            .in0(N__32567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net ),
            .ce(),
            .sr(N__62856));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIF2FF_12_LC_13_20_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIF2FF_12_LC_13_20_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIF2FF_12_LC_13_20_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIF2FF_12_LC_13_20_0  (
            .in0(N__31283),
            .in1(N__30557),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_LC_13_20_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_LC_13_20_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_LC_13_20_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_LC_13_20_1  (
            .in0(N__31086),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60127),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_0_LC_13_20_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_0_LC_13_20_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_0_LC_13_20_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_0_LC_13_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30561),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_1_0_LC_13_20_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_1_0_LC_13_20_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_1_0_LC_13_20_3 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_1_0_LC_13_20_3  (
            .in0(N__30558),
            .in1(N__31336),
            .in2(_gnd_net_),
            .in3(N__32697),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_0_0_LC_13_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_0_0_LC_13_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_0_0_LC_13_20_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_0_0_LC_13_20_4  (
            .in0(N__31284),
            .in1(N__30537),
            .in2(N__30531),
            .in3(N__31161),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_LC_13_20_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_LC_13_20_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_LC_13_20_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_LC_13_20_5  (
            .in0(N__31162),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C_net ),
            .ce(),
            .sr(N__62849));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIO27J_LC_13_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIO27J_LC_13_20_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIO27J_LC_13_20_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIO27J_LC_13_20_6  (
            .in0(N__30363),
            .in1(N__31026),
            .in2(N__30528),
            .in3(N__31160),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9_LC_13_21_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9_LC_13_21_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9_LC_13_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9_LC_13_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31173),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62845));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_10_LC_13_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_10_LC_13_21_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_10_LC_13_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_10_LC_13_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30519),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62845));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_7_LC_13_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_7_LC_13_21_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_7_LC_13_21_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_7_LC_13_21_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30379),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net ),
            .ce(),
            .sr(N__62845));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_19_LC_13_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_19_LC_13_22_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_19_LC_13_22_1 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_19_LC_13_22_1  (
            .in0(_gnd_net_),
            .in1(N__30354),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_state_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65681),
            .ce(),
            .sr(N__62838));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_LC_13_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_LC_13_22_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_LC_13_22_2 .LUT_INIT=16'b0000101110111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_LC_13_22_2  (
            .in0(N__30609),
            .in1(N__30595),
            .in2(N__31458),
            .in3(N__31478),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65681),
            .ce(),
            .sr(N__62838));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m59_i_LC_13_22_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m59_i_LC_13_22_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m59_i_LC_13_22_3 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m59_i_LC_13_22_3  (
            .in0(N__31451),
            .in1(N__31477),
            .in2(N__30597),
            .in3(N__30608),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_1816_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_7_LC_13_22_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_7_LC_13_22_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_7_LC_13_22_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_7_LC_13_22_7  (
            .in0(_gnd_net_),
            .in1(N__40111),
            .in2(_gnd_net_),
            .in3(N__40001),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_state_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65681),
            .ce(),
            .sr(N__62838));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_0_LC_13_23_0 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_0_LC_13_23_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_0_LC_13_23_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_0_LC_13_23_0  (
            .in0(_gnd_net_),
            .in1(N__34272),
            .in2(N__31590),
            .in3(N__31589),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_0 ),
            .ltout(),
            .carryin(bfn_13_23_0_),
            .carryout(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_1_LC_13_23_1 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_1_LC_13_23_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_1_LC_13_23_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_1_LC_13_23_1  (
            .in0(_gnd_net_),
            .in1(N__34190),
            .in2(_gnd_net_),
            .in3(N__30576),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_1 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0 ),
            .carryout(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_2_LC_13_23_2 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_2_LC_13_23_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_2_LC_13_23_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_2_LC_13_23_2  (
            .in0(_gnd_net_),
            .in1(N__34244),
            .in2(_gnd_net_),
            .in3(N__30573),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_2 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1 ),
            .carryout(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_3_LC_13_23_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_3_LC_13_23_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_3_LC_13_23_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_3_LC_13_23_3  (
            .in0(_gnd_net_),
            .in1(N__34217),
            .in2(_gnd_net_),
            .in3(N__30570),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetter_LC_13_24_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetter_LC_13_24_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetter_LC_13_24_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetter_LC_13_24_5  (
            .in0(N__50820),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetterZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47997),
            .ce(),
            .sr(N__62829));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_RNO_LC_13_25_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_RNO_LC_13_25_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_RNO_LC_13_25_0 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_RNO_LC_13_25_0  (
            .in0(N__30567),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35457),
            .lcout(\I2C_top_level_inst1.I2C_Control_StartUp_inst.rst_neg_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_LC_13_26_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_LC_13_26_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_LC_13_26_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_LC_13_26_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51186),
            .lcout(\I2C_top_level_inst1.s_start ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC_net ),
            .ce(),
            .sr(N__30753));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_22_LC_14_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_22_LC_14_8_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_22_LC_14_8_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_22_LC_14_8_3  (
            .in0(N__37701),
            .in1(N__42681),
            .in2(N__38304),
            .in3(N__30867),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_2_LC_14_8_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_2_LC_14_8_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_2_LC_14_8_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_2_LC_14_8_7  (
            .in0(N__30738),
            .in1(N__44675),
            .in2(N__32925),
            .in3(N__44418),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_13_LC_14_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_13_LC_14_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_13_LC_14_9_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_13_LC_14_9_0  (
            .in0(N__30720),
            .in1(N__52760),
            .in2(N__30708),
            .in3(N__52471),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_13_LC_14_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_13_LC_14_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_13_LC_14_9_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_13_LC_14_9_1  (
            .in0(_gnd_net_),
            .in1(N__52205),
            .in2(N__30690),
            .in3(N__46173),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_13_LC_14_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_13_LC_14_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_13_LC_14_9_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_13_LC_14_9_2  (
            .in0(N__30687),
            .in1(N__44663),
            .in2(N__63670),
            .in3(N__44413),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_13_LC_14_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_13_LC_14_9_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_13_LC_14_9_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_13_LC_14_9_3  (
            .in0(N__30672),
            .in1(N__51902),
            .in2(N__30657),
            .in3(N__38079),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_13_LC_14_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_13_LC_14_9_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_13_LC_14_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_13_LC_14_9_4  (
            .in0(N__35004),
            .in1(N__30654),
            .in2(N__30648),
            .in3(N__30780),
            .lcout(I2C_top_level_inst1_s_data_oreg_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65522),
            .ce(N__54514),
            .sr(N__64992));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_18_LC_14_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_18_LC_14_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_18_LC_14_10_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_18_LC_14_10_0  (
            .in0(N__30645),
            .in1(N__38373),
            .in2(N__30630),
            .in3(N__52701),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_18_LC_14_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_18_LC_14_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_18_LC_14_10_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_18_LC_14_10_1  (
            .in0(_gnd_net_),
            .in1(N__52186),
            .in2(N__30798),
            .in3(N__49173),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_18_LC_14_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_18_LC_14_10_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_18_LC_14_10_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_18_LC_14_10_2  (
            .in0(N__33498),
            .in1(N__30786),
            .in2(N__30795),
            .in3(N__30792),
            .lcout(I2C_top_level_inst1_s_data_oreg_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65529),
            .ce(N__54511),
            .sr(N__64987));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_18_LC_14_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_18_LC_14_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_18_LC_14_10_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_18_LC_14_10_3  (
            .in0(N__32412),
            .in1(N__38303),
            .in2(N__31626),
            .in3(N__48862),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_18_LC_14_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_18_LC_14_10_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_18_LC_14_10_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_18_LC_14_10_4  (
            .in0(N__53258),
            .in1(N__51438),
            .in2(N__51905),
            .in3(N__51402),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_10_LC_14_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_10_LC_14_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_10_LC_14_11_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_10_LC_14_11_0  (
            .in0(N__49340),
            .in1(N__52923),
            .in2(N__53256),
            .in3(N__49269),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_11_LC_14_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_11_LC_14_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_11_LC_14_11_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_11_LC_14_11_1  (
            .in0(N__52925),
            .in1(N__46380),
            .in2(N__53262),
            .in3(N__42527),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_13_LC_14_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_13_LC_14_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_13_LC_14_11_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_13_LC_14_11_2  (
            .in0(N__53179),
            .in1(N__46272),
            .in2(N__40896),
            .in3(N__52924),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_14_LC_14_11_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_14_LC_14_11_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_14_LC_14_11_3 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_14_LC_14_11_3  (
            .in0(N__52922),
            .in1(N__33564),
            .in2(N__53430),
            .in3(N__53175),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_15_LC_14_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_15_LC_14_11_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_15_LC_14_11_4 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_15_LC_14_11_4  (
            .in0(N__53180),
            .in1(N__52926),
            .in2(N__53382),
            .in3(N__46212),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_17_LC_14_11_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_17_LC_14_11_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_17_LC_14_11_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_17_LC_14_11_6  (
            .in0(N__53181),
            .in1(N__52927),
            .in2(N__54165),
            .in3(N__51586),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_1_LC_14_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_1_LC_14_12_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_1_LC_14_12_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_1_LC_14_12_0  (
            .in0(_gnd_net_),
            .in1(N__61861),
            .in2(_gnd_net_),
            .in3(N__59142),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_2_LC_14_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_2_LC_14_12_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_2_LC_14_12_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_2_LC_14_12_1  (
            .in0(N__59145),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61729),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_3_LC_14_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_3_LC_14_12_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_3_LC_14_12_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_3_LC_14_12_2  (
            .in0(N__63910),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59149),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_5_LC_14_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_5_LC_14_12_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_5_LC_14_12_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_5_LC_14_12_3  (
            .in0(N__59146),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63645),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_6_LC_14_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_6_LC_14_12_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_6_LC_14_12_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_6_LC_14_12_4  (
            .in0(_gnd_net_),
            .in1(N__63526),
            .in2(_gnd_net_),
            .in3(N__59143),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_7_LC_14_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_7_LC_14_12_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_7_LC_14_12_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_7_LC_14_12_5  (
            .in0(N__59147),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63467),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_8_LC_14_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_8_LC_14_12_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_8_LC_14_12_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_8_LC_14_12_6  (
            .in0(_gnd_net_),
            .in1(N__59144),
            .in2(_gnd_net_),
            .in3(N__63119),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_9_LC_14_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_9_LC_14_12_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_9_LC_14_12_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_9_LC_14_12_7  (
            .in0(N__59148),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46525),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65549),
            .ce(N__54112),
            .sr(N__62906));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMMQI1_LC_14_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMMQI1_LC_14_13_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMMQI1_LC_14_13_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMMQI1_LC_14_13_0  (
            .in0(N__55221),
            .in1(N__55399),
            .in2(N__46172),
            .in3(N__42812),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GH5_LC_14_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GH5_LC_14_13_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GH5_LC_14_13_1 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GH5_LC_14_13_1  (
            .in0(N__46271),
            .in1(N__60540),
            .in2(N__30852),
            .in3(N__30813),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOJAV5_LC_14_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOJAV5_LC_14_13_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOJAV5_LC_14_13_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOJAV5_LC_14_13_2  (
            .in0(_gnd_net_),
            .in1(N__60329),
            .in2(N__30849),
            .in3(N__30846),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13_LC_14_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13_LC_14_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13_LC_14_13_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13_LC_14_13_3  (
            .in0(_gnd_net_),
            .in1(N__41256),
            .in2(N__30840),
            .in3(N__60150),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net ),
            .ce(N__60005),
            .sr(N__62894));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI8OT76_LC_14_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI8OT76_LC_14_13_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI8OT76_LC_14_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI8OT76_LC_14_13_4  (
            .in0(N__30831),
            .in1(N__60328),
            .in2(_gnd_net_),
            .in3(N__30837),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_4_LC_14_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_4_LC_14_13_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_4_LC_14_13_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_4_LC_14_13_5  (
            .in0(N__49983),
            .in1(_gnd_net_),
            .in2(N__30825),
            .in3(N__60151),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net ),
            .ce(N__60005),
            .sr(N__62894));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU1492_17_LC_14_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU1492_17_LC_14_13_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU1492_17_LC_14_13_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU1492_17_LC_14_13_6  (
            .in0(N__57935),
            .in1(N__58157),
            .in2(N__38078),
            .in3(N__40888),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIK8FN1_LC_14_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIK8FN1_LC_14_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIK8FN1_LC_14_14_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIK8FN1_LC_14_14_0  (
            .in0(N__55183),
            .in1(N__55387),
            .in2(N__35538),
            .in3(N__33730),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7EQL2_LC_14_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7EQL2_LC_14_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7EQL2_LC_14_14_1 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7EQL2_LC_14_14_1  (
            .in0(N__35537),
            .in1(N__54953),
            .in2(N__33737),
            .in3(N__54756),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRL7_LC_14_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRL7_LC_14_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRL7_LC_14_14_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRL7_LC_14_14_2  (
            .in0(N__53976),
            .in1(N__49669),
            .in2(N__30807),
            .in3(N__40791),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI2GCO7_LC_14_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI2GCO7_LC_14_14_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI2GCO7_LC_14_14_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI2GCO7_LC_14_14_3  (
            .in0(_gnd_net_),
            .in1(N__53670),
            .in2(N__30939),
            .in3(N__30936),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3_LC_14_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3_LC_14_14_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3_LC_14_14_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3_LC_14_14_4  (
            .in0(_gnd_net_),
            .in1(N__55584),
            .in2(N__30930),
            .in3(N__55650),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net ),
            .ce(N__55521),
            .sr(N__62884));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICQCO7_LC_14_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICQCO7_LC_14_14_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICQCO7_LC_14_14_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICQCO7_LC_14_14_5  (
            .in0(N__30927),
            .in1(N__53669),
            .in2(_gnd_net_),
            .in3(N__32139),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_5_LC_14_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_5_LC_14_14_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_5_LC_14_14_6 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_5_LC_14_14_6  (
            .in0(_gnd_net_),
            .in1(N__30891),
            .in2(N__30918),
            .in3(N__55652),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net ),
            .ce(N__55521),
            .sr(N__62884));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_4_LC_14_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_4_LC_14_14_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_4_LC_14_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_4_LC_14_14_7  (
            .in0(N__55651),
            .in1(N__30915),
            .in2(_gnd_net_),
            .in3(N__30909),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net ),
            .ce(N__55521),
            .sr(N__62884));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_9_LC_14_15_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_9_LC_14_15_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_9_LC_14_15_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_9_LC_14_15_0  (
            .in0(N__38301),
            .in1(N__37706),
            .in2(N__30879),
            .in3(N__46671),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_9_LC_14_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_9_LC_14_15_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_9_LC_14_15_1 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_9_LC_14_15_1  (
            .in0(N__33939),
            .in1(N__30878),
            .in2(N__59163),
            .in3(N__46461),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_21_LC_14_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_21_LC_14_15_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_21_LC_14_15_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_21_LC_14_15_2  (
            .in0(N__61436),
            .in1(N__59023),
            .in2(N__33365),
            .in3(N__33940),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_22_LC_14_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_22_LC_14_15_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_22_LC_14_15_3 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_22_LC_14_15_3  (
            .in0(N__33936),
            .in1(N__30866),
            .in2(N__59160),
            .in3(N__61319),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_23_LC_14_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_23_LC_14_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_23_LC_14_15_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_23_LC_14_15_4  (
            .in0(N__61253),
            .in1(N__59024),
            .in2(N__37934),
            .in3(N__33941),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_24_LC_14_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_24_LC_14_15_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_24_LC_14_15_5 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_24_LC_14_15_5  (
            .in0(N__33937),
            .in1(N__61131),
            .in2(N__59161),
            .in3(N__35264),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_25_LC_14_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_25_LC_14_15_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_25_LC_14_15_6 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_25_LC_14_15_6  (
            .in0(N__35198),
            .in1(N__59025),
            .in2(N__61020),
            .in3(N__33942),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_26_LC_14_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_26_LC_14_15_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_26_LC_14_15_7 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_26_LC_14_15_7  (
            .in0(N__33938),
            .in1(N__60913),
            .in2(N__59162),
            .in3(N__30962),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65585),
            .ce(N__32489),
            .sr(N__62876));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_0_LC_14_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_0_LC_14_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_0_LC_14_16_1 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_0_LC_14_16_1  (
            .in0(N__62479),
            .in1(N__36540),
            .in2(_gnd_net_),
            .in3(N__38674),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_LC_14_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_LC_14_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_LC_14_16_2 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_LC_14_16_2  (
            .in0(_gnd_net_),
            .in1(N__38726),
            .in2(N__30948),
            .in3(N__64157),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1959_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_tz_LC_14_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_tz_LC_14_16_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_tz_LC_14_16_3 .LUT_INIT=16'b1000111111001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_tz_LC_14_16_3  (
            .in0(N__36753),
            .in1(N__38699),
            .in2(N__30945),
            .in3(N__36807),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.rdata_tri_enable_LC_14_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.rdata_tri_enable_LC_14_16_4 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.rdata_tri_enable_LC_14_16_4 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.rdata_tri_enable_LC_14_16_4  (
            .in0(N__38821),
            .in1(_gnd_net_),
            .in2(N__30942),
            .in3(N__38904),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65597),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.rdata_tri_enable_LC_14_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.rdata_tri_enable_LC_14_16_5 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.rdata_tri_enable_LC_14_16_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.rdata_tri_enable_LC_14_16_5  (
            .in0(N__38903),
            .in1(N__38820),
            .in2(_gnd_net_),
            .in3(N__32311),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65597),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_2_LC_14_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_2_LC_14_17_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_2_LC_14_17_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_2_LC_14_17_0  (
            .in0(N__31605),
            .in1(N__34280),
            .in2(_gnd_net_),
            .in3(N__34148),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net ),
            .ce(),
            .sr(N__64970));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_8_LC_14_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_8_LC_14_17_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_8_LC_14_17_1 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_8_LC_14_17_1  (
            .in0(N__41424),
            .in1(N__36651),
            .in2(_gnd_net_),
            .in3(N__34421),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net ),
            .ce(),
            .sr(N__64970));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_o2_7_LC_14_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_o2_7_LC_14_17_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_o2_7_LC_14_17_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_o2_7_LC_14_17_2  (
            .in0(_gnd_net_),
            .in1(N__56246),
            .in2(_gnd_net_),
            .in3(N__38673),
            .lcout(N_1592_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_RNO_LC_14_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_RNO_LC_14_17_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_RNO_LC_14_17_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_RNO_LC_14_17_3  (
            .in0(N__39186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Control_StartUp_inst.N_8_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1EQD_LC_14_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1EQD_LC_14_17_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1EQD_LC_14_17_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1EQD_LC_14_17_4  (
            .in0(N__31200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_0_LC_14_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_0_LC_14_17_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_0_LC_14_17_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_0_LC_14_17_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30990),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_14_17_6.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_14_17_6.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_14_17_6.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_14_17_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19_LC_14_18_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19_LC_14_18_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19_LC_14_18_0 .LUT_INIT=16'b1010101000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19_LC_14_18_0  (
            .in0(N__31041),
            .in1(N__30978),
            .in2(_gnd_net_),
            .in3(N__31263),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net ),
            .ce(),
            .sr(N__62857));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_RNIBV54_LC_14_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_RNIBV54_LC_14_18_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_RNIBV54_LC_14_18_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_RNIBV54_LC_14_18_1  (
            .in0(_gnd_net_),
            .in1(N__32646),
            .in2(_gnd_net_),
            .in3(N__31051),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIFSQ8_17_LC_14_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIFSQ8_17_LC_14_18_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIFSQ8_17_LC_14_18_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIFSQ8_17_LC_14_18_2  (
            .in0(N__32666),
            .in1(N__32696),
            .in2(N__30972),
            .in3(N__32883),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_7_LC_14_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_7_LC_14_18_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_7_LC_14_18_3 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_7_LC_14_18_3  (
            .in0(N__31262),
            .in1(_gnd_net_),
            .in2(N__31125),
            .in3(N__31131),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net ),
            .ce(),
            .sr(N__62857));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIPCFF_19_LC_14_18_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIPCFF_19_LC_14_18_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIPCFF_19_LC_14_18_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIPCFF_19_LC_14_18_4  (
            .in0(N__31052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31119),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.en_count_bits_0_i_a2_0_a2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIO9811_11_LC_14_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIO9811_11_LC_14_18_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIO9811_11_LC_14_18_5 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIO9811_11_LC_14_18_5  (
            .in0(N__31027),
            .in1(N__31384),
            .in2(N__31101),
            .in3(N__31225),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_277_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_20_LC_14_18_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_20_LC_14_18_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_20_LC_14_18_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_20_LC_14_18_6  (
            .in0(N__31053),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31261),
            .lcout(\cemf_module_64ch_ctrl_inst1.end_conf_a ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net ),
            .ce(),
            .sr(N__62857));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_18_LC_14_18_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_18_LC_14_18_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_18_LC_14_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_18_LC_14_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32667),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net ),
            .ce(),
            .sr(N__62857));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_RNILJCF_LC_14_19_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_RNILJCF_LC_14_19_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_RNILJCF_LC_14_19_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_RNILJCF_LC_14_19_0  (
            .in0(N__31035),
            .in1(N__31218),
            .in2(N__31302),
            .in3(N__31280),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_LC_14_19_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_LC_14_19_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_LC_14_19_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_LC_14_19_1  (
            .in0(N__31281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_12_LC_14_19_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_12_LC_14_19_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_12_LC_14_19_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_12_LC_14_19_2  (
            .in0(_gnd_net_),
            .in1(N__31028),
            .in2(_gnd_net_),
            .in3(N__31258),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_15_LC_14_19_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_15_LC_14_19_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_15_LC_14_19_3 .LUT_INIT=16'b1101100011011101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_15_LC_14_19_3  (
            .in0(N__31259),
            .in1(N__31290),
            .in2(N__31227),
            .in3(N__31301),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_9_LC_14_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_9_LC_14_19_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_9_LC_14_19_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_9_LC_14_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32271),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_14_LC_14_19_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_14_LC_14_19_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_14_LC_14_19_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_14_LC_14_19_5  (
            .in0(N__32272),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_13_LC_14_19_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_13_LC_14_19_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_13_LC_14_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_13_LC_14_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31282),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_16_LC_14_19_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_16_LC_14_19_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_16_LC_14_19_7 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_16_LC_14_19_7  (
            .in0(N__31260),
            .in1(_gnd_net_),
            .in2(N__31226),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net ),
            .ce(),
            .sr(N__62850));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIK0RN1_16_LC_14_20_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIK0RN1_16_LC_14_20_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIK0RN1_16_LC_14_20_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIK0RN1_16_LC_14_20_0  (
            .in0(N__31171),
            .in1(N__32698),
            .in2(N__31185),
            .in3(N__31139),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_LC_14_20_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_LC_14_20_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_LC_14_20_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_LC_14_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31203),
            .in3(N__31191),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net ),
            .ce(),
            .sr(N__62846));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIIF971_13_LC_14_20_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIIF971_13_LC_14_20_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIIF971_13_LC_14_20_2 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIIF971_13_LC_14_20_2  (
            .in0(N__32673),
            .in1(N__32566),
            .in2(N__32276),
            .in3(N__32297),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_276_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_LC_14_20_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_LC_14_20_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_LC_14_20_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_LC_14_20_3  (
            .in0(N__31140),
            .in1(N__31184),
            .in2(N__32703),
            .in3(N__31172),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net ),
            .ce(),
            .sr(N__62846));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIEJSO_0_LC_14_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIEJSO_0_LC_14_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIEJSO_0_LC_14_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIEJSO_0_LC_14_20_4  (
            .in0(_gnd_net_),
            .in1(N__32592),
            .in2(_gnd_net_),
            .in3(N__36956),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_LC_14_20_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_LC_14_20_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_LC_14_20_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_LC_14_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31395),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net ),
            .ce(),
            .sr(N__62846));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_RNI7P0A1_LC_14_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_RNI7P0A1_LC_14_20_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_RNI7P0A1_LC_14_20_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_RNI7P0A1_LC_14_20_6  (
            .in0(N__31392),
            .in1(N__31383),
            .in2(N__31365),
            .in3(N__32591),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_LC_14_20_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_LC_14_20_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_LC_14_20_7 .LUT_INIT=16'b1111010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_LC_14_20_7  (
            .in0(N__36957),
            .in1(N__31350),
            .in2(N__31343),
            .in3(N__32904),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net ),
            .ce(),
            .sr(N__62846));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIMH2I_LC_14_21_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIMH2I_LC_14_21_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIMH2I_LC_14_21_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIMH2I_LC_14_21_0  (
            .in0(N__32950),
            .in1(N__37168),
            .in2(N__34551),
            .in3(N__35755),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNI6VG51_LC_14_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNI6VG51_LC_14_21_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNI6VG51_LC_14_21_1 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNI6VG51_LC_14_21_1  (
            .in0(_gnd_net_),
            .in1(N__32782),
            .in2(N__31320),
            .in3(N__32818),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43_0_LC_14_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43_0_LC_14_21_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43_0_LC_14_21_2 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43_0_LC_14_21_2  (
            .in0(N__36696),
            .in1(N__36868),
            .in2(N__31317),
            .in3(N__39743),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIS0GS_LC_14_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIS0GS_LC_14_21_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIS0GS_LC_14_21_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIS0GS_LC_14_21_3  (
            .in0(N__39742),
            .in1(N__32949),
            .in2(_gnd_net_),
            .in3(N__32817),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_10_LC_14_21_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_10_LC_14_21_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_10_LC_14_21_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_10_LC_14_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35796),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65657),
            .ce(),
            .sr(N__62839));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_RNIIDR41_LC_14_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_RNIIDR41_LC_14_21_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_RNIIDR41_LC_14_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_RNIIDR41_LC_14_21_5  (
            .in0(N__35756),
            .in1(N__34543),
            .in2(N__32718),
            .in3(N__36695),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_RNICL4J4_LC_14_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_RNICL4J4_LC_14_21_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_RNICL4J4_LC_14_21_6 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_RNICL4J4_LC_14_21_6  (
            .in0(N__36836),
            .in1(N__31551),
            .in2(N__31539),
            .in3(N__31536),
            .lcout(N_528_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_2_LC_14_22_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_2_LC_14_22_0 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_2_LC_14_22_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_2_LC_14_22_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31413),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65672),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_1_LC_14_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_1_LC_14_22_2 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_1_LC_14_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_1_LC_14_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31503),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65672),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_2_LC_14_22_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_2_LC_14_22_3 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_2_LC_14_22_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_2_LC_14_22_3  (
            .in0(N__31488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65672),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_RNI5H26_2_LC_14_22_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_RNI5H26_2_LC_14_22_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_RNI5H26_2_LC_14_22_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_RNI5H26_2_LC_14_22_4  (
            .in0(_gnd_net_),
            .in1(N__31494),
            .in2(_gnd_net_),
            .in3(N__31487),
            .lcout(\cemf_module_64ch_ctrl_inst1.n_state41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_li_0_i_i_a2_0_a2_1_LC_14_22_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_li_0_i_i_a2_0_a2_1_LC_14_22_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_li_0_i_i_a2_0_a2_1_LC_14_22_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_li_0_i_i_a2_0_a2_1_LC_14_22_5  (
            .in0(N__36904),
            .in1(N__32951),
            .in2(N__31457),
            .in3(N__34512),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_li_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_1_LC_14_22_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_1_LC_14_22_6 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_1_LC_14_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_1_LC_14_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50790),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65672),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0_LC_14_23_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0_LC_14_23_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0_LC_14_23_0 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0_LC_14_23_0  (
            .in0(N__34331),
            .in1(N__32540),
            .in2(N__63301),
            .in3(N__31407),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ),
            .ce(),
            .sr(N__64991));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_1_LC_14_23_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_1_LC_14_23_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_1_LC_14_23_1 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_1_LC_14_23_1  (
            .in0(N__32538),
            .in1(N__34332),
            .in2(N__63273),
            .in3(N__31401),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ),
            .ce(),
            .sr(N__64991));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_3_LC_14_23_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_3_LC_14_23_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_3_LC_14_23_2 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_3_LC_14_23_2  (
            .in0(N__34334),
            .in1(N__32541),
            .in2(N__63302),
            .in3(N__31617),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ),
            .ce(),
            .sr(N__64991));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_2_LC_14_23_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_2_LC_14_23_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_2_LC_14_23_3 .LUT_INIT=16'b1111011100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_2_LC_14_23_3  (
            .in0(N__32539),
            .in1(N__34333),
            .in2(N__63274),
            .in3(N__31611),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ),
            .ce(),
            .sr(N__64991));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIH7DQ_3_LC_14_23_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIH7DQ_3_LC_14_23_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIH7DQ_3_LC_14_23_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIH7DQ_3_LC_14_23_4  (
            .in0(N__34216),
            .in1(N__34240),
            .in2(_gnd_net_),
            .in3(N__34189),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_275_0 ),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_275_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNI7FJ71_0_LC_14_23_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNI7FJ71_0_LC_14_23_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNI7FJ71_0_LC_14_23_5 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNI7FJ71_0_LC_14_23_5  (
            .in0(N__34116),
            .in1(_gnd_net_),
            .in2(N__31596),
            .in3(N__34276),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_1_LC_14_23_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_1_LC_14_23_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_1_LC_14_23_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_1_LC_14_23_6  (
            .in0(N__34335),
            .in1(N__63231),
            .in2(N__31593),
            .in3(N__36573),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net ),
            .ce(),
            .sr(N__64991));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI344J1_1_LC_14_23_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI344J1_1_LC_14_23_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI344J1_1_LC_14_23_7 .LUT_INIT=16'b1111101111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI344J1_1_LC_14_23_7  (
            .in0(N__63230),
            .in1(N__34330),
            .in2(N__34125),
            .in3(N__34299),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_13_LC_14_24_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_13_LC_14_24_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_13_LC_14_24_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_13_LC_14_24_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37116),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65696),
            .ce(),
            .sr(N__62823));
    defparam \serializer_mod_inst.current_state_1_LC_14_26_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_1_LC_14_26_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.current_state_1_LC_14_26_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \serializer_mod_inst.current_state_1_LC_14_26_7  (
            .in0(_gnd_net_),
            .in1(N__45174),
            .in2(_gnd_net_),
            .in3(N__45064),
            .lcout(\serializer_mod_inst.current_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65724),
            .ce(),
            .sr(N__62813));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_2_LC_15_7_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_2_LC_15_7_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_2_LC_15_7_1 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_2_LC_15_7_1  (
            .in0(N__33087),
            .in1(N__31575),
            .in2(N__51926),
            .in3(N__49752),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_2_LC_15_8_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_2_LC_15_8_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_2_LC_15_8_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_2_LC_15_8_1  (
            .in0(N__31569),
            .in1(N__52769),
            .in2(N__31764),
            .in3(N__52513),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_2_LC_15_8_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_2_LC_15_8_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_2_LC_15_8_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_2_LC_15_8_2  (
            .in0(_gnd_net_),
            .in1(N__52204),
            .in2(N__31746),
            .in3(N__43005),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_2_LC_15_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_2_LC_15_8_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_2_LC_15_8_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_2_LC_15_8_3  (
            .in0(N__35280),
            .in1(N__33297),
            .in2(N__31743),
            .in3(N__31740),
            .lcout(I2C_top_level_inst1_s_data_oreg_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65514),
            .ce(N__54515),
            .sr(N__65002));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_10_LC_15_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_10_LC_15_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_10_LC_15_9_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_10_LC_15_9_0  (
            .in0(N__31734),
            .in1(N__52674),
            .in2(N__31716),
            .in3(N__52494),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_10_LC_15_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_10_LC_15_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_10_LC_15_9_1 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_10_LC_15_9_1  (
            .in0(N__42738),
            .in1(_gnd_net_),
            .in2(N__31698),
            .in3(N__52123),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_10_LC_15_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_10_LC_15_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_10_LC_15_9_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_10_LC_15_9_2  (
            .in0(N__44640),
            .in1(N__31695),
            .in2(N__61712),
            .in3(N__44414),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_10_LC_15_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_10_LC_15_9_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_10_LC_15_9_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_10_LC_15_9_3  (
            .in0(N__31677),
            .in1(N__51791),
            .in2(N__31668),
            .in3(N__49307),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_10_LC_15_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_10_LC_15_9_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_10_LC_15_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_10_LC_15_9_4  (
            .in0(N__31665),
            .in1(N__37890),
            .in2(N__31653),
            .in3(N__31650),
            .lcout(I2C_top_level_inst1_s_data_oreg_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65519),
            .ce(N__54512),
            .sr(N__64998));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_18_LC_15_9_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_18_LC_15_9_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_18_LC_15_9_5 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_18_LC_15_9_5  (
            .in0(N__52495),
            .in1(N__31644),
            .in2(N__58766),
            .in3(N__44639),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_11_LC_15_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_11_LC_15_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_11_LC_15_10_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_11_LC_15_10_0  (
            .in0(N__31935),
            .in1(N__52673),
            .in2(N__31914),
            .in3(N__52493),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_11_LC_15_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_11_LC_15_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_11_LC_15_10_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_11_LC_15_10_1  (
            .in0(_gnd_net_),
            .in1(N__52122),
            .in2(N__31893),
            .in3(N__42915),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_11_LC_15_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_11_LC_15_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_11_LC_15_10_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_11_LC_15_10_2  (
            .in0(N__44409),
            .in1(N__63905),
            .in2(N__44660),
            .in3(N__31890),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_11_LC_15_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_11_LC_15_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_11_LC_15_10_3 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_11_LC_15_10_3  (
            .in0(N__51790),
            .in1(N__31872),
            .in2(N__31857),
            .in3(N__42558),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_11_LC_15_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_11_LC_15_10_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_11_LC_15_10_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_11_LC_15_10_4  (
            .in0(N__31854),
            .in1(N__31848),
            .in2(N__31842),
            .in3(N__35079),
            .lcout(I2C_top_level_inst1_s_data_oreg_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65523),
            .ce(N__54508),
            .sr(N__64993));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_19_LC_15_10_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_19_LC_15_10_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_19_LC_15_10_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_19_LC_15_10_5  (
            .in0(N__31839),
            .in1(N__44628),
            .in2(N__58634),
            .in3(N__44408),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_20_LC_15_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_20_LC_15_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_20_LC_15_11_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_20_LC_15_11_0  (
            .in0(N__31821),
            .in1(N__52676),
            .in2(N__31803),
            .in3(N__52381),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_20_LC_15_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_20_LC_15_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_20_LC_15_11_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_20_LC_15_11_1  (
            .in0(_gnd_net_),
            .in1(N__52124),
            .in2(N__31785),
            .in3(N__35691),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_20_LC_15_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_20_LC_15_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_20_LC_15_11_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_20_LC_15_11_2  (
            .in0(N__31782),
            .in1(N__38374),
            .in2(N__58593),
            .in3(N__44664),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_20_LC_15_11_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_20_LC_15_11_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_20_LC_15_11_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_20_LC_15_11_3  (
            .in0(N__32028),
            .in1(N__38278),
            .in2(N__32013),
            .in3(N__42423),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_20_LC_15_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_20_LC_15_11_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_20_LC_15_11_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_20_LC_15_11_4  (
            .in0(N__38034),
            .in1(N__33465),
            .in2(N__32010),
            .in3(N__32007),
            .lcout(I2C_top_level_inst1_s_data_oreg_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65530),
            .ce(N__54504),
            .sr(N__64988));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQEFN1_LC_15_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQEFN1_LC_15_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQEFN1_LC_15_12_0 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQEFN1_LC_15_12_0  (
            .in0(N__33673),
            .in1(N__55217),
            .in2(N__41088),
            .in3(N__55431),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIDKQL2_LC_15_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIDKQL2_LC_15_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIDKQL2_LC_15_12_1 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIDKQL2_LC_15_12_1  (
            .in0(N__55001),
            .in1(N__33674),
            .in2(N__54836),
            .in3(N__41087),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRL7_LC_15_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRL7_LC_15_12_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRL7_LC_15_12_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRL7_LC_15_12_2  (
            .in0(N__53949),
            .in1(N__31981),
            .in2(N__31965),
            .in3(N__33747),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRLZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SL7_LC_15_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SL7_LC_15_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SL7_LC_15_12_3 .LUT_INIT=16'b0011101111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SL7_LC_15_12_3  (
            .in0(N__40510),
            .in1(N__45513),
            .in2(N__53994),
            .in3(N__40560),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIM4DO7_LC_15_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIM4DO7_LC_15_12_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIM4DO7_LC_15_12_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIM4DO7_LC_15_12_4  (
            .in0(N__32058),
            .in1(_gnd_net_),
            .in2(N__31962),
            .in3(N__53695),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHVCO7_LC_15_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHVCO7_LC_15_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHVCO7_LC_15_12_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHVCO7_LC_15_12_5  (
            .in0(N__53694),
            .in1(N__31953),
            .in2(_gnd_net_),
            .in3(N__31959),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6_LC_15_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6_LC_15_12_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6_LC_15_12_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6_LC_15_12_6  (
            .in0(N__31947),
            .in1(_gnd_net_),
            .in2(N__31938),
            .in3(N__55693),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net ),
            .ce(N__55522),
            .sr(N__62895));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_7_LC_15_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_7_LC_15_12_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_7_LC_15_12_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_7_LC_15_12_7  (
            .in0(N__55694),
            .in1(N__32064),
            .in2(_gnd_net_),
            .in3(N__32057),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net ),
            .ce(N__55522),
            .sr(N__62895));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_6_LC_15_13_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_6_LC_15_13_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_6_LC_15_13_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_6_LC_15_13_0  (
            .in0(N__38269),
            .in1(N__37694),
            .in2(N__32040),
            .in3(N__41083),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_6_LC_15_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_6_LC_15_13_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_6_LC_15_13_1 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_6_LC_15_13_1  (
            .in0(N__33946),
            .in1(N__32039),
            .in2(N__59544),
            .in3(N__63543),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_16_LC_15_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_16_LC_15_13_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_16_LC_15_13_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_16_LC_15_13_2  (
            .in0(N__57632),
            .in1(N__59333),
            .in2(N__34910),
            .in3(N__33947),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_17_LC_15_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_17_LC_15_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_17_LC_15_13_3 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_17_LC_15_13_3  (
            .in0(N__33943),
            .in1(N__35330),
            .in2(N__59541),
            .in3(N__57423),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_18_LC_15_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_18_LC_15_13_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_18_LC_15_13_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_18_LC_15_13_4  (
            .in0(N__59850),
            .in1(N__59334),
            .in2(N__33521),
            .in3(N__33948),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_19_LC_15_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_19_LC_15_13_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_19_LC_15_13_5 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_19_LC_15_13_5  (
            .in0(N__33944),
            .in1(N__35234),
            .in2(N__59542),
            .in3(N__61639),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_2_LC_15_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_2_LC_15_13_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_2_LC_15_13_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_2_LC_15_13_6  (
            .in0(N__61711),
            .in1(N__59335),
            .in2(N__35303),
            .in3(N__33949),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_20_LC_15_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_20_LC_15_13_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_20_LC_15_13_7 .LUT_INIT=16'b0100111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_20_LC_15_13_7  (
            .in0(N__33945),
            .in1(N__33479),
            .in2(N__59543),
            .in3(N__61526),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65550),
            .ce(N__32512),
            .sr(N__62885));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2HK93_LC_15_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2HK93_LC_15_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2HK93_LC_15_14_1 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2HK93_LC_15_14_1  (
            .in0(N__45842),
            .in1(N__46013),
            .in2(N__32208),
            .in3(N__42212),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRL7_LC_15_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRL7_LC_15_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRL7_LC_15_14_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRL7_LC_15_14_2  (
            .in0(N__53969),
            .in1(N__32170),
            .in2(N__32142),
            .in3(N__32133),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRLZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBIQL2_LC_15_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBIQL2_LC_15_14_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBIQL2_LC_15_14_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBIQL2_LC_15_14_3  (
            .in0(N__54928),
            .in1(N__54736),
            .in2(N__41126),
            .in3(N__32110),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_5_LC_15_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_5_LC_15_14_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_5_LC_15_14_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_5_LC_15_14_4  (
            .in0(_gnd_net_),
            .in1(N__63677),
            .in2(_gnd_net_),
            .in3(N__59141),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65562),
            .ce(N__49059),
            .sr(N__62877));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOOQI1_LC_15_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOOQI1_LC_15_14_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOOQI1_LC_15_14_5 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOOQI1_LC_15_14_5  (
            .in0(N__55154),
            .in1(N__55386),
            .in2(N__42644),
            .in3(N__32080),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_14_LC_15_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_14_LC_15_14_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_14_LC_15_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_14_LC_15_14_6  (
            .in0(_gnd_net_),
            .in1(N__58496),
            .in2(_gnd_net_),
            .in3(N__59140),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65562),
            .ce(N__49059),
            .sr(N__62877));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBU5H2_LC_15_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBU5H2_LC_15_14_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBU5H2_LC_15_14_7 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBU5H2_LC_15_14_7  (
            .in0(N__54929),
            .in1(N__54735),
            .in2(N__42645),
            .in3(N__32081),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_7_LC_15_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_7_LC_15_15_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_7_LC_15_15_0 .LUT_INIT=16'b1000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_7_LC_15_15_0  (
            .in0(N__34092),
            .in1(N__50449),
            .in2(N__63472),
            .in3(N__33798),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65575),
            .ce(N__32488),
            .sr(N__62870));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_m2_0_LC_15_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_m2_0_LC_15_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_m2_0_LC_15_15_1 .LUT_INIT=16'b0111000011111000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_m2_0_LC_15_15_1  (
            .in0(N__36306),
            .in1(N__34844),
            .in2(N__34671),
            .in3(N__38665),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_242_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_i_0_LC_15_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_i_0_LC_15_15_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_i_0_LC_15_15_2 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_i_0_LC_15_15_2  (
            .in0(N__38706),
            .in1(N__34670),
            .in2(N__32067),
            .in3(N__62481),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_1_LC_15_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_1_LC_15_15_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_1_LC_15_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_1_LC_15_15_3  (
            .in0(_gnd_net_),
            .in1(N__61863),
            .in2(_gnd_net_),
            .in3(N__34091),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65575),
            .ce(N__32488),
            .sr(N__62870));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_0_a2_0_LC_15_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_0_a2_0_LC_15_15_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_0_a2_0_LC_15_15_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_0_a2_0_LC_15_15_5  (
            .in0(N__36272),
            .in1(N__34843),
            .in2(_gnd_net_),
            .in3(N__38664),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_15_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_15_15_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_15_15_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_15_15_6  (
            .in0(N__38666),
            .in1(N__34851),
            .in2(_gnd_net_),
            .in3(N__36324),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_27_LC_15_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_27_LC_15_15_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_27_LC_15_15_7 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_27_LC_15_15_7  (
            .in0(N__35177),
            .in1(N__59139),
            .in2(N__60816),
            .in3(N__33922),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65575),
            .ce(N__32488),
            .sr(N__62870));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_5_LC_15_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_5_LC_15_16_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_5_LC_15_16_1 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_5_LC_15_16_1  (
            .in0(N__33919),
            .in1(N__32222),
            .in2(N__63697),
            .in3(N__59016),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_10_LC_15_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_10_LC_15_16_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_10_LC_15_16_2 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_10_LC_15_16_2  (
            .in0(N__58783),
            .in1(N__37904),
            .in2(N__33950),
            .in3(N__59012),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_11_LC_15_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_11_LC_15_16_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_11_LC_15_16_3 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_11_LC_15_16_3  (
            .in0(N__33916),
            .in1(N__58660),
            .in2(N__35099),
            .in3(N__59013),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_12_LC_15_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_12_LC_15_16_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_12_LC_15_16_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_12_LC_15_16_4  (
            .in0(N__58596),
            .in1(N__59010),
            .in2(N__35060),
            .in3(N__33920),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_13_LC_15_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_13_LC_15_16_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_13_LC_15_16_5 .LUT_INIT=16'b0100010011100100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_13_LC_15_16_5  (
            .in0(N__33917),
            .in1(N__35018),
            .in2(N__58357),
            .in3(N__59014),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_14_LC_15_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_14_LC_15_16_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_14_LC_15_16_6 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_14_LC_15_16_6  (
            .in0(N__58500),
            .in1(N__59011),
            .in2(N__34988),
            .in3(N__33921),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_15_LC_15_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_15_LC_15_16_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_15_LC_15_16_7 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_15_LC_15_16_7  (
            .in0(N__33918),
            .in1(N__57520),
            .in2(N__34943),
            .in3(N__59015),
            .lcout(cemf_module_64ch_ctrl_inst1_s_data_system_o_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65586),
            .ce(N__32490),
            .sr(N__62862));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_16_LC_15_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_16_LC_15_17_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_16_LC_15_17_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_16_LC_15_17_1  (
            .in0(N__64071),
            .in1(N__32451),
            .in2(N__43431),
            .in3(N__37803),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_764 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_18_LC_15_17_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_18_LC_15_17_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_18_LC_15_17_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_18_LC_15_17_2  (
            .in0(N__32336),
            .in1(N__43370),
            .in2(N__32433),
            .in3(N__64072),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1911 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_0_LC_15_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_0_LC_15_17_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_0_LC_15_17_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_0_LC_15_17_3  (
            .in0(_gnd_net_),
            .in1(N__66799),
            .in2(_gnd_net_),
            .in3(N__57238),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_8_LC_15_17_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_8_LC_15_17_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_8_LC_15_17_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_8_LC_15_17_4  (
            .in0(N__32337),
            .in1(N__32400),
            .in2(N__32385),
            .in3(N__64070),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1920 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.rdata_tri_enable_LC_15_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.rdata_tri_enable_LC_15_17_5 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.rdata_tri_enable_LC_15_17_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.rdata_tri_enable_LC_15_17_5  (
            .in0(N__38893),
            .in1(N__38808),
            .in2(_gnd_net_),
            .in3(N__32313),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65598),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.rdata_tri_enable_LC_15_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.rdata_tri_enable_LC_15_17_7 .SEQ_MODE=4'b1000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.rdata_tri_enable_LC_15_17_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.rdata_tri_enable_LC_15_17_7  (
            .in0(N__38892),
            .in1(N__38807),
            .in2(_gnd_net_),
            .in3(N__32312),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65598),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_LC_15_18_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_LC_15_18_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_LC_15_18_0 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_LC_15_18_0  (
            .in0(N__32557),
            .in1(N__32298),
            .in2(N__32277),
            .in3(N__32671),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net ),
            .ce(),
            .sr(N__62851));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_17_LC_15_18_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_17_LC_15_18_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_17_LC_15_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_17_LC_15_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32702),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net ),
            .ce(),
            .sr(N__62851));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_LC_15_18_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_LC_15_18_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_LC_15_18_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_LC_15_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32672),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net ),
            .ce(),
            .sr(N__62851));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_1_LC_15_18_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_1_LC_15_18_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_1_LC_15_18_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_1_LC_15_18_3  (
            .in0(N__32602),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36967),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net ),
            .ce(),
            .sr(N__62851));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_RNIETUR_1_LC_15_18_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_RNIETUR_1_LC_15_18_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_RNIETUR_1_LC_15_18_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_RNIETUR_1_LC_15_18_4  (
            .in0(N__36477),
            .in1(N__36435),
            .in2(_gnd_net_),
            .in3(N__66274),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1372_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI216D_2_LC_15_18_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI216D_2_LC_15_18_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI216D_2_LC_15_18_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI216D_2_LC_15_18_5  (
            .in0(N__43813),
            .in1(N__36595),
            .in2(_gnd_net_),
            .in3(N__34420),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1379_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI2QEM_0_LC_15_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI2QEM_0_LC_15_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI2QEM_0_LC_15_18_6 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI2QEM_0_LC_15_18_6  (
            .in0(N__50881),
            .in1(N__43671),
            .in2(_gnd_net_),
            .in3(N__34170),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_113_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI35U51_14_LC_15_18_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI35U51_14_LC_15_18_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI35U51_14_LC_15_18_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI35U51_14_LC_15_18_7  (
            .in0(N__34147),
            .in1(N__34359),
            .in2(_gnd_net_),
            .in3(N__34295),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_11_0_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_14_LC_15_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_14_LC_15_19_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_14_LC_15_19_0 .LUT_INIT=16'b0100010111001111;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_14_LC_15_19_0  (
            .in0(N__32751),
            .in1(N__50865),
            .in2(N__34358),
            .in3(N__43931),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_12_LC_15_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_12_LC_15_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_12_LC_15_19_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_12_LC_15_19_1  (
            .in0(N__43902),
            .in1(N__48256),
            .in2(_gnd_net_),
            .in3(N__36676),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1394_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_12_LC_15_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_12_LC_15_19_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_12_LC_15_19_2 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_12_LC_15_19_2  (
            .in0(N__36638),
            .in1(N__63197),
            .in2(N__32520),
            .in3(N__32727),
            .lcout(\I2C_top_level_inst1.s_enable_desp_tx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net ),
            .ce(),
            .sr(N__64980));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_12_LC_15_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_12_LC_15_19_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_12_LC_15_19_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_12_LC_15_19_3  (
            .in0(N__43932),
            .in1(N__32750),
            .in2(_gnd_net_),
            .in3(N__34375),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_13_LC_15_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_13_LC_15_19_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_13_LC_15_19_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_13_LC_15_19_4  (
            .in0(N__36639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63198),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net ),
            .ce(),
            .sr(N__64980));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_LC_15_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_LC_15_19_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_LC_15_19_5 .LUT_INIT=16'b1111110010001100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_LC_15_19_5  (
            .in0(N__50864),
            .in1(N__34354),
            .in2(N__43686),
            .in3(N__36677),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net ),
            .ce(),
            .sr(N__64980));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_4_LC_15_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_4_LC_15_19_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_4_LC_15_19_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_4_LC_15_19_6  (
            .in0(N__36675),
            .in1(N__43903),
            .in2(_gnd_net_),
            .in3(N__48257),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1381_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_4_LC_15_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_4_LC_15_19_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_4_LC_15_19_7 .LUT_INIT=16'b1011101110110000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_4_LC_15_19_7  (
            .in0(N__43904),
            .in1(N__36640),
            .in2(N__32721),
            .in3(N__36599),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net ),
            .ce(),
            .sr(N__64980));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO59R_2_LC_15_20_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO59R_2_LC_15_20_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO59R_2_LC_15_20_0 .LUT_INIT=16'b0000000000100011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO59R_2_LC_15_20_0  (
            .in0(N__32899),
            .in1(N__36958),
            .in2(N__32862),
            .in3(N__35725),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_LC_15_20_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_LC_15_20_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_LC_15_20_1 .LUT_INIT=16'b0000001100000001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_LC_15_20_1  (
            .in0(N__32857),
            .in1(N__35748),
            .in2(N__36968),
            .in3(N__32903),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65631),
            .ce(),
            .sr(N__62840));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_4_LC_15_20_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_4_LC_15_20_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_4_LC_15_20_2 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_4_LC_15_20_2  (
            .in0(N__32902),
            .in1(N__36960),
            .in2(_gnd_net_),
            .in3(N__32858),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_state_i_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65631),
            .ce(),
            .sr(N__62840));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_3_LC_15_20_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_3_LC_15_20_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_3_LC_15_20_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_3_LC_15_20_3  (
            .in0(_gnd_net_),
            .in1(N__32709),
            .in2(_gnd_net_),
            .in3(N__32901),
            .lcout(\cemf_module_64ch_ctrl_inst1.start_conf_b ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65631),
            .ce(),
            .sr(N__62840));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNI2QTM_20_LC_15_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNI2QTM_20_LC_15_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNI2QTM_20_LC_15_20_4 .LUT_INIT=16'b0010001000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNI2QTM_20_LC_15_20_4  (
            .in0(N__32900),
            .in1(N__36959),
            .in2(_gnd_net_),
            .in3(N__32856),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_1817_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_2_LC_15_20_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_2_LC_15_20_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_2_LC_15_20_5 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_2_LC_15_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32865),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65631),
            .ce(),
            .sr(N__62840));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIM2JK_2_LC_15_20_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIM2JK_2_LC_15_20_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIM2JK_2_LC_15_20_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIM2JK_2_LC_15_20_6  (
            .in0(_gnd_net_),
            .in1(N__35818),
            .in2(_gnd_net_),
            .in3(N__32855),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_4_LC_15_20_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_4_LC_15_20_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_4_LC_15_20_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_4_LC_15_20_7  (
            .in0(N__35819),
            .in1(N__35881),
            .in2(_gnd_net_),
            .in3(N__32993),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65631),
            .ce(),
            .sr(N__62840));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_RNI3S391_LC_15_21_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_RNI3S391_LC_15_21_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_RNI3S391_LC_15_21_0 .LUT_INIT=16'b0000001100000111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_RNI3S391_LC_15_21_0  (
            .in0(N__32838),
            .in1(N__36955),
            .in2(N__32826),
            .in3(N__37083),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1874_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNISDQ71_10_LC_15_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNISDQ71_10_LC_15_21_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNISDQ71_10_LC_15_21_1 .LUT_INIT=16'b0101000001110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNISDQ71_10_LC_15_21_1  (
            .in0(N__36954),
            .in1(N__37161),
            .in2(N__36909),
            .in3(N__36717),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1873_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIP3H21_LC_15_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIP3H21_LC_15_21_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIP3H21_LC_15_21_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIP3H21_LC_15_21_2  (
            .in0(N__36837),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32783),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_RNIAUPM2_LC_15_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_RNIAUPM2_LC_15_21_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_RNIAUPM2_LC_15_21_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_RNIAUPM2_LC_15_21_3  (
            .in0(N__37082),
            .in1(N__34521),
            .in2(N__32799),
            .in3(N__32796),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1950 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIVHBV1_LC_15_21_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIVHBV1_LC_15_21_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIVHBV1_LC_15_21_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIVHBV1_LC_15_21_4  (
            .in0(N__32790),
            .in1(N__32784),
            .in2(_gnd_net_),
            .in3(N__34511),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIUA133_LC_15_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIUA133_LC_15_21_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIUA133_LC_15_21_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIUA133_LC_15_21_5  (
            .in0(N__39757),
            .in1(N__32952),
            .in2(N__33027),
            .in3(N__36900),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1949_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNII03U6_LC_15_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNII03U6_LC_15_21_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNII03U6_LC_15_21_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNII03U6_LC_15_21_6  (
            .in0(N__34599),
            .in1(N__33024),
            .in2(N__33018),
            .in3(N__35400),
            .lcout(stop_fpga2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_5_LC_15_22_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_5_LC_15_22_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_5_LC_15_22_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_5_LC_15_22_0  (
            .in0(_gnd_net_),
            .in1(N__35888),
            .in2(_gnd_net_),
            .in3(N__32997),
            .lcout(\cemf_module_64ch_ctrl_inst1.clr_sys_reg ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_1_LC_15_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_1_LC_15_22_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_1_LC_15_22_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_1_LC_15_22_1  (
            .in0(_gnd_net_),
            .in1(N__34629),
            .in2(_gnd_net_),
            .in3(N__35396),
            .lcout(\cemf_module_64ch_ctrl_inst1.start_conf_a ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_LC_15_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_LC_15_22_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_LC_15_22_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_LC_15_22_2  (
            .in0(N__35367),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35922),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \serializer_mod_inst.shift_reg_55_LC_15_22_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_55_LC_15_22_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_55_LC_15_22_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_55_LC_15_22_4  (
            .in0(N__47883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40122),
            .lcout(\serializer_mod_inst.shift_regZ0Z_55 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \serializer_mod_inst.shift_reg_113_LC_15_22_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_113_LC_15_22_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_113_LC_15_22_5 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_113_LC_15_22_5  (
            .in0(N__32931),
            .in1(N__45389),
            .in2(_gnd_net_),
            .in3(N__44901),
            .lcout(\serializer_mod_inst.shift_regZ0Z_113 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_0_LC_15_22_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_0_LC_15_22_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_0_LC_15_22_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_0_LC_15_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34494),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \serializer_mod_inst.shift_reg_112_LC_15_22_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_112_LC_15_22_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_112_LC_15_22_7 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_112_LC_15_22_7  (
            .in0(N__33060),
            .in1(N__45388),
            .in2(_gnd_net_),
            .in3(N__44900),
            .lcout(\serializer_mod_inst.shift_regZ0Z_112 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65658),
            .ce(),
            .sr(N__62830));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_2_LC_15_23_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_2_LC_15_23_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_2_LC_15_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_2_LC_15_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48105),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65673),
            .ce(N__44088),
            .sr(N__64997));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_4_LC_15_23_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_4_LC_15_23_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_4_LC_15_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_4_LC_15_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41376),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65673),
            .ce(N__44088),
            .sr(N__64997));
    defparam \serializer_mod_inst.shift_reg_111_LC_15_24_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_111_LC_15_24_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_111_LC_15_24_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_111_LC_15_24_0  (
            .in0(N__47879),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34740),
            .lcout(\serializer_mod_inst.shift_regZ0Z_111 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65682),
            .ce(),
            .sr(N__62818));
    defparam \serializer_mod_inst.shift_reg_119_LC_15_24_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_119_LC_15_24_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_119_LC_15_24_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_119_LC_15_24_1  (
            .in0(_gnd_net_),
            .in1(N__33033),
            .in2(_gnd_net_),
            .in3(N__47880),
            .lcout(\serializer_mod_inst.shift_regZ0Z_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65682),
            .ce(),
            .sr(N__62818));
    defparam \serializer_mod_inst.shift_reg_39_LC_15_24_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_39_LC_15_24_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_39_LC_15_24_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_39_LC_15_24_2  (
            .in0(N__47882),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33183),
            .lcout(\serializer_mod_inst.shift_regZ0Z_39 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65682),
            .ce(),
            .sr(N__62818));
    defparam \serializer_mod_inst.shift_reg_121_LC_15_24_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_121_LC_15_24_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_121_LC_15_24_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_121_LC_15_24_5  (
            .in0(_gnd_net_),
            .in1(N__33045),
            .in2(_gnd_net_),
            .in3(N__47881),
            .lcout(\serializer_mod_inst.shift_regZ0Z_121 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65682),
            .ce(),
            .sr(N__62818));
    defparam \serializer_mod_inst.shift_reg_120_LC_15_24_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_120_LC_15_24_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_120_LC_15_24_7 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_120_LC_15_24_7  (
            .in0(N__44964),
            .in1(N__33051),
            .in2(_gnd_net_),
            .in3(N__45247),
            .lcout(\serializer_mod_inst.shift_regZ0Z_120 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65682),
            .ce(),
            .sr(N__62818));
    defparam \serializer_mod_inst.shift_reg_36_LC_15_25_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_36_LC_15_25_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_36_LC_15_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_36_LC_15_25_0  (
            .in0(N__47878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33165),
            .lcout(\serializer_mod_inst.shift_regZ0Z_36 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65697),
            .ce(),
            .sr(N__62814));
    defparam \serializer_mod_inst.shift_reg_37_LC_15_25_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_37_LC_15_25_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_37_LC_15_25_4 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_37_LC_15_25_4  (
            .in0(N__45031),
            .in1(N__33039),
            .in2(_gnd_net_),
            .in3(N__45177),
            .lcout(\serializer_mod_inst.shift_regZ0Z_37 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65697),
            .ce(),
            .sr(N__62814));
    defparam \serializer_mod_inst.shift_reg_118_LC_15_25_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_118_LC_15_25_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_118_LC_15_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_118_LC_15_25_5  (
            .in0(_gnd_net_),
            .in1(N__34863),
            .in2(_gnd_net_),
            .in3(N__47877),
            .lcout(\serializer_mod_inst.shift_regZ0Z_118 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65697),
            .ce(),
            .sr(N__62814));
    defparam \serializer_mod_inst.shift_reg_33_LC_15_25_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_33_LC_15_25_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_33_LC_15_25_6 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_33_LC_15_25_6  (
            .in0(N__45030),
            .in1(N__34563),
            .in2(_gnd_net_),
            .in3(N__45176),
            .lcout(\serializer_mod_inst.shift_regZ0Z_33 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65697),
            .ce(),
            .sr(N__62814));
    defparam \serializer_mod_inst.shift_reg_38_LC_15_25_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_38_LC_15_25_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_38_LC_15_25_7 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_38_LC_15_25_7  (
            .in0(N__45178),
            .in1(N__33189),
            .in2(_gnd_net_),
            .in3(N__45032),
            .lcout(\serializer_mod_inst.shift_regZ0Z_38 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65697),
            .ce(),
            .sr(N__62814));
    defparam \serializer_mod_inst.shift_reg_76_LC_15_26_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_76_LC_15_26_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_76_LC_15_26_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_76_LC_15_26_0  (
            .in0(N__47870),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40245),
            .lcout(\serializer_mod_inst.shift_regZ0Z_76 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65715),
            .ce(),
            .sr(N__62810));
    defparam \serializer_mod_inst.shift_reg_34_LC_15_26_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_34_LC_15_26_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_34_LC_15_26_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_34_LC_15_26_1  (
            .in0(N__33177),
            .in1(N__45175),
            .in2(_gnd_net_),
            .in3(N__45057),
            .lcout(\serializer_mod_inst.shift_regZ0Z_34 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65715),
            .ce(),
            .sr(N__62810));
    defparam \serializer_mod_inst.shift_reg_35_LC_15_26_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_35_LC_15_26_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_35_LC_15_26_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_35_LC_15_26_5  (
            .in0(_gnd_net_),
            .in1(N__33171),
            .in2(_gnd_net_),
            .in3(N__47869),
            .lcout(\serializer_mod_inst.shift_regZ0Z_35 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65715),
            .ce(),
            .sr(N__62810));
    defparam \serializer_mod_inst.shift_reg_77_LC_15_26_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_77_LC_15_26_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_77_LC_15_26_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_77_LC_15_26_7  (
            .in0(_gnd_net_),
            .in1(N__33159),
            .in2(_gnd_net_),
            .in3(N__47871),
            .lcout(\serializer_mod_inst.shift_regZ0Z_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65715),
            .ce(),
            .sr(N__62810));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_17_LC_16_8_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_17_LC_16_8_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_17_LC_16_8_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_17_LC_16_8_0  (
            .in0(N__64246),
            .in1(N__33153),
            .in2(N__43572),
            .in3(N__37878),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_753 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_19_LC_16_8_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_19_LC_16_8_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_19_LC_16_8_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_19_LC_16_8_1  (
            .in0(N__37879),
            .in1(N__43529),
            .in2(N__33123),
            .in3(N__64249),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_731 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_2_LC_16_8_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_2_LC_16_8_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_2_LC_16_8_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_2_LC_16_8_2  (
            .in0(N__64248),
            .in1(N__33102),
            .in2(N__43574),
            .in3(N__37877),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_918 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_22_LC_16_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_22_LC_16_8_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_22_LC_16_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_22_LC_16_8_3  (
            .in0(N__37874),
            .in1(N__43519),
            .in2(N__33345),
            .in3(N__64245),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_698 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_23_LC_16_8_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_23_LC_16_8_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_23_LC_16_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_23_LC_16_8_4  (
            .in0(N__64247),
            .in1(N__33312),
            .in2(N__43573),
            .in3(N__37880),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_687 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_2_LC_16_8_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_2_LC_16_8_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_2_LC_16_8_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_2_LC_16_8_5  (
            .in0(N__52983),
            .in1(N__53792),
            .in2(N__53318),
            .in3(N__49965),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_25_LC_16_8_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_25_LC_16_8_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_25_LC_16_8_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_25_LC_16_8_6  (
            .in0(N__64243),
            .in1(N__33291),
            .in2(N__43571),
            .in3(N__37875),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_665 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_27_LC_16_8_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_27_LC_16_8_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_27_LC_16_8_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_27_LC_16_8_7  (
            .in0(N__37876),
            .in1(N__43518),
            .in2(N__33273),
            .in3(N__64244),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_654 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_19_LC_16_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_19_LC_16_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_19_LC_16_9_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_19_LC_16_9_0  (
            .in0(N__33255),
            .in1(N__52672),
            .in2(N__33237),
            .in3(N__52440),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_19_LC_16_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_19_LC_16_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_19_LC_16_9_1 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_19_LC_16_9_1  (
            .in0(N__33216),
            .in1(N__33210),
            .in2(N__51867),
            .in3(N__51510),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_19_LC_16_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_19_LC_16_9_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_19_LC_16_9_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_19_LC_16_9_2  (
            .in0(N__35217),
            .in1(N__33438),
            .in2(N__33204),
            .in3(N__33195),
            .lcout(I2C_top_level_inst1_s_data_oreg_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65513),
            .ce(N__54509),
            .sr(N__65003));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_19_LC_16_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_19_LC_16_9_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_19_LC_16_9_3 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_19_LC_16_9_3  (
            .in0(N__52145),
            .in1(N__33201),
            .in2(_gnd_net_),
            .in3(N__48681),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_19_LC_16_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_19_LC_16_9_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_19_LC_16_9_4 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_19_LC_16_9_4  (
            .in0(N__52982),
            .in1(N__57330),
            .in2(N__53324),
            .in3(N__51477),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_1_LC_16_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_1_LC_16_10_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_1_LC_16_10_0 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_1_LC_16_10_0  (
            .in0(N__56606),
            .in1(N__47415),
            .in2(N__47307),
            .in3(N__42888),
            .lcout(s_paddr_I2C_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65517),
            .ce(N__50091),
            .sr(N__64999));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_2_LC_16_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_2_LC_16_10_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_2_LC_16_10_1 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_2_LC_16_10_1  (
            .in0(N__47414),
            .in1(N__56607),
            .in2(N__47271),
            .in3(N__42870),
            .lcout(s_paddr_I2C_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65517),
            .ce(N__50091),
            .sr(N__64999));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_1_0_LC_16_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_1_0_LC_16_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_1_0_LC_16_10_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_1_0_LC_16_10_3  (
            .in0(N__35989),
            .in1(N__36268),
            .in2(N__43514),
            .in3(N__64172),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_0_LC_16_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_0_LC_16_10_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_0_LC_16_10_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_0_LC_16_10_4  (
            .in0(N__64174),
            .in1(N__43436),
            .in2(N__36273),
            .in3(N__35988),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIRQ9DD_0_LC_16_10_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIRQ9DD_0_LC_16_10_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIRQ9DD_0_LC_16_10_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIRQ9DD_0_LC_16_10_5  (
            .in0(N__43435),
            .in1(N__33431),
            .in2(_gnd_net_),
            .in3(N__64173),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1319_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_0_LC_16_10_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_0_LC_16_10_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_0_LC_16_10_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_0_LC_16_10_6  (
            .in0(N__33408),
            .in1(N__33393),
            .in2(N__33375),
            .in3(N__52441),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_0_LC_16_10_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_0_LC_16_10_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_0_LC_16_10_7 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_0_LC_16_10_7  (
            .in0(_gnd_net_),
            .in1(N__52054),
            .in2(N__33372),
            .in3(N__48921),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_21_LC_16_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_21_LC_16_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_21_LC_16_11_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_21_LC_16_11_0  (
            .in0(N__52903),
            .in1(N__37642),
            .in2(N__33369),
            .in3(N__46317),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_1_LC_16_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_1_LC_16_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_1_LC_16_11_1 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_1_LC_16_11_1  (
            .in0(N__37641),
            .in1(N__52901),
            .in2(N__34641),
            .in3(N__60710),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIH49MI_2_LC_16_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIH49MI_2_LC_16_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIH49MI_2_LC_16_11_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIH49MI_2_LC_16_11_2  (
            .in0(N__64235),
            .in1(N__35987),
            .in2(N__43581),
            .in3(N__36305),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_18_LC_16_11_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_18_LC_16_11_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_18_LC_16_11_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_18_LC_16_11_3  (
            .in0(N__33525),
            .in1(N__52902),
            .in2(N__33501),
            .in3(N__51368),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_20_LC_16_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_20_LC_16_11_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_20_LC_16_11_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_20_LC_16_11_4  (
            .in0(N__52904),
            .in1(N__37643),
            .in2(N__33486),
            .in3(N__40986),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_LC_16_11_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_LC_16_11_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_LC_16_11_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_LC_16_11_5  (
            .in0(N__35986),
            .in1(N__36362),
            .in2(N__43582),
            .in3(N__64236),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_7_LC_16_11_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_7_LC_16_11_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_7_LC_16_11_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_7_LC_16_11_6  (
            .in0(N__45534),
            .in1(N__33825),
            .in2(N__33459),
            .in3(N__37640),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15_LC_16_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15_LC_16_12_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15_LC_16_12_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15_LC_16_12_0  (
            .in0(N__60158),
            .in1(_gnd_net_),
            .in2(N__33600),
            .in3(N__33635),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net ),
            .ce(N__60004),
            .sr(N__62881));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI26492_17_LC_16_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI26492_17_LC_16_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI26492_17_LC_16_12_1 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI26492_17_LC_16_12_1  (
            .in0(N__53375),
            .in1(N__58190),
            .in2(N__48585),
            .in3(N__58005),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGH5_LC_16_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGH5_LC_16_12_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGH5_LC_16_12_2 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGH5_LC_16_12_2  (
            .in0(N__60565),
            .in1(N__42396),
            .in2(N__33441),
            .in3(N__46211),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI2UAV5_LC_16_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI2UAV5_LC_16_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI2UAV5_LC_16_12_3 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI2UAV5_LC_16_12_3  (
            .in0(N__33636),
            .in1(_gnd_net_),
            .in2(N__33639),
            .in3(N__60381),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITOAV5_LC_16_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITOAV5_LC_16_12_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITOAV5_LC_16_12_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITOAV5_LC_16_12_4  (
            .in0(N__33627),
            .in1(N__60380),
            .in2(_gnd_net_),
            .in3(N__33579),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_14_LC_16_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_14_LC_16_12_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_14_LC_16_12_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_14_LC_16_12_5  (
            .in0(_gnd_net_),
            .in1(N__33621),
            .in2(N__33603),
            .in3(N__60157),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net ),
            .ce(N__60004),
            .sr(N__62881));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI04492_17_LC_16_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI04492_17_LC_16_12_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI04492_17_LC_16_12_6 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI04492_17_LC_16_12_6  (
            .in0(N__58004),
            .in1(N__38479),
            .in2(N__58198),
            .in3(N__53420),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGH5_LC_16_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGH5_LC_16_12_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGH5_LC_16_12_7 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGH5_LC_16_12_7  (
            .in0(N__60558),
            .in1(N__33557),
            .in2(N__33591),
            .in3(N__33588),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGHZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2TV43_LC_16_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2TV43_LC_16_13_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2TV43_LC_16_13_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2TV43_LC_16_13_0  (
            .in0(N__45990),
            .in1(N__45832),
            .in2(N__38480),
            .in3(N__33556),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8D7_LC_16_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8D7_LC_16_13_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8D7_LC_16_13_1 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8D7_LC_16_13_1  (
            .in0(N__53419),
            .in1(N__53978),
            .in2(N__33573),
            .in3(N__33570),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8DZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_14_LC_16_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_14_LC_16_13_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_14_LC_16_13_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_14_LC_16_13_2  (
            .in0(_gnd_net_),
            .in1(N__58497),
            .in2(_gnd_net_),
            .in3(N__59382),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65536),
            .ce(N__58869),
            .sr(N__62873));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2V153_LC_16_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2V153_LC_16_13_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2V153_LC_16_13_3 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2V153_LC_16_13_3  (
            .in0(N__45991),
            .in1(N__48964),
            .in2(N__45868),
            .in3(N__49003),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDD7_LC_16_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDD7_LC_16_13_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDD7_LC_16_13_4 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDD7_LC_16_13_4  (
            .in0(N__53979),
            .in1(N__42777),
            .in2(N__33792),
            .in3(N__51251),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDDZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISQUF7_LC_16_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISQUF7_LC_16_13_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISQUF7_LC_16_13_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISQUF7_LC_16_13_5  (
            .in0(N__36141),
            .in1(_gnd_net_),
            .in2(N__33789),
            .in3(N__53691),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_23_LC_16_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_23_LC_16_13_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_23_LC_16_13_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_23_LC_16_13_6  (
            .in0(_gnd_net_),
            .in1(N__61247),
            .in2(_gnd_net_),
            .in3(N__59383),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65536),
            .ce(N__58869),
            .sr(N__62873));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4JK93_LC_16_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4JK93_LC_16_13_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4JK93_LC_16_13_7 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4JK93_LC_16_13_7  (
            .in0(N__45831),
            .in1(N__45989),
            .in2(N__42176),
            .in3(N__33775),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_1_LC_16_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_1_LC_16_14_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_1_LC_16_14_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_1_LC_16_14_0  (
            .in0(_gnd_net_),
            .in1(N__61867),
            .in2(_gnd_net_),
            .in3(N__59188),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_3_LC_16_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_3_LC_16_14_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_3_LC_16_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_3_LC_16_14_1  (
            .in0(N__59185),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63939),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_4_LC_16_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_4_LC_16_14_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_4_LC_16_14_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_4_LC_16_14_2  (
            .in0(_gnd_net_),
            .in1(N__63809),
            .in2(_gnd_net_),
            .in3(N__59190),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_6_LC_16_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_6_LC_16_14_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_6_LC_16_14_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_6_LC_16_14_3  (
            .in0(N__59186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63580),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_26_LC_16_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_26_LC_16_14_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_26_LC_16_14_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_26_LC_16_14_4  (
            .in0(_gnd_net_),
            .in1(N__60921),
            .in2(_gnd_net_),
            .in3(N__59189),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_0Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_20_LC_16_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_20_LC_16_14_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_20_LC_16_14_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_20_LC_16_14_5  (
            .in0(N__59183),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61525),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_12_LC_16_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_12_LC_16_14_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_12_LC_16_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_12_LC_16_14_6  (
            .in0(_gnd_net_),
            .in1(N__58589),
            .in2(_gnd_net_),
            .in3(N__59187),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_30_LC_16_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_30_LC_16_14_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_30_LC_16_14_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_30_LC_16_14_7  (
            .in0(N__59184),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62184),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65546),
            .ce(N__49033),
            .sr(N__62865));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_15_LC_16_15_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_15_LC_16_15_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_15_LC_16_15_0 .LUT_INIT=16'b1110001011000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_15_LC_16_15_0  (
            .in0(N__64312),
            .in1(N__55927),
            .in2(N__50625),
            .in3(N__64081),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1654_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_15_LC_16_15_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_15_LC_16_15_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_15_LC_16_15_1 .LUT_INIT=16'b1100000011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_15_LC_16_15_1  (
            .in0(_gnd_net_),
            .in1(N__50592),
            .in2(N__34011),
            .in3(N__49875),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65556),
            .ce(),
            .sr(N__64975));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNI6TP01_7_LC_16_15_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNI6TP01_7_LC_16_15_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNI6TP01_7_LC_16_15_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNI6TP01_7_LC_16_15_2  (
            .in0(N__63448),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59164),
            .lcout(N_12_0),
            .ltout(N_12_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_7_LC_16_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_7_LC_16_15_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_7_LC_16_15_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_7_LC_16_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34008),
            .in3(N__64073),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_o2_LC_16_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_o2_LC_16_15_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_o2_LC_16_15_4 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_o2_LC_16_15_4  (
            .in0(N__36294),
            .in1(N__36785),
            .in2(_gnd_net_),
            .in3(N__34852),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_RNO_0_7_LC_16_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_RNO_0_7_LC_16_15_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_RNO_0_7_LC_16_15_5 .LUT_INIT=16'b0101001111110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_RNO_0_7_LC_16_15_5  (
            .in0(N__36396),
            .in1(N__33821),
            .in2(N__33807),
            .in3(N__33804),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_5_LC_16_15_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_5_LC_16_15_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_5_LC_16_15_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_5_LC_16_15_6  (
            .in0(N__50558),
            .in1(N__56308),
            .in2(_gnd_net_),
            .in3(N__38657),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_a3_2_7_LC_16_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_a3_2_7_LC_16_15_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_a3_2_7_LC_16_15_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_a3_2_7_LC_16_15_7  (
            .in0(N__59165),
            .in1(N__34856),
            .in2(N__36789),
            .in3(N__36295),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_1786_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_26_LC_16_16_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_26_LC_16_16_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_26_LC_16_16_1 .LUT_INIT=16'b0000000000001011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_26_LC_16_16_1  (
            .in0(N__34083),
            .in1(N__34074),
            .in2(N__66813),
            .in3(N__64074),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_4093_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.N_536_i_i_o2_LC_16_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.N_536_i_i_o2_LC_16_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.N_536_i_i_o2_LC_16_16_2 .LUT_INIT=16'b0011000000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.N_536_i_i_o2_LC_16_16_2  (
            .in0(N__46807),
            .in1(N__64117),
            .in2(N__39660),
            .in3(N__39145),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISBI9D_0_LC_16_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISBI9D_0_LC_16_16_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISBI9D_0_LC_16_16_3 .LUT_INIT=16'b1000000010000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISBI9D_0_LC_16_16_3  (
            .in0(N__43366),
            .in1(N__37804),
            .in2(N__64209),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1320 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_LC_16_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_LC_16_16_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_LC_16_16_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_LC_16_16_4  (
            .in0(N__47111),
            .in1(N__34062),
            .in2(_gnd_net_),
            .in3(N__39144),
            .lcout(N_409),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_2_LC_16_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_2_LC_16_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_2_LC_16_16_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_2_LC_16_16_5  (
            .in0(N__47172),
            .in1(N__54334),
            .in2(N__56151),
            .in3(N__41609),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2),
            .ltout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIAC0UC_7_LC_16_16_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIAC0UC_7_LC_16_16_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIAC0UC_7_LC_16_16_6 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIAC0UC_7_LC_16_16_6  (
            .in0(N__47110),
            .in1(N__50244),
            .in2(N__34056),
            .in3(N__39143),
            .lcout(N_1838_0),
            .ltout(N_1838_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ91HD_0_LC_16_16_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ91HD_0_LC_16_16_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ91HD_0_LC_16_16_7 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ91HD_0_LC_16_16_7  (
            .in0(N__43365),
            .in1(_gnd_net_),
            .in2(N__34053),
            .in3(N__34049),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1314 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE6LS1_15_LC_16_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE6LS1_15_LC_16_17_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE6LS1_15_LC_16_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE6LS1_15_LC_16_17_0  (
            .in0(N__43235),
            .in1(N__43268),
            .in2(N__43205),
            .in3(N__43034),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_12_LC_16_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_12_LC_16_17_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_12_LC_16_17_3 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_12_LC_16_17_3  (
            .in0(N__64574),
            .in1(N__47411),
            .in2(N__41487),
            .in3(N__43023),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65582),
            .ce(N__50087),
            .sr(N__64976));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_13_LC_16_17_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_13_LC_16_17_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_13_LC_16_17_4 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_13_LC_16_17_4  (
            .in0(N__47409),
            .in1(N__64576),
            .in2(N__41469),
            .in3(N__43257),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65582),
            .ce(N__50087),
            .sr(N__64976));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_14_LC_16_17_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_14_LC_16_17_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_14_LC_16_17_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_14_LC_16_17_5  (
            .in0(N__64575),
            .in1(N__47412),
            .in2(N__41454),
            .in3(N__43224),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65582),
            .ce(N__50087),
            .sr(N__64976));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_15_LC_16_17_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_15_LC_16_17_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_15_LC_16_17_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_15_LC_16_17_6  (
            .in0(N__47410),
            .in1(N__64577),
            .in2(N__41439),
            .in3(N__43185),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65582),
            .ce(N__50087),
            .sr(N__64976));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_0_LC_16_18_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_0_LC_16_18_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_0_LC_16_18_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_0_LC_16_18_0  (
            .in0(N__57685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.s_data_ireg_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(N__36503),
            .sr(N__62843));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_1_LC_16_18_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_1_LC_16_18_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_1_LC_16_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_1_LC_16_18_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48262),
            .lcout(\I2C_top_level_inst1.s_data_ireg_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(N__36503),
            .sr(N__62843));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_7_LC_16_18_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_7_LC_16_18_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_7_LC_16_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_7_LC_16_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41733),
            .lcout(\I2C_top_level_inst1.s_data_ireg_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(N__36503),
            .sr(N__62843));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_5_LC_16_18_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_5_LC_16_18_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_5_LC_16_18_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_5_LC_16_18_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41375),
            .lcout(\I2C_top_level_inst1.s_data_ireg_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(N__36503),
            .sr(N__62843));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_2_LC_16_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_2_LC_16_18_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_2_LC_16_18_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_2_LC_16_18_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48140),
            .lcout(\I2C_top_level_inst1.s_data_ireg_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(N__36503),
            .sr(N__62843));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_4_LC_16_18_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_4_LC_16_18_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_4_LC_16_18_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_4_LC_16_18_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48032),
            .lcout(\I2C_top_level_inst1.s_data_ireg_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47983),
            .ce(N__36503),
            .sr(N__62843));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIEDSM_1_LC_16_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIEDSM_1_LC_16_19_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIEDSM_1_LC_16_19_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIEDSM_1_LC_16_19_0  (
            .in0(N__34167),
            .in1(N__34449),
            .in2(N__34149),
            .in3(N__34313),
            .lcout(\I2C_top_level_inst1.N_327_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_6_LC_16_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_6_LC_16_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_6_LC_16_19_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_6_LC_16_19_1  (
            .in0(N__50874),
            .in1(N__36634),
            .in2(_gnd_net_),
            .in3(N__34168),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1400_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_6_LC_16_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_6_LC_16_19_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_6_LC_16_19_2 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_6_LC_16_19_2  (
            .in0(N__36657),
            .in1(N__34404),
            .in2(N__34302),
            .in3(N__34381),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net ),
            .ce(),
            .sr(N__64984));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNILBK01_6_LC_16_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNILBK01_6_LC_16_19_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNILBK01_6_LC_16_19_3 .LUT_INIT=16'b0000101110101011;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNILBK01_6_LC_16_19_3  (
            .in0(N__50873),
            .in1(N__34166),
            .in2(N__34458),
            .in3(N__41574),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1374_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIAT631_3_LC_16_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIAT631_3_LC_16_19_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIAT631_3_LC_16_19_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIAT631_3_LC_16_19_4  (
            .in0(N__34281),
            .in1(N__34248),
            .in2(N__34224),
            .in3(N__34197),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0 ),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1354_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_7_LC_16_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_7_LC_16_19_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_7_LC_16_19_5 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_7_LC_16_19_5  (
            .in0(N__50872),
            .in1(_gnd_net_),
            .in2(N__34173),
            .in3(N__34169),
            .lcout(\I2C_top_level_inst1.s_load_addr1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net ),
            .ce(),
            .sr(N__64984));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_11_LC_16_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_11_LC_16_19_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_11_LC_16_19_6 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_11_LC_16_19_6  (
            .in0(N__41576),
            .in1(N__50871),
            .in2(N__36647),
            .in3(N__34454),
            .lcout(\I2C_top_level_inst1.s_load_wdata ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net ),
            .ce(),
            .sr(N__64984));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_1_LC_16_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_1_LC_16_19_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_1_LC_16_19_7 .LUT_INIT=16'b0101010011111100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_1_LC_16_19_7  (
            .in0(N__34453),
            .in1(N__34146),
            .in2(N__50885),
            .in3(N__41575),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_10_LC_16_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_10_LC_16_20_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_10_LC_16_20_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_10_LC_16_20_0  (
            .in0(N__34455),
            .in1(N__41521),
            .in2(N__43733),
            .in3(N__66275),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1399_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_10_LC_16_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_10_LC_16_20_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_10_LC_16_20_1 .LUT_INIT=16'b0000111100001011;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_10_LC_16_20_1  (
            .in0(N__43720),
            .in1(N__50884),
            .in2(N__34473),
            .in3(N__41577),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIIMIE_11_LC_16_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIIMIE_11_LC_16_20_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIIMIE_11_LC_16_20_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIIMIE_11_LC_16_20_2  (
            .in0(N__50883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50979),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1373_0 ),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1373_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_10_LC_16_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_10_LC_16_20_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_10_LC_16_20_3 .LUT_INIT=16'b0001000100000001;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_10_LC_16_20_3  (
            .in0(N__43721),
            .in1(N__34456),
            .in2(N__34470),
            .in3(N__34382),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1395_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_10_LC_16_20_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_10_LC_16_20_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_10_LC_16_20_4 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_10_LC_16_20_4  (
            .in0(N__34457),
            .in1(N__36643),
            .in2(N__34467),
            .in3(N__34464),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net ),
            .ce(),
            .sr(N__64989));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_9_LC_16_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_9_LC_16_20_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_9_LC_16_20_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_9_LC_16_20_5  (
            .in0(N__36642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34428),
            .lcout(\I2C_top_level_inst1.s_load_addr0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net ),
            .ce(),
            .sr(N__64989));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_14_LC_16_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_14_LC_16_20_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_14_LC_16_20_6 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_14_LC_16_20_6  (
            .in0(N__34403),
            .in1(N__41522),
            .in2(_gnd_net_),
            .in3(N__66276),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1409_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_14_LC_16_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_14_LC_16_20_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_14_LC_16_20_7 .LUT_INIT=16'b1111110111110101;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_14_LC_16_20_7  (
            .in0(N__34392),
            .in1(N__43938),
            .in2(N__34386),
            .in3(N__34383),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net ),
            .ce(),
            .sr(N__64989));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_2_LC_16_21_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_2_LC_16_21_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_2_LC_16_21_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_2_LC_16_21_0  (
            .in0(N__37149),
            .in1(N__37108),
            .in2(N__34557),
            .in3(N__36735),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_14_LC_16_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_14_LC_16_21_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_14_LC_16_21_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_14_LC_16_21_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34556),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65626),
            .ce(),
            .sr(N__62828));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_LC_16_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_LC_16_21_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_LC_16_21_2 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_LC_16_21_2  (
            .in0(N__34555),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36736),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1880 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65626),
            .ce(),
            .sr(N__62828));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_10_LC_16_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_10_LC_16_21_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_10_LC_16_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_10_LC_16_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37032),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65626),
            .ce(),
            .sr(N__62828));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI6HM8_10_LC_16_21_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI6HM8_10_LC_16_21_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI6HM8_10_LC_16_21_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI6HM8_10_LC_16_21_4  (
            .in0(_gnd_net_),
            .in1(N__36734),
            .in2(_gnd_net_),
            .in3(N__36714),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_1848_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_1848_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIVI6G_15_LC_16_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIVI6G_15_LC_16_21_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIVI6G_15_LC_16_21_5 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIVI6G_15_LC_16_21_5  (
            .in0(_gnd_net_),
            .in1(N__37148),
            .in2(N__34515),
            .in3(N__35724),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1884_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_15_LC_16_21_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_15_LC_16_21_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_15_LC_16_21_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_15_LC_16_21_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36737),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65626),
            .ce(),
            .sr(N__62828));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_11_LC_16_21_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_11_LC_16_21_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_11_LC_16_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_11_LC_16_21_7  (
            .in0(N__36715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65626),
            .ce(),
            .sr(N__62828));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI2MBM1_5_LC_16_22_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI2MBM1_5_LC_16_22_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI2MBM1_5_LC_16_22_0 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI2MBM1_5_LC_16_22_0  (
            .in0(N__34654),
            .in1(N__35394),
            .in2(N__34639),
            .in3(N__34597),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_0_LC_16_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_0_LC_16_22_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_0_LC_16_22_1 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_0_LC_16_22_1  (
            .in0(_gnd_net_),
            .in1(N__37031),
            .in2(N__34488),
            .in3(N__37064),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0_a2_6_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_LC_16_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_LC_16_22_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_LC_16_22_2 .LUT_INIT=16'b1101010111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_LC_16_22_2  (
            .in0(N__35795),
            .in1(N__34485),
            .in2(N__34476),
            .in3(N__34701),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65642),
            .ce(),
            .sr(N__62822));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_1_LC_16_22_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_1_LC_16_22_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_1_LC_16_22_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_1_LC_16_22_3  (
            .in0(N__35360),
            .in1(N__35915),
            .in2(N__34710),
            .in3(N__37019),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNIDMPS1_LC_16_22_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNIDMPS1_LC_16_22_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNIDMPS1_LC_16_22_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNIDMPS1_LC_16_22_4  (
            .in0(N__34695),
            .in1(N__34680),
            .in2(_gnd_net_),
            .in3(N__34689),
            .lcout(c_state_ret_12_RNIDMPS1_0),
            .ltout(c_state_ret_12_RNIDMPS1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.current_state_0_LC_16_22_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_0_LC_16_22_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.current_state_0_LC_16_22_5 .LUT_INIT=16'b0011001000010000;
    LogicCell40 \serializer_mod_inst.current_state_0_LC_16_22_5  (
            .in0(N__45469),
            .in1(N__44899),
            .in2(N__34674),
            .in3(N__45498),
            .lcout(\serializer_mod_inst.current_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65642),
            .ce(),
            .sr(N__62822));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_LC_16_22_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_LC_16_22_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_LC_16_22_6 .LUT_INIT=16'b0000000001010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_LC_16_22_6  (
            .in0(N__34655),
            .in1(N__35395),
            .in2(N__34640),
            .in3(N__34598),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65642),
            .ce(),
            .sr(N__62822));
    defparam \serializer_mod_inst.shift_reg_7_LC_16_23_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_7_LC_16_23_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_7_LC_16_23_1 .LUT_INIT=16'b0101101000001010;
    LogicCell40 \serializer_mod_inst.shift_reg_7_LC_16_23_1  (
            .in0(N__44894),
            .in1(_gnd_net_),
            .in2(N__45464),
            .in3(N__41847),
            .lcout(\serializer_mod_inst.shift_regZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65653),
            .ce(),
            .sr(N__62817));
    defparam \serializer_mod_inst.shift_reg_11_LC_16_23_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_11_LC_16_23_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_11_LC_16_23_2 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_11_LC_16_23_2  (
            .in0(N__37239),
            .in1(N__45422),
            .in2(_gnd_net_),
            .in3(N__44895),
            .lcout(\serializer_mod_inst.shift_regZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65653),
            .ce(),
            .sr(N__62817));
    defparam \serializer_mod_inst.shift_reg_8_LC_16_23_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_8_LC_16_23_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_8_LC_16_23_4 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_8_LC_16_23_4  (
            .in0(N__34575),
            .in1(N__45426),
            .in2(_gnd_net_),
            .in3(N__44896),
            .lcout(\serializer_mod_inst.shift_regZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65653),
            .ce(),
            .sr(N__62817));
    defparam \serializer_mod_inst.shift_reg_31_LC_16_24_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_31_LC_16_24_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_31_LC_16_24_0 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_31_LC_16_24_0  (
            .in0(N__44214),
            .in1(N__45411),
            .in2(_gnd_net_),
            .in3(N__45033),
            .lcout(\serializer_mod_inst.shift_regZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65668),
            .ce(),
            .sr(N__62812));
    defparam \serializer_mod_inst.shift_reg_32_LC_16_24_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_32_LC_16_24_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_32_LC_16_24_1 .LUT_INIT=16'b0011110000001100;
    LogicCell40 \serializer_mod_inst.shift_reg_32_LC_16_24_1  (
            .in0(_gnd_net_),
            .in1(N__44949),
            .in2(N__45462),
            .in3(N__34569),
            .lcout(\serializer_mod_inst.shift_regZ0Z_32 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65668),
            .ce(),
            .sr(N__62812));
    defparam \serializer_mod_inst.shift_reg_48_LC_16_24_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_48_LC_16_24_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_48_LC_16_24_2 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_48_LC_16_24_2  (
            .in0(N__37347),
            .in1(N__45415),
            .in2(_gnd_net_),
            .in3(N__45034),
            .lcout(\serializer_mod_inst.shift_regZ0Z_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65668),
            .ce(),
            .sr(N__62812));
    defparam \serializer_mod_inst.shift_reg_115_LC_16_24_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_115_LC_16_24_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_115_LC_16_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_115_LC_16_24_3  (
            .in0(_gnd_net_),
            .in1(N__34746),
            .in2(_gnd_net_),
            .in3(N__47876),
            .lcout(\serializer_mod_inst.shift_regZ0Z_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65668),
            .ce(),
            .sr(N__62812));
    defparam \serializer_mod_inst.shift_reg_114_LC_16_24_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_114_LC_16_24_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_114_LC_16_24_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_114_LC_16_24_5  (
            .in0(_gnd_net_),
            .in1(N__34755),
            .in2(_gnd_net_),
            .in3(N__47875),
            .lcout(\serializer_mod_inst.shift_regZ0Z_114 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65668),
            .ce(),
            .sr(N__62812));
    defparam \serializer_mod_inst.shift_reg_79_LC_16_25_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_79_LC_16_25_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_79_LC_16_25_0 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_79_LC_16_25_0  (
            .in0(N__45027),
            .in1(N__34722),
            .in2(_gnd_net_),
            .in3(N__45406),
            .lcout(\serializer_mod_inst.shift_regZ0Z_79 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65680),
            .ce(),
            .sr(N__62809));
    defparam \serializer_mod_inst.shift_reg_110_LC_16_25_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_110_LC_16_25_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_110_LC_16_25_1 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_110_LC_16_25_1  (
            .in0(N__45403),
            .in1(N__41922),
            .in2(_gnd_net_),
            .in3(N__45028),
            .lcout(\serializer_mod_inst.shift_regZ0Z_110 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65680),
            .ce(),
            .sr(N__62809));
    defparam \serializer_mod_inst.shift_reg_40_LC_16_25_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_40_LC_16_25_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_40_LC_16_25_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_40_LC_16_25_2  (
            .in0(N__45026),
            .in1(N__34734),
            .in2(_gnd_net_),
            .in3(N__45404),
            .lcout(\serializer_mod_inst.shift_regZ0Z_40 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65680),
            .ce(),
            .sr(N__62809));
    defparam \serializer_mod_inst.shift_reg_78_LC_16_25_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_78_LC_16_25_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_78_LC_16_25_3 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_78_LC_16_25_3  (
            .in0(N__45405),
            .in1(N__34728),
            .in2(_gnd_net_),
            .in3(N__45029),
            .lcout(\serializer_mod_inst.shift_regZ0Z_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65680),
            .ce(),
            .sr(N__62809));
    defparam \serializer_mod_inst.shift_reg_41_LC_16_25_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_41_LC_16_25_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_41_LC_16_25_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_41_LC_16_25_7  (
            .in0(_gnd_net_),
            .in1(N__34716),
            .in2(_gnd_net_),
            .in3(N__47874),
            .lcout(\serializer_mod_inst.shift_regZ0Z_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65680),
            .ce(),
            .sr(N__62809));
    defparam \serializer_mod_inst.shift_reg_67_LC_16_26_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_67_LC_16_26_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_67_LC_16_26_0 .LUT_INIT=16'b0011110000001100;
    LogicCell40 \serializer_mod_inst.shift_reg_67_LC_16_26_0  (
            .in0(_gnd_net_),
            .in1(N__45058),
            .in2(N__45357),
            .in3(N__40176),
            .lcout(\serializer_mod_inst.shift_regZ0Z_67 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65692),
            .ce(),
            .sr(N__62806));
    defparam \serializer_mod_inst.shift_reg_69_LC_16_26_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_69_LC_16_26_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_69_LC_16_26_2 .LUT_INIT=16'b0011110000001100;
    LogicCell40 \serializer_mod_inst.shift_reg_69_LC_16_26_2  (
            .in0(_gnd_net_),
            .in1(N__45059),
            .in2(N__45358),
            .in3(N__34884),
            .lcout(\serializer_mod_inst.shift_regZ0Z_69 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65692),
            .ce(),
            .sr(N__62806));
    defparam \serializer_mod_inst.shift_reg_68_LC_16_26_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_68_LC_16_26_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_68_LC_16_26_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_68_LC_16_26_4  (
            .in0(N__47812),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34890),
            .lcout(\serializer_mod_inst.shift_regZ0Z_68 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65692),
            .ce(),
            .sr(N__62806));
    defparam \serializer_mod_inst.shift_reg_116_LC_16_26_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_116_LC_16_26_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_116_LC_16_26_5 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \serializer_mod_inst.shift_reg_116_LC_16_26_5  (
            .in0(N__34878),
            .in1(N__47811),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\serializer_mod_inst.shift_regZ0Z_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65692),
            .ce(),
            .sr(N__62806));
    defparam \serializer_mod_inst.shift_reg_117_LC_16_26_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_117_LC_16_26_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_117_LC_16_26_7 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_117_LC_16_26_7  (
            .in0(N__34869),
            .in1(N__45232),
            .in2(_gnd_net_),
            .in3(N__45060),
            .lcout(\serializer_mod_inst.shift_regZ0Z_117 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65692),
            .ce(),
            .sr(N__62806));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_0_a2_0_LC_16_27_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_0_a2_0_LC_16_27_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_0_a2_0_LC_16_27_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_0_a2_0_LC_16_27_6  (
            .in0(N__38679),
            .in1(N__36366),
            .in2(_gnd_net_),
            .in3(N__34857),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_n_ibuf_RNIBNDC_LC_16_32_2.C_ON=1'b0;
    defparam rst_n_ibuf_RNIBNDC_LC_16_32_2.SEQ_MODE=4'b0000;
    defparam rst_n_ibuf_RNIBNDC_LC_16_32_2.LUT_INIT=16'b0000000011111111;
    LogicCell40 rst_n_ibuf_RNIBNDC_LC_16_32_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35464),
            .lcout(rst_n_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_12_LC_17_8_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_12_LC_17_8_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_12_LC_17_8_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_12_LC_17_8_6  (
            .in0(N__52146),
            .in1(N__41234),
            .in2(N__53317),
            .in3(N__40961),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_12_LC_17_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_12_LC_17_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_12_LC_17_9_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_12_LC_17_9_0  (
            .in0(N__34800),
            .in1(N__52675),
            .in2(N__34779),
            .in3(N__52484),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_12_LC_17_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_12_LC_17_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_12_LC_17_9_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_12_LC_17_9_1  (
            .in0(_gnd_net_),
            .in1(N__53000),
            .in2(N__34758),
            .in3(N__46350),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_12_LC_17_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_12_LC_17_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_12_LC_17_9_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_12_LC_17_9_2  (
            .in0(N__35154),
            .in1(N__44661),
            .in2(N__63831),
            .in3(N__44427),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_12_LC_17_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_12_LC_17_9_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_12_LC_17_9_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_12_LC_17_9_3  (
            .in0(N__35136),
            .in1(N__51824),
            .in2(N__35124),
            .in3(N__41202),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_12_LC_17_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_12_LC_17_9_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_12_LC_17_9_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_12_LC_17_9_4  (
            .in0(N__35037),
            .in1(N__35121),
            .in2(N__35115),
            .in3(N__35112),
            .lcout(I2C_top_level_inst1_s_data_oreg_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65520),
            .ce(N__54505),
            .sr(N__65005));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_11_LC_17_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_11_LC_17_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_11_LC_17_10_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_11_LC_17_10_1  (
            .in0(N__38220),
            .in1(N__37649),
            .in2(N__35106),
            .in3(N__42951),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_12_LC_17_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_12_LC_17_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_12_LC_17_10_2 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_12_LC_17_10_2  (
            .in0(N__37650),
            .in1(N__38221),
            .in2(N__35070),
            .in3(N__42705),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_13_LC_17_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_13_LC_17_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_13_LC_17_10_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_13_LC_17_10_3  (
            .in0(N__38216),
            .in1(N__37645),
            .in2(N__35031),
            .in3(N__42813),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_14_LC_17_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_14_LC_17_10_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_14_LC_17_10_4 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_14_LC_17_10_4  (
            .in0(N__37644),
            .in1(N__38215),
            .in2(N__34992),
            .in3(N__42643),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_15_LC_17_10_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_15_LC_17_10_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_15_LC_17_10_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_15_LC_17_10_5  (
            .in0(N__38218),
            .in1(N__37648),
            .in2(N__34953),
            .in3(N__42612),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_16_LC_17_10_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_16_LC_17_10_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_16_LC_17_10_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_16_LC_17_10_6  (
            .in0(N__37647),
            .in1(N__38219),
            .in2(N__34914),
            .in3(N__42582),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_17_LC_17_10_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_17_LC_17_10_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_17_LC_17_10_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_17_LC_17_10_7  (
            .in0(N__38217),
            .in1(N__37646),
            .in2(N__35340),
            .in3(N__45617),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_3_0_LC_17_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_3_0_LC_17_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_3_0_LC_17_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_3_0_LC_17_11_0  (
            .in0(N__36355),
            .in1(N__35996),
            .in2(N__43583),
            .in3(N__64234),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_2_LC_17_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_2_LC_17_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_2_LC_17_11_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_2_LC_17_11_1  (
            .in0(N__37656),
            .in1(N__35304),
            .in2(N__35283),
            .in3(N__42975),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_24_LC_17_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_24_LC_17_11_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_24_LC_17_11_4 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_24_LC_17_11_4  (
            .in0(N__38238),
            .in1(N__35268),
            .in2(N__35250),
            .in3(N__37657),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_24_LC_17_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_24_LC_17_11_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_24_LC_17_11_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_24_LC_17_11_5  (
            .in0(N__61103),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59388),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65531),
            .ce(N__45570),
            .sr(N__62907));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_19_LC_17_11_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_19_LC_17_11_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_19_LC_17_11_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_19_LC_17_11_6  (
            .in0(N__38237),
            .in1(N__37655),
            .in2(N__35241),
            .in3(N__48705),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_25_LC_17_11_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_25_LC_17_11_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_25_LC_17_11_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_25_LC_17_11_7  (
            .in0(N__37658),
            .in1(N__38239),
            .in2(N__44238),
            .in3(N__35205),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_27_LC_17_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_27_LC_17_12_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_27_LC_17_12_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_27_LC_17_12_0  (
            .in0(N__35184),
            .in1(N__38214),
            .in2(N__35163),
            .in3(N__37654),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_27_LC_17_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_27_LC_17_12_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_27_LC_17_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_27_LC_17_12_1  (
            .in0(_gnd_net_),
            .in1(N__60797),
            .in2(_gnd_net_),
            .in3(N__59384),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65541),
            .ce(N__45568),
            .sr(N__62896));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_28_LC_17_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_28_LC_17_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_28_LC_17_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_28_LC_17_12_2  (
            .in0(N__35655),
            .in1(N__38213),
            .in2(N__35619),
            .in3(N__37653),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_28_LC_17_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_28_LC_17_12_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_28_LC_17_12_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_28_LC_17_12_3  (
            .in0(_gnd_net_),
            .in1(N__62336),
            .in2(_gnd_net_),
            .in3(N__59385),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65541),
            .ce(N__45568),
            .sr(N__62896));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_29_LC_17_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_29_LC_17_12_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_29_LC_17_12_4 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_29_LC_17_12_4  (
            .in0(N__35610),
            .in1(N__38211),
            .in2(N__35589),
            .in3(N__37652),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_29_LC_17_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_29_LC_17_12_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_29_LC_17_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_29_LC_17_12_5  (
            .in0(N__62264),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59386),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65541),
            .ce(N__45568),
            .sr(N__62896));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_3_LC_17_12_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_3_LC_17_12_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_3_LC_17_12_6 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_3_LC_17_12_6  (
            .in0(N__35580),
            .in1(N__37651),
            .in2(N__35533),
            .in3(N__38212),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_3_LC_17_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_3_LC_17_12_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_3_LC_17_12_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_3_LC_17_12_7  (
            .in0(_gnd_net_),
            .in1(N__63923),
            .in2(_gnd_net_),
            .in3(N__59387),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65541),
            .ce(N__45568),
            .sr(N__62896));
    defparam \serializer_mod_inst.serial_out_test_e_0_LC_17_13_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.serial_out_test_e_0_LC_17_13_0 .SEQ_MODE=4'b1000;
    defparam \serializer_mod_inst.serial_out_test_e_0_LC_17_13_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \serializer_mod_inst.serial_out_test_e_0_LC_17_13_0  (
            .in0(N__44007),
            .in1(N__45485),
            .in2(_gnd_net_),
            .in3(N__45090),
            .lcout(serial_out_testing_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65551),
            .ce(N__35481),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIIO3I_0_LC_17_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIIO3I_0_LC_17_13_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIIO3I_0_LC_17_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIIO3I_0_LC_17_13_1  (
            .in0(_gnd_net_),
            .in1(N__40096),
            .in2(_gnd_net_),
            .in3(N__39791),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1965 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_6_LC_17_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_6_LC_17_13_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_6_LC_17_13_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_6_LC_17_13_2  (
            .in0(N__40097),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40002),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_522_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIMEFF_LC_17_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIMEFF_LC_17_13_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIMEFF_LC_17_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIMEFF_LC_17_13_3  (
            .in0(_gnd_net_),
            .in1(N__40041),
            .in2(_gnd_net_),
            .in3(N__40098),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO4JK_4_LC_17_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO4JK_4_LC_17_13_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO4JK_4_LC_17_13_4 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO4JK_4_LC_17_13_4  (
            .in0(N__35892),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35862),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIP1G7_15_LC_17_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIP1G7_15_LC_17_13_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIP1G7_15_LC_17_13_5 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIP1G7_15_LC_17_13_5  (
            .in0(_gnd_net_),
            .in1(N__37169),
            .in2(_gnd_net_),
            .in3(N__35761),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_1854_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIGUF7_LC_17_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIGUF7_LC_17_13_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIGUF7_LC_17_13_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIGUF7_LC_17_13_6  (
            .in0(N__36183),
            .in1(N__53692),
            .in2(_gnd_net_),
            .in3(N__45708),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINLUF7_LC_17_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINLUF7_LC_17_13_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINLUF7_LC_17_13_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINLUF7_LC_17_13_7  (
            .in0(N__53693),
            .in1(N__38403),
            .in2(_gnd_net_),
            .in3(N__36159),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIKSI1_LC_17_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIKSI1_LC_17_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIKSI1_LC_17_14_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIKSI1_LC_17_14_0  (
            .in0(N__55155),
            .in1(N__42412),
            .in2(N__55451),
            .in3(N__35680),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5Q7H2_LC_17_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5Q7H2_LC_17_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5Q7H2_LC_17_14_1 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5Q7H2_LC_17_14_1  (
            .in0(N__35681),
            .in1(N__55010),
            .in2(N__42419),
            .in3(N__54802),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DD7_LC_17_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DD7_LC_17_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DD7_LC_17_14_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DD7_LC_17_14_2  (
            .in0(N__53977),
            .in1(N__38566),
            .in2(N__35667),
            .in3(N__40800),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DDZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIDBUF7_LC_17_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIDBUF7_LC_17_14_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIDBUF7_LC_17_14_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIDBUF7_LC_17_14_3  (
            .in0(N__53671),
            .in1(_gnd_net_),
            .in2(N__35664),
            .in3(N__35661),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20_LC_17_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20_LC_17_14_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20_LC_17_14_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20_LC_17_14_4  (
            .in0(_gnd_net_),
            .in1(N__49191),
            .in2(N__36192),
            .in3(N__55686),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net ),
            .ce(N__55563),
            .sr(N__62878));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_21_LC_17_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_21_LC_17_14_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_21_LC_17_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_21_LC_17_14_5  (
            .in0(N__55687),
            .in1(N__36189),
            .in2(_gnd_net_),
            .in3(N__36182),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net ),
            .ce(N__55563),
            .sr(N__62878));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_22_LC_17_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_22_LC_17_14_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_22_LC_17_14_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_22_LC_17_14_6  (
            .in0(N__36171),
            .in1(N__55688),
            .in2(_gnd_net_),
            .in3(N__36158),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net ),
            .ce(N__55563),
            .sr(N__62878));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_23_LC_17_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_23_LC_17_14_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_23_LC_17_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_23_LC_17_14_7  (
            .in0(N__55689),
            .in1(N__36147),
            .in2(_gnd_net_),
            .in3(N__36140),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_conf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net ),
            .ce(N__55563),
            .sr(N__62878));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_2_0_LC_17_15_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_2_0_LC_17_15_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_2_0_LC_17_15_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_2_0_LC_17_15_0  (
            .in0(N__35990),
            .in1(N__36317),
            .in2(N__43569),
            .in3(N__64066),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_1_LC_17_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_1_LC_17_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_1_LC_17_15_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_1_LC_17_15_1  (
            .in0(N__64067),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35991),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1831_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_2 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_2  (
            .in0(N__36259),
            .in1(N__38656),
            .in2(N__35997),
            .in3(N__64068),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPOSB_11_LC_17_15_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPOSB_11_LC_17_15_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPOSB_11_LC_17_15_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPOSB_11_LC_17_15_3  (
            .in0(_gnd_net_),
            .in1(N__56868),
            .in2(_gnd_net_),
            .in3(N__57718),
            .lcout(N_1841_0),
            .ltout(N_1841_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_4 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_4  (
            .in0(N__35992),
            .in1(N__36354),
            .in2(N__35925),
            .in3(N__64069),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_12_LC_17_15_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_12_LC_17_15_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_12_LC_17_15_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_12_LC_17_15_5  (
            .in0(_gnd_net_),
            .in1(N__66184),
            .in2(_gnd_net_),
            .in3(N__57719),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65576),
            .ce(),
            .sr(N__64981));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_11_LC_17_15_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_11_LC_17_15_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_11_LC_17_15_6 .LUT_INIT=16'b0111000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_11_LC_17_15_6  (
            .in0(N__50943),
            .in1(N__50559),
            .in2(N__50490),
            .in3(N__47517),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65576),
            .ce(),
            .sr(N__64981));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_13_LC_17_15_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_13_LC_17_15_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_13_LC_17_15_7 .LUT_INIT=16'b0000000011101100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_13_LC_17_15_7  (
            .in0(N__43173),
            .in1(N__56869),
            .in2(N__56245),
            .in3(N__66185),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65576),
            .ce(),
            .sr(N__64981));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNINHAS1_0_LC_17_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNINHAS1_0_LC_17_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNINHAS1_0_LC_17_16_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNINHAS1_0_LC_17_16_0  (
            .in0(N__39036),
            .in1(N__46764),
            .in2(_gnd_net_),
            .in3(N__39113),
            .lcout(N_1613),
            .ltout(N_1613_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_1 .LUT_INIT=16'b0000101000001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_1  (
            .in0(N__39612),
            .in1(N__46900),
            .in2(N__36369),
            .in3(N__39132),
            .lcout(N_1860_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_2 .LUT_INIT=16'b0010001000001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_2  (
            .in0(N__36219),
            .in1(N__39611),
            .in2(N__46910),
            .in3(N__39116),
            .lcout(N_202_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII7LO3_2_LC_17_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII7LO3_2_LC_17_16_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII7LO3_2_LC_17_16_3 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII7LO3_2_LC_17_16_3  (
            .in0(N__39114),
            .in1(N__46896),
            .in2(N__39617),
            .in3(N__36218),
            .lcout(N_1859_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_4 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_4  (
            .in0(N__36220),
            .in1(N__39613),
            .in2(N__46909),
            .in3(N__39115),
            .lcout(N_1861_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_0_LC_17_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_0_LC_17_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_0_LC_17_16_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_0_LC_17_16_5  (
            .in0(N__48519),
            .in1(N__45588),
            .in2(_gnd_net_),
            .in3(N__36221),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_604 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI7T453_9_LC_17_16_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI7T453_9_LC_17_16_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI7T453_9_LC_17_16_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI7T453_9_LC_17_16_6  (
            .in0(N__47043),
            .in1(N__47013),
            .in2(N__46950),
            .in3(N__47456),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE7FP3_4_LC_17_16_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE7FP3_4_LC_17_16_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE7FP3_4_LC_17_16_7 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE7FP3_4_LC_17_16_7  (
            .in0(_gnd_net_),
            .in1(N__47243),
            .in2(N__36417),
            .in3(N__47206),
            .lcout(N_396),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_6_0_a3_0_o2_LC_17_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_6_0_a3_0_o2_LC_17_17_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_6_0_a3_0_o2_LC_17_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_6_0_a3_0_o2_LC_17_17_0  (
            .in0(N__36402),
            .in1(N__36408),
            .in2(N__36384),
            .in3(N__36414),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_4_LC_17_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_4_LC_17_17_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_4_LC_17_17_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_4_LC_17_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41377),
            .lcout(\I2C_top_level_inst1.s_command_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__47921),
            .sr(N__62858));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_5_LC_17_17_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_5_LC_17_17_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_5_LC_17_17_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_5_LC_17_17_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41796),
            .lcout(\I2C_top_level_inst1.s_command_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__47921),
            .sr(N__62858));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_6_LC_17_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_6_LC_17_17_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_6_LC_17_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_6_LC_17_17_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41734),
            .lcout(\I2C_top_level_inst1.s_command_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__47921),
            .sr(N__62858));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIFO5I1_7_LC_17_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIFO5I1_7_LC_17_17_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIFO5I1_7_LC_17_17_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIFO5I1_7_LC_17_17_4  (
            .in0(_gnd_net_),
            .in1(N__39455),
            .in2(_gnd_net_),
            .in3(N__39109),
            .lcout(N_1803),
            .ltout(N_1803_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_26_LC_17_17_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_26_LC_17_17_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_26_LC_17_17_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_26_LC_17_17_5  (
            .in0(N__37182),
            .in1(N__36519),
            .in2(N__36387),
            .in3(N__36375),
            .lcout(N_410),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_7_LC_17_17_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_7_LC_17_17_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_7_LC_17_17_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_7_LC_17_17_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41688),
            .lcout(\I2C_top_level_inst1.s_command_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47978),
            .ce(N__47921),
            .sr(N__62858));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6_26_LC_17_17_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6_26_LC_17_17_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6_26_LC_17_17_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6_26_LC_17_17_7  (
            .in0(N__39512),
            .in1(N__39536),
            .in2(N__39486),
            .in3(N__39566),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_a2_6_0_LC_17_18_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_a2_6_0_LC_17_18_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_a2_6_0_LC_17_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_a2_6_0_LC_17_18_0  (
            .in0(N__41729),
            .in1(N__41786),
            .in2(N__41658),
            .in3(N__41348),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_300_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_6_LC_17_18_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_6_LC_17_18_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_6_LC_17_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_6_LC_17_18_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41787),
            .lcout(\I2C_top_level_inst1.s_data_ireg_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47980),
            .ce(N__36510),
            .sr(N__62852));
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_3_LC_17_18_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_3_LC_17_18_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_3_LC_17_18_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_3_LC_17_18_5  (
            .in0(N__48081),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.s_data_ireg_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47980),
            .ce(N__36510),
            .sr(N__62852));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_a2_1_0_LC_17_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_a2_1_0_LC_17_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_a2_1_0_LC_17_18_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_a2_1_0_LC_17_18_6  (
            .in0(N__48020),
            .in1(N__48132),
            .in2(_gnd_net_),
            .in3(N__48080),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1425_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0_LC_17_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0_LC_17_19_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0_LC_17_19_0 .LUT_INIT=16'b1000100001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0_LC_17_19_0  (
            .in0(N__36486),
            .in1(N__36449),
            .in2(_gnd_net_),
            .in3(N__36472),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .ce(),
            .sr(N__64990));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIUAQ1_11_LC_17_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIUAQ1_11_LC_17_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIUAQ1_11_LC_17_19_1 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIUAQ1_11_LC_17_19_1  (
            .in0(_gnd_net_),
            .in1(N__50983),
            .in2(_gnd_net_),
            .in3(N__43954),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1367_0 ),
            .ltout(\I2C_top_level_inst1.I2C_FSM_inst.N_1367_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_1_LC_17_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_1_LC_17_19_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_1_LC_17_19_2 .LUT_INIT=16'b1100011000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_1_LC_17_19_2  (
            .in0(N__36473),
            .in1(N__36431),
            .in2(N__36453),
            .in3(N__36450),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .ce(),
            .sr(N__64990));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_r_w_LC_17_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_r_w_LC_17_19_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_r_w_LC_17_19_3 .LUT_INIT=16'b0101010000000100;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_r_w_LC_17_19_3  (
            .in0(N__43664),
            .in1(N__51299),
            .in2(N__43901),
            .in3(N__48258),
            .lcout(\I2C_top_level_inst1.s_r_w ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .ce(),
            .sr(N__64990));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_0_LC_17_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_0_LC_17_19_4 .SEQ_MODE=4'b1011;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_0_LC_17_19_4 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_0_LC_17_19_4  (
            .in0(N__43790),
            .in1(N__43665),
            .in2(N__43638),
            .in3(N__43852),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .ce(),
            .sr(N__64990));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_3_LC_17_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_3_LC_17_19_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_3_LC_17_19_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_3_LC_17_19_5  (
            .in0(N__43853),
            .in1(N__43828),
            .in2(_gnd_net_),
            .in3(N__43789),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .ce(),
            .sr(N__64990));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_6_LC_17_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_6_LC_17_19_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_6_LC_17_19_6 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_6_LC_17_19_6  (
            .in0(N__36678),
            .in1(N__47914),
            .in2(_gnd_net_),
            .in3(N__43887),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_5_LC_17_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_5_LC_17_19_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_5_LC_17_19_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_5_LC_17_19_7  (
            .in0(_gnd_net_),
            .in1(N__36641),
            .in2(_gnd_net_),
            .in3(N__36600),
            .lcout(\I2C_top_level_inst1.s_load_command ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net ),
            .ce(),
            .sr(N__64990));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_1_LC_17_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_1_LC_17_20_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_1_LC_17_20_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_1_LC_17_20_0  (
            .in0(N__36579),
            .in1(N__36561),
            .in2(N__43748),
            .in3(N__43956),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_1_LC_17_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_1_LC_17_20_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_1_LC_17_20_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_1_LC_17_20_1  (
            .in0(N__47912),
            .in1(N__41406),
            .in2(_gnd_net_),
            .in3(N__43885),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI8SIH_3_LC_17_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI8SIH_3_LC_17_20_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI8SIH_3_LC_17_20_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI8SIH_3_LC_17_20_2  (
            .in0(N__43886),
            .in1(N__47913),
            .in2(N__43749),
            .in3(N__41413),
            .lcout(),
            .ltout(\I2C_top_level_inst1.N_4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.s_sda_o_tx_RNITO2M_LC_17_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.s_sda_o_tx_RNITO2M_LC_17_20_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.s_sda_o_tx_RNITO2M_LC_17_20_3 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \I2C_top_level_inst1.s_sda_o_tx_RNITO2M_LC_17_20_3  (
            .in0(N__63292),
            .in1(N__36981),
            .in2(N__36555),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.N_259 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_552_i_0_a2_LC_17_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_552_i_0_a2_LC_17_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_552_i_0_a2_LC_17_20_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_552_i_0_a2_LC_17_20_4  (
            .in0(N__36530),
            .in1(N__62456),
            .in2(_gnd_net_),
            .in3(N__56878),
            .lcout(N_552_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7_26_LC_17_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7_26_LC_17_20_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7_26_LC_17_20_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7_26_LC_17_20_5  (
            .in0(N__39878),
            .in1(N__39893),
            .in2(N__39711),
            .in3(N__39908),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.s_sda_o_q_1_LC_17_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.s_sda_o_q_1_LC_17_20_6 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.s_sda_o_q_1_LC_17_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.s_sda_o_q_1_LC_17_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36975),
            .lcout(\I2C_top_level_inst1.s_sda_o_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65632),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.s_sda_o_tx_LC_17_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.s_sda_o_tx_LC_17_20_7 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.s_sda_o_tx_LC_17_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.s_sda_o_tx_LC_17_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36987),
            .lcout(\I2C_top_level_inst1.s_sda_o_txZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65632),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.s_sda_o_q_0_LC_17_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.s_sda_o_q_0_LC_17_21_0 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.s_sda_o_q_0_LC_17_21_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.s_sda_o_q_0_LC_17_21_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61989),
            .lcout(\I2C_top_level_inst1.s_sda_o_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65648),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_RNI8HA01_1_LC_17_21_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_RNI8HA01_1_LC_17_21_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_RNI8HA01_1_LC_17_21_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_RNI8HA01_1_LC_17_21_1  (
            .in0(_gnd_net_),
            .in1(N__36969),
            .in2(_gnd_net_),
            .in3(N__36908),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_1855_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_1855_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_RNI6LR22_LC_17_21_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_RNI6LR22_LC_17_21_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_RNI6LR22_LC_17_21_2 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_RNI6LR22_LC_17_21_2  (
            .in0(_gnd_net_),
            .in1(N__37005),
            .in2(N__36846),
            .in3(N__36838),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_1857_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.N_1857_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_a2_LC_17_21_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_a2_LC_17_21_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_a2_LC_17_21_3 .LUT_INIT=16'b0100111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_a2_LC_17_21_3  (
            .in0(N__36770),
            .in1(N__36689),
            .in2(N__36792),
            .in3(N__39146),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_384 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_2_o2_0_LC_17_21_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_2_o2_0_LC_17_21_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_2_o2_0_LC_17_21_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_2_o2_0_LC_17_21_4  (
            .in0(N__36771),
            .in1(N__37048),
            .in2(_gnd_net_),
            .in3(N__37107),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1840_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI1ITL_8_LC_17_21_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI1ITL_8_LC_17_21_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI1ITL_8_LC_17_21_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI1ITL_8_LC_17_21_5  (
            .in0(N__37106),
            .in1(N__36738),
            .in2(N__37050),
            .in3(N__36716),
            .lcout(\cemf_module_64ch_ctrl_inst1.N_383 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8_26_LC_17_21_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8_26_LC_17_21_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8_26_LC_17_21_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8_26_LC_17_21_6  (
            .in0(N__39848),
            .in1(N__39863),
            .in2(N__39834),
            .in3(N__39421),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_12_LC_17_22_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_12_LC_17_22_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_12_LC_17_22_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_12_LC_17_22_0  (
            .in0(N__37160),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_state_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65659),
            .ce(),
            .sr(N__62831));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_9_LC_17_22_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_9_LC_17_22_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_9_LC_17_22_1 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_9_LC_17_22_1  (
            .in0(_gnd_net_),
            .in1(N__37159),
            .in2(_gnd_net_),
            .in3(N__37109),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1862 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65659),
            .ce(),
            .sr(N__62831));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_8_LC_17_22_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_8_LC_17_22_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_8_LC_17_22_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_8_LC_17_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37068),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_state_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65659),
            .ce(),
            .sr(N__62831));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_9_LC_17_22_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_9_LC_17_22_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_9_LC_17_22_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_9_LC_17_22_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37049),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65659),
            .ce(),
            .sr(N__62831));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_LC_17_22_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_LC_17_22_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_LC_17_22_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_LC_17_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37020),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65659),
            .ce(),
            .sr(N__62831));
    defparam \serializer_mod_inst.shift_reg_1_LC_17_23_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_1_LC_17_23_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_1_LC_17_23_0 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \serializer_mod_inst.shift_reg_1_LC_17_23_0  (
            .in0(N__44898),
            .in1(N__45427),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\serializer_mod_inst.shift_regZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65674),
            .ce(),
            .sr(N__62824));
    defparam \serializer_mod_inst.shift_reg_12_LC_17_23_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_12_LC_17_23_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_12_LC_17_23_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_12_LC_17_23_1  (
            .in0(_gnd_net_),
            .in1(N__36999),
            .in2(_gnd_net_),
            .in3(N__47857),
            .lcout(\serializer_mod_inst.shift_regZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65674),
            .ce(),
            .sr(N__62824));
    defparam \serializer_mod_inst.shift_reg_49_LC_17_23_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_49_LC_17_23_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_49_LC_17_23_2 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_49_LC_17_23_2  (
            .in0(N__36993),
            .in1(N__45428),
            .in2(_gnd_net_),
            .in3(N__44902),
            .lcout(\serializer_mod_inst.shift_regZ0Z_49 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65674),
            .ce(),
            .sr(N__62824));
    defparam \serializer_mod_inst.shift_reg_91_LC_17_23_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_91_LC_17_23_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_91_LC_17_23_3 .LUT_INIT=16'b0011110000001100;
    LogicCell40 \serializer_mod_inst.shift_reg_91_LC_17_23_3  (
            .in0(_gnd_net_),
            .in1(N__44897),
            .in2(N__45465),
            .in3(N__39915),
            .lcout(\serializer_mod_inst.shift_regZ0Z_91 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65674),
            .ce(),
            .sr(N__62824));
    defparam \serializer_mod_inst.shift_reg_51_LC_17_23_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_51_LC_17_23_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_51_LC_17_23_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \serializer_mod_inst.shift_reg_51_LC_17_23_4  (
            .in0(N__47858),
            .in1(_gnd_net_),
            .in2(N__39930),
            .in3(_gnd_net_),
            .lcout(\serializer_mod_inst.shift_regZ0Z_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65674),
            .ce(),
            .sr(N__62824));
    defparam \serializer_mod_inst.shift_reg_52_LC_17_23_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_52_LC_17_23_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_52_LC_17_23_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_52_LC_17_23_6  (
            .in0(N__47859),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37245),
            .lcout(\serializer_mod_inst.shift_regZ0Z_52 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65674),
            .ce(),
            .sr(N__62824));
    defparam \serializer_mod_inst.shift_reg_10_LC_17_24_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_10_LC_17_24_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_10_LC_17_24_0 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_10_LC_17_24_0  (
            .in0(N__37188),
            .in1(N__45416),
            .in2(_gnd_net_),
            .in3(N__45083),
            .lcout(\serializer_mod_inst.shift_regZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_56_LC_17_24_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_56_LC_17_24_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_56_LC_17_24_1 .LUT_INIT=16'b0011110000001100;
    LogicCell40 \serializer_mod_inst.shift_reg_56_LC_17_24_1  (
            .in0(_gnd_net_),
            .in1(N__44948),
            .in2(N__45463),
            .in3(N__37233),
            .lcout(\serializer_mod_inst.shift_regZ0Z_56 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_15_LC_17_24_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_15_LC_17_24_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_15_LC_17_24_2 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_15_LC_17_24_2  (
            .in0(N__37212),
            .in1(N__45418),
            .in2(_gnd_net_),
            .in3(N__45085),
            .lcout(\serializer_mod_inst.shift_regZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_122_LC_17_24_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_122_LC_17_24_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_122_LC_17_24_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_122_LC_17_24_3  (
            .in0(_gnd_net_),
            .in1(N__37221),
            .in2(_gnd_net_),
            .in3(N__47851),
            .lcout(\serializer_mod_inst.shift_regZ0Z_122 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_14_LC_17_24_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_14_LC_17_24_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_14_LC_17_24_4 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_14_LC_17_24_4  (
            .in0(N__37200),
            .in1(N__45417),
            .in2(_gnd_net_),
            .in3(N__45084),
            .lcout(\serializer_mod_inst.shift_regZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_13_LC_17_24_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_13_LC_17_24_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_13_LC_17_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_13_LC_17_24_5  (
            .in0(N__37206),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__47852),
            .lcout(\serializer_mod_inst.shift_regZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_9_LC_17_24_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_9_LC_17_24_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_9_LC_17_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_9_LC_17_24_7  (
            .in0(_gnd_net_),
            .in1(N__37194),
            .in2(_gnd_net_),
            .in3(N__47853),
            .lcout(\serializer_mod_inst.shift_regZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65683),
            .ce(),
            .sr(N__62819));
    defparam \serializer_mod_inst.shift_reg_18_LC_17_25_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_18_LC_17_25_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_18_LC_17_25_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_18_LC_17_25_0  (
            .in0(N__47850),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37269),
            .lcout(\serializer_mod_inst.shift_regZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65698),
            .ce(),
            .sr(N__62815));
    defparam \serializer_mod_inst.shift_reg_16_LC_17_25_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_16_LC_17_25_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_16_LC_17_25_1 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_16_LC_17_25_1  (
            .in0(N__45066),
            .in1(N__37287),
            .in2(_gnd_net_),
            .in3(N__45407),
            .lcout(\serializer_mod_inst.shift_regZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65698),
            .ce(),
            .sr(N__62815));
    defparam \serializer_mod_inst.shift_reg_80_LC_17_25_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_80_LC_17_25_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_80_LC_17_25_2 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_80_LC_17_25_2  (
            .in0(N__45410),
            .in1(N__37281),
            .in2(_gnd_net_),
            .in3(N__45069),
            .lcout(\serializer_mod_inst.shift_regZ0Z_80 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65698),
            .ce(),
            .sr(N__62815));
    defparam \serializer_mod_inst.shift_reg_108_LC_17_25_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_108_LC_17_25_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_108_LC_17_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_108_LC_17_25_5  (
            .in0(_gnd_net_),
            .in1(N__37257),
            .in2(_gnd_net_),
            .in3(N__47849),
            .lcout(\serializer_mod_inst.shift_regZ0Z_108 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65698),
            .ce(),
            .sr(N__62815));
    defparam \serializer_mod_inst.shift_reg_17_LC_17_25_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_17_LC_17_25_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_17_LC_17_25_6 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_17_LC_17_25_6  (
            .in0(N__45408),
            .in1(N__37275),
            .in2(_gnd_net_),
            .in3(N__45068),
            .lcout(\serializer_mod_inst.shift_regZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65698),
            .ce(),
            .sr(N__62815));
    defparam \serializer_mod_inst.shift_reg_19_LC_17_25_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_19_LC_17_25_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_19_LC_17_25_7 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_19_LC_17_25_7  (
            .in0(N__45067),
            .in1(N__37263),
            .in2(_gnd_net_),
            .in3(N__45409),
            .lcout(\serializer_mod_inst.shift_regZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65698),
            .ce(),
            .sr(N__62815));
    defparam \serializer_mod_inst.shift_reg_107_LC_17_26_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_107_LC_17_26_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_107_LC_17_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_107_LC_17_26_0  (
            .in0(_gnd_net_),
            .in1(N__37353),
            .in2(_gnd_net_),
            .in3(N__47810),
            .lcout(\serializer_mod_inst.shift_regZ0Z_107 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65716),
            .ce(),
            .sr(N__62811));
    defparam \serializer_mod_inst.shift_reg_70_LC_17_26_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_70_LC_17_26_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_70_LC_17_26_1 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_70_LC_17_26_1  (
            .in0(N__45076),
            .in1(N__37251),
            .in2(_gnd_net_),
            .in3(N__45241),
            .lcout(\serializer_mod_inst.shift_regZ0Z_70 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65716),
            .ce(),
            .sr(N__62811));
    defparam \serializer_mod_inst.shift_reg_104_LC_17_26_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_104_LC_17_26_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_104_LC_17_26_3 .LUT_INIT=16'b0101000010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_104_LC_17_26_3  (
            .in0(N__45074),
            .in1(_gnd_net_),
            .in2(N__40158),
            .in3(N__45239),
            .lcout(\serializer_mod_inst.shift_regZ0Z_104 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65716),
            .ce(),
            .sr(N__62811));
    defparam \serializer_mod_inst.shift_reg_106_LC_17_26_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_106_LC_17_26_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_106_LC_17_26_7 .LUT_INIT=16'b0101000010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_106_LC_17_26_7  (
            .in0(N__45075),
            .in1(_gnd_net_),
            .in2(N__37323),
            .in3(N__45240),
            .lcout(\serializer_mod_inst.shift_regZ0Z_106 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65716),
            .ce(),
            .sr(N__62811));
    defparam \serializer_mod_inst.shift_reg_47_LC_17_27_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_47_LC_17_27_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_47_LC_17_27_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_47_LC_17_27_0  (
            .in0(N__47864),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37314),
            .lcout(\serializer_mod_inst.shift_regZ0Z_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65725),
            .ce(),
            .sr(N__62807));
    defparam \serializer_mod_inst.shift_reg_95_LC_17_27_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_95_LC_17_27_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_95_LC_17_27_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_95_LC_17_27_2  (
            .in0(N__45047),
            .in1(N__37335),
            .in2(_gnd_net_),
            .in3(N__45360),
            .lcout(\serializer_mod_inst.shift_regZ0Z_95 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65725),
            .ce(),
            .sr(N__62807));
    defparam \serializer_mod_inst.shift_reg_94_LC_17_27_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_94_LC_17_27_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_94_LC_17_27_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_94_LC_17_27_4  (
            .in0(N__47865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37293),
            .lcout(\serializer_mod_inst.shift_regZ0Z_94 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65725),
            .ce(),
            .sr(N__62807));
    defparam \serializer_mod_inst.shift_reg_105_LC_17_27_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_105_LC_17_27_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_105_LC_17_27_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_105_LC_17_27_5  (
            .in0(_gnd_net_),
            .in1(N__37329),
            .in2(_gnd_net_),
            .in3(N__47863),
            .lcout(\serializer_mod_inst.shift_regZ0Z_105 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65725),
            .ce(),
            .sr(N__62807));
    defparam \serializer_mod_inst.shift_reg_46_LC_17_27_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_46_LC_17_27_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_46_LC_17_27_7 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_46_LC_17_27_7  (
            .in0(N__40272),
            .in1(N__45359),
            .in2(_gnd_net_),
            .in3(N__45048),
            .lcout(\serializer_mod_inst.shift_regZ0Z_46 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65725),
            .ce(),
            .sr(N__62807));
    defparam \serializer_mod_inst.shift_reg_97_LC_17_28_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_97_LC_17_28_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_97_LC_17_28_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_97_LC_17_28_1  (
            .in0(N__37461),
            .in1(N__45442),
            .in2(_gnd_net_),
            .in3(N__45053),
            .lcout(\serializer_mod_inst.shift_regZ0Z_97 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65736),
            .ce(),
            .sr(N__62805));
    defparam \serializer_mod_inst.shift_reg_92_LC_17_28_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_92_LC_17_28_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_92_LC_17_28_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_92_LC_17_28_2  (
            .in0(_gnd_net_),
            .in1(N__37308),
            .in2(_gnd_net_),
            .in3(N__47867),
            .lcout(\serializer_mod_inst.shift_regZ0Z_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65736),
            .ce(),
            .sr(N__62805));
    defparam \serializer_mod_inst.shift_reg_93_LC_17_28_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_93_LC_17_28_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_93_LC_17_28_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_93_LC_17_28_3  (
            .in0(N__47868),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37299),
            .lcout(\serializer_mod_inst.shift_regZ0Z_93 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65736),
            .ce(),
            .sr(N__62805));
    defparam \serializer_mod_inst.shift_reg_96_LC_17_28_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_96_LC_17_28_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_96_LC_17_28_7 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_96_LC_17_28_7  (
            .in0(N__37467),
            .in1(N__45441),
            .in2(_gnd_net_),
            .in3(N__45052),
            .lcout(\serializer_mod_inst.shift_regZ0Z_96 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65736),
            .ce(),
            .sr(N__62805));
    defparam \serializer_mod_inst.shift_reg_98_LC_17_29_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_98_LC_17_29_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_98_LC_17_29_0 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_98_LC_17_29_0  (
            .in0(N__45049),
            .in1(N__37455),
            .in2(_gnd_net_),
            .in3(N__45445),
            .lcout(\serializer_mod_inst.shift_regZ0Z_98 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65745),
            .ce(),
            .sr(N__62804));
    defparam \serializer_mod_inst.enable_config_LC_17_29_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.enable_config_LC_17_29_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.enable_config_LC_17_29_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \serializer_mod_inst.enable_config_LC_17_29_5  (
            .in0(_gnd_net_),
            .in1(N__45443),
            .in2(_gnd_net_),
            .in3(N__45051),
            .lcout(enable_config_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65745),
            .ce(),
            .sr(N__62804));
    defparam \serializer_mod_inst.serial_out_LC_17_29_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.serial_out_LC_17_29_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.serial_out_LC_17_29_6 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \serializer_mod_inst.serial_out_LC_17_29_6  (
            .in0(N__45050),
            .in1(N__44003),
            .in2(_gnd_net_),
            .in3(N__45444),
            .lcout(elec_config_out_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65745),
            .ce(),
            .sr(N__62804));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_24_LC_18_8_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_24_LC_18_8_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_24_LC_18_8_0 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_24_LC_18_8_0  (
            .in0(N__37713),
            .in1(N__51891),
            .in2(N__48537),
            .in3(N__42291),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_24_LC_18_8_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_24_LC_18_8_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_24_LC_18_8_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_24_LC_18_8_1  (
            .in0(N__37422),
            .in1(N__37407),
            .in2(N__37410),
            .in3(N__37359),
            .lcout(I2C_top_level_inst1_s_data_oreg_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65521),
            .ce(N__54506),
            .sr(N__65016));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_24_LC_18_8_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_24_LC_18_8_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_24_LC_18_8_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_24_LC_18_8_2  (
            .in0(N__54222),
            .in1(N__53286),
            .in2(N__40437),
            .in3(N__52989),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_24_LC_18_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_24_LC_18_8_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_24_LC_18_8_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_24_LC_18_8_3  (
            .in0(N__37401),
            .in1(N__52756),
            .in2(N__37383),
            .in3(N__52512),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_24_LC_18_8_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_24_LC_18_8_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_24_LC_18_8_4 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_24_LC_18_8_4  (
            .in0(N__46578),
            .in1(_gnd_net_),
            .in2(N__37362),
            .in3(N__52199),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_23_LC_18_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_23_LC_18_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_23_LC_18_9_0 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_23_LC_18_9_0  (
            .in0(N__37700),
            .in1(N__38311),
            .in2(N__37938),
            .in3(N__49497),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_10_LC_18_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_10_LC_18_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_10_LC_18_9_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_10_LC_18_9_1  (
            .in0(N__37914),
            .in1(N__37699),
            .in2(N__38318),
            .in3(N__42765),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_24_LC_18_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_24_LC_18_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_24_LC_18_9_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_24_LC_18_9_2  (
            .in0(N__37843),
            .in1(N__43584),
            .in2(N__37731),
            .in3(N__64250),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_676 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_0_LC_18_9_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_0_LC_18_9_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_0_LC_18_9_7 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_0_LC_18_9_7  (
            .in0(N__40113),
            .in1(N__37698),
            .in2(N__38317),
            .in3(N__48942),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_23_LC_18_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_23_LC_18_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_23_LC_18_10_0 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_23_LC_18_10_0  (
            .in0(N__51846),
            .in1(N__37557),
            .in2(N__37548),
            .in3(N__49004),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_23_LC_18_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_23_LC_18_10_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_23_LC_18_10_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_23_LC_18_10_1  (
            .in0(N__37524),
            .in1(N__37533),
            .in2(N__37527),
            .in3(N__37473),
            .lcout(I2C_top_level_inst1_s_data_oreg_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65532),
            .ce(N__54498),
            .sr(N__65006));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_23_LC_18_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_23_LC_18_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_23_LC_18_10_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_23_LC_18_10_2  (
            .in0(N__52988),
            .in1(N__48974),
            .in2(N__53306),
            .in3(N__51252),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_23_LC_18_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_23_LC_18_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_23_LC_18_10_3 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_23_LC_18_10_3  (
            .in0(N__37518),
            .in1(N__52738),
            .in2(N__37497),
            .in3(N__52496),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_23_LC_18_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_23_LC_18_10_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_23_LC_18_10_4 .LUT_INIT=16'b0111000001110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_23_LC_18_10_4  (
            .in0(N__49464),
            .in1(N__52191),
            .in2(N__37476),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_20_LC_18_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_20_LC_18_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_20_LC_18_11_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_20_LC_18_11_0  (
            .in0(N__53194),
            .in1(N__42447),
            .in2(N__51915),
            .in3(N__38576),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_21_LC_18_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_21_LC_18_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_21_LC_18_11_1 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_21_LC_18_11_1  (
            .in0(N__45744),
            .in1(N__53195),
            .in2(N__45768),
            .in3(N__51871),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQV592_17_LC_18_11_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQV592_17_LC_18_11_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQV592_17_LC_18_11_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQV592_17_LC_18_11_2  (
            .in0(N__58165),
            .in1(N__58015),
            .in2(N__38577),
            .in3(N__42446),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJJFV5_LC_18_11_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJJFV5_LC_18_11_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJJFV5_LC_18_11_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJJFV5_LC_18_11_3  (
            .in0(N__60353),
            .in1(N__38025),
            .in2(_gnd_net_),
            .in3(N__46086),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21_LC_18_11_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21_LC_18_11_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21_LC_18_11_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21_LC_18_11_4  (
            .in0(_gnd_net_),
            .in1(N__37986),
            .in2(N__38019),
            .in3(N__60187),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net ),
            .ce(N__60009),
            .sr(N__62915));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LH5_LC_18_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LH5_LC_18_11_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LH5_LC_18_11_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LH5_LC_18_11_5  (
            .in0(N__60604),
            .in1(N__40985),
            .in2(N__38016),
            .in3(N__38007),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIEEFV5_LC_18_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIEEFV5_LC_18_11_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIEEFV5_LC_18_11_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIEEFV5_LC_18_11_6  (
            .in0(N__60358),
            .in1(_gnd_net_),
            .in2(N__37998),
            .in3(N__37995),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_20_LC_18_11_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_20_LC_18_11_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_20_LC_18_11_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_20_LC_18_11_7  (
            .in0(N__60186),
            .in1(_gnd_net_),
            .in2(N__37989),
            .in3(N__51525),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net ),
            .ce(N__60009),
            .sr(N__62915));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_21_LC_18_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_21_LC_18_12_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_21_LC_18_12_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_21_LC_18_12_0  (
            .in0(N__37980),
            .in1(N__52755),
            .in2(N__37959),
            .in3(N__52446),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_21_LC_18_12_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_21_LC_18_12_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_21_LC_18_12_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_21_LC_18_12_1  (
            .in0(_gnd_net_),
            .in1(N__52198),
            .in2(N__38397),
            .in3(N__45678),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_21_LC_18_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_21_LC_18_12_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_21_LC_18_12_2 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_21_LC_18_12_2  (
            .in0(N__38394),
            .in1(N__58350),
            .in2(N__44647),
            .in3(N__38375),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_21_LC_18_12_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_21_LC_18_12_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_21_LC_18_12_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_21_LC_18_12_3  (
            .in0(N__38328),
            .in1(N__38222),
            .in2(N__38127),
            .in3(N__45699),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_21_LC_18_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_21_LC_18_12_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_21_LC_18_12_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_21_LC_18_12_4  (
            .in0(N__38124),
            .in1(N__38118),
            .in2(N__38106),
            .in3(N__38103),
            .lcout(I2C_top_level_inst1_s_data_oreg_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65552),
            .ce(N__54496),
            .sr(N__65000));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_12_LC_18_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_12_LC_18_13_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_12_LC_18_13_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_12_LC_18_13_0  (
            .in0(N__59636),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58595),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_21_LC_18_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_21_LC_18_13_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_21_LC_18_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_21_LC_18_13_1  (
            .in0(_gnd_net_),
            .in1(N__59633),
            .in2(_gnd_net_),
            .in3(N__61406),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_30_LC_18_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_30_LC_18_13_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_30_LC_18_13_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_30_LC_18_13_2  (
            .in0(N__59638),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62165),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_13_LC_18_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_13_LC_18_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_13_LC_18_13_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_13_LC_18_13_3  (
            .in0(_gnd_net_),
            .in1(N__59632),
            .in2(_gnd_net_),
            .in3(N__58351),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_22_LC_18_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_22_LC_18_13_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_22_LC_18_13_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_22_LC_18_13_4  (
            .in0(N__59639),
            .in1(N__61352),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_31_LC_18_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_31_LC_18_13_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_31_LC_18_13_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_31_LC_18_13_5  (
            .in0(_gnd_net_),
            .in1(N__59635),
            .in2(_gnd_net_),
            .in3(N__62070),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_14_LC_18_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_14_LC_18_13_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_14_LC_18_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_14_LC_18_13_6  (
            .in0(N__59637),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58498),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_23_LC_18_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_23_LC_18_13_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_23_LC_18_13_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_23_LC_18_13_7  (
            .in0(_gnd_net_),
            .in1(N__59634),
            .in2(_gnd_net_),
            .in3(N__61193),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65564),
            .ce(N__48723),
            .sr(N__62897));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMOSI1_LC_18_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMOSI1_LC_18_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMOSI1_LC_18_14_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMOSI1_LC_18_14_0  (
            .in0(N__55163),
            .in1(N__55423),
            .in2(N__42674),
            .in3(N__38596),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALH5_LC_18_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALH5_LC_18_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALH5_LC_18_14_1 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALH5_LC_18_14_1  (
            .in0(N__60557),
            .in1(N__42277),
            .in2(N__38445),
            .in3(N__38442),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALHZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU3692_17_LC_18_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU3692_17_LC_18_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU3692_17_LC_18_14_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU3692_17_LC_18_14_2  (
            .in0(N__57914),
            .in1(N__58120),
            .in2(N__38429),
            .in3(N__38518),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_22_LC_18_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_22_LC_18_14_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_22_LC_18_14_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_22_LC_18_14_3  (
            .in0(_gnd_net_),
            .in1(N__61353),
            .in2(_gnd_net_),
            .in3(N__59553),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65577),
            .ce(N__49034),
            .sr(N__62886));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0T153_LC_18_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0T153_LC_18_14_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0T153_LC_18_14_4 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0T153_LC_18_14_4  (
            .in0(N__42278),
            .in1(N__46050),
            .in2(N__45915),
            .in3(N__38425),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDD7_LC_18_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDD7_LC_18_14_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDD7_LC_18_14_5 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDD7_LC_18_14_5  (
            .in0(N__38519),
            .in1(N__54005),
            .in2(N__38406),
            .in3(N__38583),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDDZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9U7H2_LC_18_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9U7H2_LC_18_14_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9U7H2_LC_18_14_6 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9U7H2_LC_18_14_6  (
            .in0(N__54798),
            .in1(N__42670),
            .in2(N__55035),
            .in3(N__38597),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_10_LC_18_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_10_LC_18_15_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_10_LC_18_15_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_10_LC_18_15_0  (
            .in0(_gnd_net_),
            .in1(N__59647),
            .in2(_gnd_net_),
            .in3(N__58787),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_11_LC_18_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_11_LC_18_15_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_11_LC_18_15_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_11_LC_18_15_1  (
            .in0(N__59643),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58692),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_20_LC_18_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_20_LC_18_15_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_20_LC_18_15_2 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_20_LC_18_15_2  (
            .in0(N__61530),
            .in1(N__59650),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_12_LC_18_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_12_LC_18_15_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_12_LC_18_15_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_12_LC_18_15_3  (
            .in0(N__59644),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58594),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_21_LC_18_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_21_LC_18_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_21_LC_18_15_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_21_LC_18_15_4  (
            .in0(_gnd_net_),
            .in1(N__59649),
            .in2(_gnd_net_),
            .in3(N__61421),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_30_LC_18_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_30_LC_18_15_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_30_LC_18_15_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_30_LC_18_15_5  (
            .in0(N__59646),
            .in1(N__62179),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_13_LC_18_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_13_LC_18_15_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_13_LC_18_15_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_13_LC_18_15_6  (
            .in0(_gnd_net_),
            .in1(N__59648),
            .in2(_gnd_net_),
            .in3(N__58349),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_22_LC_18_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_22_LC_18_15_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_22_LC_18_15_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_22_LC_18_15_7  (
            .in0(N__59645),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61354),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65587),
            .ce(N__54114),
            .sr(N__62879));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_26_LC_18_16_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_26_LC_18_16_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_26_LC_18_16_0 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_26_LC_18_16_0  (
            .in0(N__56407),
            .in1(N__47546),
            .in2(N__66192),
            .in3(N__56593),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65599),
            .ce(),
            .sr(N__64977));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBDJD_23_LC_18_16_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBDJD_23_LC_18_16_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBDJD_23_LC_18_16_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBDJD_23_LC_18_16_1  (
            .in0(N__57242),
            .in1(N__56406),
            .in2(_gnd_net_),
            .in3(N__56733),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_8_0_m2_ns_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI3S672_1_LC_18_16_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI3S672_1_LC_18_16_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI3S672_1_LC_18_16_2 .LUT_INIT=16'b0000001101000111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI3S672_1_LC_18_16_2  (
            .in0(N__48329),
            .in1(N__56592),
            .in2(N__38709),
            .in3(N__50145),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_322 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_5_LC_18_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_5_LC_18_16_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_5_LC_18_16_3 .LUT_INIT=16'b0000000011011100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_5_LC_18_16_3  (
            .in0(N__47547),
            .in1(N__56949),
            .in2(N__43142),
            .in3(N__66191),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65599),
            .ce(),
            .sr(N__64977));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_6_LC_18_16_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_6_LC_18_16_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_6_LC_18_16_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_6_LC_18_16_4  (
            .in0(N__66187),
            .in1(N__47545),
            .in2(_gnd_net_),
            .in3(N__43135),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65599),
            .ce(),
            .sr(N__64977));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_21_LC_18_16_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_21_LC_18_16_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_21_LC_18_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_21_LC_18_16_5  (
            .in0(_gnd_net_),
            .in1(N__66186),
            .in2(_gnd_net_),
            .in3(N__56916),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65599),
            .ce(),
            .sr(N__64977));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_o2_0_LC_18_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_o2_0_LC_18_16_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_o2_0_LC_18_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_o2_0_LC_18_16_6  (
            .in0(N__56915),
            .in1(N__43134),
            .in2(N__43612),
            .in3(N__56948),
            .lcout(N_1842_0),
            .ltout(N_1842_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.psel_1_N_680_i_i_a2_LC_18_16_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.psel_1_N_680_i_i_a2_LC_18_16_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.psel_1_N_680_i_i_a2_LC_18_16_7 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.psel_1_N_680_i_i_a2_LC_18_16_7  (
            .in0(N__65945),
            .in1(N__56828),
            .in2(N__38682),
            .in3(N__38637),
            .lcout(N_1975),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9_LC_18_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9_LC_18_17_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9_LC_18_17_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9_LC_18_17_0  (
            .in0(N__63045),
            .in1(N__63246),
            .in2(_gnd_net_),
            .in3(N__46524),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C_net ),
            .ce(N__63029),
            .sr(N__62863));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI1SAS1_5_LC_18_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI1SAS1_5_LC_18_17_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI1SAS1_5_LC_18_17_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI1SAS1_5_LC_18_17_1  (
            .in0(N__39513),
            .in1(N__47246),
            .in2(_gnd_net_),
            .in3(N__39106),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI3UAS1_6_LC_18_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI3UAS1_6_LC_18_17_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI3UAS1_6_LC_18_17_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI3UAS1_6_LC_18_17_3  (
            .in0(N__39485),
            .in1(N__47164),
            .in2(_gnd_net_),
            .in3(N__39107),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_addr_RNI3UAS1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI50BS1_7_LC_18_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI50BS1_7_LC_18_17_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI50BS1_7_LC_18_17_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI50BS1_7_LC_18_17_4  (
            .in0(N__39108),
            .in1(N__47093),
            .in2(_gnd_net_),
            .in3(N__39456),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_addr_RNI50BS1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIVPAS1_4_LC_18_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIVPAS1_4_LC_18_17_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIVPAS1_4_LC_18_17_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIVPAS1_4_LC_18_17_5  (
            .in0(N__47196),
            .in1(N__39537),
            .in2(_gnd_net_),
            .in3(N__39105),
            .lcout(\cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_LC_18_18_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_LC_18_18_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_LC_18_18_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_LC_18_18_0  (
            .in0(_gnd_net_),
            .in1(N__39042),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_18_18_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_LUT4_0_LC_18_18_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_LUT4_0_LC_18_18_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_LUT4_0_LC_18_18_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_LUT4_0_LC_18_18_1  (
            .in0(_gnd_net_),
            .in1(N__39282),
            .in2(N__39011),
            .in3(N__38976),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_LUT4_0_LC_18_18_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_LUT4_0_LC_18_18_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_LUT4_0_LC_18_18_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_LUT4_0_LC_18_18_2  (
            .in0(_gnd_net_),
            .in1(N__38960),
            .in2(N__39315),
            .in3(N__38931),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPT1_LC_18_18_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPT1_LC_18_18_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPT1_LC_18_18_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPT1_LC_18_18_3  (
            .in0(_gnd_net_),
            .in1(N__39286),
            .in2(N__38928),
            .in3(N__38835),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQT1_LC_18_18_4 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQT1_LC_18_18_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQT1_LC_18_18_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQT1_LC_18_18_4  (
            .in0(_gnd_net_),
            .in1(N__39253),
            .in2(N__38832),
            .in3(N__38742),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93ST1_LC_18_18_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93ST1_LC_18_18_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93ST1_LC_18_18_5 .LUT_INIT=16'b1100101000110101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93ST1_LC_18_18_5  (
            .in0(N__56147),
            .in1(N__39426),
            .in2(N__39147),
            .in3(N__38739),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93STZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_LC_18_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_LC_18_18_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_LC_18_18_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_LC_18_18_6  (
            .in0(N__39281),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rstZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47984),
            .ce(),
            .sr(N__39174));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNIJHC9_1_LC_18_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNIJHC9_1_LC_18_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNIJHC9_1_LC_18_19_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNIJHC9_1_LC_18_19_1  (
            .in0(_gnd_net_),
            .in1(N__55968),
            .in2(_gnd_net_),
            .in3(N__56352),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_3_LC_18_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_3_LC_18_19_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_3_LC_18_19_2 .LUT_INIT=16'b1010101011110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_3_LC_18_19_2  (
            .in0(N__41385),
            .in1(N__47433),
            .in2(N__39153),
            .in3(N__64570),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_3_LC_18_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_3_LC_18_19_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_3_LC_18_19_3 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_3_LC_18_19_3  (
            .in0(N__54289),
            .in1(N__47384),
            .in2(N__39150),
            .in3(N__42852),
            .lcout(s_paddr_I2C_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65633),
            .ce(N__50080),
            .sr(N__64994));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNO_LC_18_19_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNO_LC_18_19_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNO_LC_18_19_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNO_LC_18_19_4  (
            .in0(N__39564),
            .in1(N__54288),
            .in2(_gnd_net_),
            .in3(N__39133),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_5_LC_18_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_5_LC_18_19_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_5_LC_18_19_5 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_5_LC_18_19_5  (
            .in0(N__64571),
            .in1(N__47382),
            .in2(N__41766),
            .in3(N__43116),
            .lcout(s_paddr_I2C_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65633),
            .ce(N__50080),
            .sr(N__64994));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_6_LC_18_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_6_LC_18_19_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_6_LC_18_19_6 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_6_LC_18_19_6  (
            .in0(N__47381),
            .in1(N__64573),
            .in2(N__41703),
            .in3(N__43101),
            .lcout(s_paddr_I2C_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65633),
            .ce(N__50080),
            .sr(N__64994));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_7_LC_18_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_7_LC_18_19_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_7_LC_18_19_7 .LUT_INIT=16'b1011001110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_7_LC_18_19_7  (
            .in0(N__64572),
            .in1(N__47383),
            .in2(N__41628),
            .in3(N__43086),
            .lcout(s_paddr_I2C_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65633),
            .ce(N__50080),
            .sr(N__64994));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_0_LC_18_20_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_0_LC_18_20_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_0_LC_18_20_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_0_LC_18_20_0  (
            .in0(N__39813),
            .in1(N__39032),
            .in2(_gnd_net_),
            .in3(N__39018),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0 ),
            .ltout(),
            .carryin(bfn_18_20_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_1_LC_18_20_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_1_LC_18_20_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_1_LC_18_20_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_1_LC_18_20_1  (
            .in0(N__39809),
            .in1(N__39646),
            .in2(_gnd_net_),
            .in3(N__39624),
            .lcout(\cemf_module_64ch_ctrl_inst1.paddr_fsm_1 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_2_LC_18_20_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_2_LC_18_20_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_2_LC_18_20_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_2_LC_18_20_2  (
            .in0(N__39814),
            .in1(N__39595),
            .in2(_gnd_net_),
            .in3(N__39579),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_2),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_3_LC_18_20_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_3_LC_18_20_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_3_LC_18_20_3 .LUT_INIT=16'b1011101111101110;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_3_LC_18_20_3  (
            .in0(N__39810),
            .in1(N__39565),
            .in2(_gnd_net_),
            .in3(N__39540),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_3),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_4_LC_18_20_4 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_4_LC_18_20_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_4_LC_18_20_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_4_LC_18_20_4  (
            .in0(N__39815),
            .in1(N__39535),
            .in2(_gnd_net_),
            .in3(N__39516),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_4),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_5_LC_18_20_5 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_5_LC_18_20_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_5_LC_18_20_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_5_LC_18_20_5  (
            .in0(N__39811),
            .in1(N__39505),
            .in2(_gnd_net_),
            .in3(N__39489),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_5),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_6_LC_18_20_6 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_6_LC_18_20_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_6_LC_18_20_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_6_LC_18_20_6  (
            .in0(N__39816),
            .in1(N__39475),
            .in2(_gnd_net_),
            .in3(N__39459),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_6),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_7_LC_18_20_7 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_7_LC_18_20_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_7_LC_18_20_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_7_LC_18_20_7  (
            .in0(N__39812),
            .in1(N__39448),
            .in2(_gnd_net_),
            .in3(N__39429),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7 ),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_7 ),
            .clk(N__65649),
            .ce(N__39696),
            .sr(N__62847));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_8_LC_18_21_0 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_8_LC_18_21_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_8_LC_18_21_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_8_LC_18_21_0  (
            .in0(N__39799),
            .in1(N__39425),
            .in2(_gnd_net_),
            .in3(N__39405),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_8),
            .ltout(),
            .carryin(bfn_18_21_0_),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_9_LC_18_21_1 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_9_LC_18_21_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_9_LC_18_21_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_9_LC_18_21_1  (
            .in0(N__39794),
            .in1(N__39909),
            .in2(_gnd_net_),
            .in3(N__39897),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_9),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_10_LC_18_21_2 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_10_LC_18_21_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_10_LC_18_21_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_10_LC_18_21_2  (
            .in0(N__39796),
            .in1(N__39894),
            .in2(_gnd_net_),
            .in3(N__39882),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_10),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_11_LC_18_21_3 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_11_LC_18_21_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_11_LC_18_21_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_11_LC_18_21_3  (
            .in0(N__39792),
            .in1(N__39879),
            .in2(_gnd_net_),
            .in3(N__39867),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_11),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_12_LC_18_21_4 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_12_LC_18_21_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_12_LC_18_21_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_12_LC_18_21_4  (
            .in0(N__39797),
            .in1(N__39864),
            .in2(_gnd_net_),
            .in3(N__39852),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_12),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_13_LC_18_21_5 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_13_LC_18_21_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_13_LC_18_21_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_13_LC_18_21_5  (
            .in0(N__39793),
            .in1(N__39849),
            .in2(_gnd_net_),
            .in3(N__39837),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_13),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_14_LC_18_21_6 .C_ON=1'b1;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_14_LC_18_21_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_14_LC_18_21_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_14_LC_18_21_6  (
            .in0(N__39798),
            .in1(N__39833),
            .in2(_gnd_net_),
            .in3(N__39819),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_14),
            .ltout(),
            .carryin(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13 ),
            .carryout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_14 ),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_15_LC_18_21_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_15_LC_18_21_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_15_LC_18_21_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_15_LC_18_21_7  (
            .in0(N__39795),
            .in1(N__39710),
            .in2(_gnd_net_),
            .in3(N__39714),
            .lcout(cemf_module_64ch_ctrl_inst1_paddr_fsm_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65660),
            .ce(N__39695),
            .sr(N__62841));
    defparam \serializer_mod_inst.shift_reg_86_LC_18_22_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_86_LC_18_22_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_86_LC_18_22_0 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \serializer_mod_inst.shift_reg_86_LC_18_22_0  (
            .in0(N__47873),
            .in1(N__40197),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\serializer_mod_inst.shift_regZ0Z_86 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65675),
            .ce(),
            .sr(N__62835));
    defparam \serializer_mod_inst.shift_reg_87_LC_18_22_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_87_LC_18_22_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_87_LC_18_22_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_87_LC_18_22_2  (
            .in0(N__44929),
            .in1(N__39666),
            .in2(_gnd_net_),
            .in3(N__45459),
            .lcout(\serializer_mod_inst.shift_regZ0Z_87 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65675),
            .ce(),
            .sr(N__62835));
    defparam \serializer_mod_inst.shift_reg_54_LC_18_22_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_54_LC_18_22_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_54_LC_18_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_54_LC_18_22_3  (
            .in0(_gnd_net_),
            .in1(N__39957),
            .in2(_gnd_net_),
            .in3(N__47872),
            .lcout(\serializer_mod_inst.shift_regZ0Z_54 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65675),
            .ce(),
            .sr(N__62835));
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_6_LC_18_22_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_6_LC_18_22_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_6_LC_18_22_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_6_LC_18_22_5  (
            .in0(N__40112),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40033),
            .lcout(\cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65675),
            .ce(),
            .sr(N__62835));
    defparam \serializer_mod_inst.shift_reg_53_LC_18_22_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_53_LC_18_22_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_53_LC_18_22_7 .LUT_INIT=16'b0101010110100000;
    LogicCell40 \serializer_mod_inst.shift_reg_53_LC_18_22_7  (
            .in0(N__45458),
            .in1(_gnd_net_),
            .in2(N__39966),
            .in3(N__44930),
            .lcout(\serializer_mod_inst.shift_regZ0Z_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65675),
            .ce(),
            .sr(N__62835));
    defparam \serializer_mod_inst.shift_reg_88_LC_18_23_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_88_LC_18_23_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_88_LC_18_23_0 .LUT_INIT=16'b0011000011001100;
    LogicCell40 \serializer_mod_inst.shift_reg_88_LC_18_23_0  (
            .in0(_gnd_net_),
            .in1(N__45065),
            .in2(N__39951),
            .in3(N__45391),
            .lcout(\serializer_mod_inst.shift_regZ0Z_88 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65684),
            .ce(),
            .sr(N__62832));
    defparam \serializer_mod_inst.shift_reg_101_LC_18_23_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_101_LC_18_23_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_101_LC_18_23_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_101_LC_18_23_1  (
            .in0(N__40131),
            .in1(N__45390),
            .in2(_gnd_net_),
            .in3(N__45082),
            .lcout(\serializer_mod_inst.shift_regZ0Z_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65684),
            .ce(),
            .sr(N__62832));
    defparam \serializer_mod_inst.shift_reg_89_LC_18_23_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_89_LC_18_23_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_89_LC_18_23_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_89_LC_18_23_4  (
            .in0(_gnd_net_),
            .in1(N__39942),
            .in2(_gnd_net_),
            .in3(N__47855),
            .lcout(\serializer_mod_inst.shift_regZ0Z_89 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65684),
            .ce(),
            .sr(N__62832));
    defparam \serializer_mod_inst.shift_reg_50_LC_18_23_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_50_LC_18_23_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_50_LC_18_23_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_50_LC_18_23_6  (
            .in0(_gnd_net_),
            .in1(N__39936),
            .in2(_gnd_net_),
            .in3(N__47854),
            .lcout(\serializer_mod_inst.shift_regZ0Z_50 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65684),
            .ce(),
            .sr(N__62832));
    defparam \serializer_mod_inst.shift_reg_90_LC_18_23_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_90_LC_18_23_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_90_LC_18_23_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_90_LC_18_23_7  (
            .in0(N__47856),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__39921),
            .lcout(\serializer_mod_inst.shift_regZ0Z_90 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65684),
            .ce(),
            .sr(N__62832));
    defparam \serializer_mod_inst.shift_reg_85_LC_18_24_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_85_LC_18_24_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_85_LC_18_24_0 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_85_LC_18_24_0  (
            .in0(N__45071),
            .in1(N__40146),
            .in2(_gnd_net_),
            .in3(N__45451),
            .lcout(\serializer_mod_inst.shift_regZ0Z_85 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65699),
            .ce(),
            .sr(N__62825));
    defparam \serializer_mod_inst.shift_reg_2_LC_18_24_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_2_LC_18_24_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_2_LC_18_24_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_2_LC_18_24_2  (
            .in0(N__45070),
            .in1(N__40188),
            .in2(_gnd_net_),
            .in3(N__45449),
            .lcout(\serializer_mod_inst.shift_regZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65699),
            .ce(),
            .sr(N__62825));
    defparam \serializer_mod_inst.shift_reg_102_LC_18_24_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_102_LC_18_24_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_102_LC_18_24_3 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_102_LC_18_24_3  (
            .in0(N__45448),
            .in1(N__40182),
            .in2(_gnd_net_),
            .in3(N__45072),
            .lcout(\serializer_mod_inst.shift_regZ0Z_102 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65699),
            .ce(),
            .sr(N__62825));
    defparam \serializer_mod_inst.shift_reg_66_LC_18_24_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_66_LC_18_24_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_66_LC_18_24_5 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_66_LC_18_24_5  (
            .in0(N__45450),
            .in1(N__44019),
            .in2(_gnd_net_),
            .in3(N__45073),
            .lcout(\serializer_mod_inst.shift_regZ0Z_66 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65699),
            .ce(),
            .sr(N__62825));
    defparam \serializer_mod_inst.shift_reg_103_LC_18_24_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_103_LC_18_24_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_103_LC_18_24_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_103_LC_18_24_7  (
            .in0(_gnd_net_),
            .in1(N__40164),
            .in2(_gnd_net_),
            .in3(N__47848),
            .lcout(\serializer_mod_inst.shift_regZ0Z_103 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65699),
            .ce(),
            .sr(N__62825));
    defparam \serializer_mod_inst.shift_reg_44_LC_18_25_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_44_LC_18_25_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_44_LC_18_25_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_44_LC_18_25_1  (
            .in0(_gnd_net_),
            .in1(N__40284),
            .in2(_gnd_net_),
            .in3(N__47845),
            .lcout(\serializer_mod_inst.shift_regZ0Z_44 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_84_LC_18_25_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_84_LC_18_25_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_84_LC_18_25_2 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \serializer_mod_inst.shift_reg_84_LC_18_25_2  (
            .in0(N__47847),
            .in1(_gnd_net_),
            .in2(N__40206),
            .in3(_gnd_net_),
            .lcout(\serializer_mod_inst.shift_regZ0Z_84 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_22_LC_18_25_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_22_LC_18_25_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_22_LC_18_25_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_22_LC_18_25_3  (
            .in0(_gnd_net_),
            .in1(N__41814),
            .in2(_gnd_net_),
            .in3(N__47843),
            .lcout(\serializer_mod_inst.shift_regZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_42_LC_18_25_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_42_LC_18_25_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_42_LC_18_25_4 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_42_LC_18_25_4  (
            .in0(N__40140),
            .in1(N__45447),
            .in2(_gnd_net_),
            .in3(N__45086),
            .lcout(\serializer_mod_inst.shift_regZ0Z_42 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_100_LC_18_25_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_100_LC_18_25_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_100_LC_18_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_100_LC_18_25_5  (
            .in0(_gnd_net_),
            .in1(N__40227),
            .in2(_gnd_net_),
            .in3(N__47842),
            .lcout(\serializer_mod_inst.shift_regZ0Z_100 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_43_LC_18_25_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_43_LC_18_25_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_43_LC_18_25_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_43_LC_18_25_6  (
            .in0(N__47844),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40290),
            .lcout(\serializer_mod_inst.shift_regZ0Z_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_45_LC_18_25_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_45_LC_18_25_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_45_LC_18_25_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_45_LC_18_25_7  (
            .in0(_gnd_net_),
            .in1(N__40278),
            .in2(_gnd_net_),
            .in3(N__47846),
            .lcout(\serializer_mod_inst.shift_regZ0Z_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65717),
            .ce(),
            .sr(N__62820));
    defparam \serializer_mod_inst.shift_reg_72_LC_18_26_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_72_LC_18_26_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_72_LC_18_26_0 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_72_LC_18_26_0  (
            .in0(N__45077),
            .in1(N__40257),
            .in2(_gnd_net_),
            .in3(N__45245),
            .lcout(\serializer_mod_inst.shift_regZ0Z_72 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_71_LC_18_26_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_71_LC_18_26_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_71_LC_18_26_1 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_71_LC_18_26_1  (
            .in0(N__40263),
            .in1(N__45242),
            .in2(_gnd_net_),
            .in3(N__45079),
            .lcout(\serializer_mod_inst.shift_regZ0Z_71 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_74_LC_18_26_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_74_LC_18_26_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_74_LC_18_26_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_74_LC_18_26_2  (
            .in0(N__45078),
            .in1(N__40212),
            .in2(_gnd_net_),
            .in3(N__45246),
            .lcout(\serializer_mod_inst.shift_regZ0Z_74 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_75_LC_18_26_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_75_LC_18_26_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_75_LC_18_26_3 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_75_LC_18_26_3  (
            .in0(N__40251),
            .in1(N__45243),
            .in2(_gnd_net_),
            .in3(N__45080),
            .lcout(\serializer_mod_inst.shift_regZ0Z_75 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_99_LC_18_26_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_99_LC_18_26_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_99_LC_18_26_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_99_LC_18_26_4  (
            .in0(N__47742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__40236),
            .lcout(\serializer_mod_inst.shift_regZ0Z_99 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_73_LC_18_26_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_73_LC_18_26_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_73_LC_18_26_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_73_LC_18_26_5  (
            .in0(_gnd_net_),
            .in1(N__47741),
            .in2(_gnd_net_),
            .in3(N__40218),
            .lcout(\serializer_mod_inst.shift_regZ0Z_73 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_83_LC_18_26_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_83_LC_18_26_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_83_LC_18_26_7 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_83_LC_18_26_7  (
            .in0(N__40422),
            .in1(N__45244),
            .in2(_gnd_net_),
            .in3(N__45081),
            .lcout(\serializer_mod_inst.shift_regZ0Z_83 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65726),
            .ce(),
            .sr(N__62816));
    defparam \serializer_mod_inst.shift_reg_82_LC_18_28_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_82_LC_18_28_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_82_LC_18_28_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_82_LC_18_28_1  (
            .in0(_gnd_net_),
            .in1(N__40401),
            .in2(_gnd_net_),
            .in3(N__47866),
            .lcout(\serializer_mod_inst.shift_regZ0Z_82 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65746),
            .ce(),
            .sr(N__62808));
    defparam \serializer_mod_inst.shift_reg_81_LC_18_28_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_81_LC_18_28_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_81_LC_18_28_2 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_81_LC_18_28_2  (
            .in0(N__40413),
            .in1(N__45457),
            .in2(_gnd_net_),
            .in3(N__45089),
            .lcout(\serializer_mod_inst.shift_regZ0Z_81 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65746),
            .ce(),
            .sr(N__62808));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_27_LC_19_8_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_27_LC_19_8_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_27_LC_19_8_4 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_27_LC_19_8_4  (
            .in0(N__53008),
            .in1(N__51279),
            .in2(N__40584),
            .in3(N__53282),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_29_LC_19_9_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_29_LC_19_9_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_29_LC_19_9_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_29_LC_19_9_0  (
            .in0(N__51264),
            .in1(N__53296),
            .in2(N__59748),
            .in3(N__52999),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_29_LC_19_9_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_29_LC_19_9_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_29_LC_19_9_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_29_LC_19_9_1  (
            .in0(N__40395),
            .in1(N__52770),
            .in2(N__40374),
            .in3(N__52485),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_29_LC_19_9_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_29_LC_19_9_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_29_LC_19_9_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_29_LC_19_9_2  (
            .in0(_gnd_net_),
            .in1(N__49110),
            .in2(N__40353),
            .in3(N__52214),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_29_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_29_LC_19_9_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_29_LC_19_9_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_29_LC_19_9_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_29_LC_19_9_3  (
            .in0(N__40350),
            .in1(N__40335),
            .in2(N__40329),
            .in3(N__40296),
            .lcout(I2C_top_level_inst1_s_data_oreg_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65533),
            .ce(N__54499),
            .sr(N__65017));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_29_LC_19_9_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_29_LC_19_9_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_29_LC_19_9_4 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_29_LC_19_9_4  (
            .in0(N__40326),
            .in1(N__51890),
            .in2(N__48774),
            .in3(N__40311),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI4TB92_17_LC_19_10_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI4TB92_17_LC_19_10_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI4TB92_17_LC_19_10_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI4TB92_17_LC_19_10_0  (
            .in0(N__58016),
            .in1(N__58185),
            .in2(N__40530),
            .in3(N__48749),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6VB92_17_LC_19_10_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6VB92_17_LC_19_10_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6VB92_17_LC_19_10_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6VB92_17_LC_19_10_1  (
            .in0(N__58186),
            .in1(N__58017),
            .in2(N__40773),
            .in3(N__40696),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3Q5_LC_19_10_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3Q5_LC_19_10_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3Q5_LC_19_10_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3Q5_LC_19_10_2  (
            .in0(N__60591),
            .in1(N__40717),
            .in2(N__40491),
            .in3(N__40782),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNISCU76_LC_19_10_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNISCU76_LC_19_10_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNISCU76_LC_19_10_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNISCU76_LC_19_10_3  (
            .in0(_gnd_net_),
            .in1(N__60357),
            .in2(N__40488),
            .in3(N__40485),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8_LC_19_10_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8_LC_19_10_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8_LC_19_10_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8_LC_19_10_4  (
            .in0(N__60203),
            .in1(_gnd_net_),
            .in2(N__40479),
            .in3(N__40443),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net ),
            .ce(N__59994),
            .sr(N__62933));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3Q5_LC_19_10_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3Q5_LC_19_10_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3Q5_LC_19_10_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3Q5_LC_19_10_5  (
            .in0(N__60517),
            .in1(N__45529),
            .in2(N__40476),
            .in3(N__40569),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIN7U76_LC_19_10_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIN7U76_LC_19_10_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIN7U76_LC_19_10_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIN7U76_LC_19_10_6  (
            .in0(N__60356),
            .in1(_gnd_net_),
            .in2(N__40467),
            .in3(N__40464),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_7_LC_19_10_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_7_LC_19_10_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_7_LC_19_10_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_7_LC_19_10_7  (
            .in0(N__40458),
            .in1(_gnd_net_),
            .in2(N__40446),
            .in3(N__60202),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net ),
            .ce(N__59994),
            .sr(N__62933));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_24_LC_19_11_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_24_LC_19_11_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_24_LC_19_11_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_24_LC_19_11_0  (
            .in0(N__61125),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59702),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_16_LC_19_11_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_16_LC_19_11_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_16_LC_19_11_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_16_LC_19_11_1  (
            .in0(N__59696),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57601),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_28_LC_19_11_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_28_LC_19_11_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_28_LC_19_11_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_28_LC_19_11_2  (
            .in0(N__62369),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59704),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_8_LC_19_11_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_8_LC_19_11_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_8_LC_19_11_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_8_LC_19_11_3  (
            .in0(N__63149),
            .in1(_gnd_net_),
            .in2(N__59728),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_26_LC_19_11_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_26_LC_19_11_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_26_LC_19_11_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_26_LC_19_11_4  (
            .in0(_gnd_net_),
            .in1(N__59695),
            .in2(_gnd_net_),
            .in3(N__60914),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_1Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_18_LC_19_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_18_LC_19_11_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_18_LC_19_11_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_18_LC_19_11_5  (
            .in0(N__59697),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59852),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_27_LC_19_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_27_LC_19_11_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_27_LC_19_11_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_27_LC_19_11_6  (
            .in0(N__60776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59703),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_1_LC_19_11_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_1_LC_19_11_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_1_LC_19_11_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_1_LC_19_11_7  (
            .in0(N__59698),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61859),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65553),
            .ce(N__58879),
            .sr(N__62924));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISGFN1_LC_19_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISGFN1_LC_19_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISGFN1_LC_19_12_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISGFN1_LC_19_12_0  (
            .in0(N__55256),
            .in1(N__55447),
            .in2(N__41053),
            .in3(N__40543),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIFMQL2_LC_19_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIFMQL2_LC_19_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIFMQL2_LC_19_12_1 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIFMQL2_LC_19_12_1  (
            .in0(N__40544),
            .in1(N__55031),
            .in2(N__41054),
            .in3(N__54820),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_7_LC_19_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_7_LC_19_12_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_7_LC_19_12_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_7_LC_19_12_2  (
            .in0(N__59706),
            .in1(N__63476),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65565),
            .ce(N__49083),
            .sr(N__62916));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISSQI1_LC_19_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISSQI1_LC_19_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISSQI1_LC_19_12_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISSQI1_LC_19_12_3  (
            .in0(N__55446),
            .in1(N__55257),
            .in2(N__42010),
            .in3(N__42577),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_16_LC_19_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_16_LC_19_12_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_16_LC_19_12_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_16_LC_19_12_4  (
            .in0(N__59705),
            .in1(N__57619),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65565),
            .ce(N__49083),
            .sr(N__62916));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIF26H2_LC_19_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIF26H2_LC_19_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIF26H2_LC_19_12_5 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIF26H2_LC_19_12_5  (
            .in0(N__54963),
            .in1(N__54819),
            .in2(N__42011),
            .in3(N__42578),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUIFN1_LC_19_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUIFN1_LC_19_12_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUIFN1_LC_19_12_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUIFN1_LC_19_12_6  (
            .in0(N__55258),
            .in1(N__55448),
            .in2(N__41021),
            .in3(N__40822),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_8_LC_19_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_8_LC_19_12_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_8_LC_19_12_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_8_LC_19_12_7  (
            .in0(_gnd_net_),
            .in1(N__59707),
            .in2(_gnd_net_),
            .in3(N__63150),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65565),
            .ce(N__49083),
            .sr(N__62916));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI8NK93_LC_19_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI8NK93_LC_19_13_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI8NK93_LC_19_13_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI8NK93_LC_19_13_0  (
            .in0(N__45869),
            .in1(N__40766),
            .in2(N__46068),
            .in3(N__40721),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SL7_LC_19_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SL7_LC_19_13_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SL7_LC_19_13_1 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SL7_LC_19_13_1  (
            .in0(N__54004),
            .in1(N__40697),
            .in2(N__40653),
            .in3(N__40806),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIR9DO7_LC_19_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIR9DO7_LC_19_13_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIR9DO7_LC_19_13_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIR9DO7_LC_19_13_2  (
            .in0(_gnd_net_),
            .in1(N__53690),
            .in2(N__40650),
            .in3(N__40647),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8_LC_19_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8_LC_19_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8_LC_19_13_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8_LC_19_13_3  (
            .in0(_gnd_net_),
            .in1(N__40641),
            .in2(N__40626),
            .in3(N__55723),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net ),
            .ce(N__55539),
            .sr(N__62908));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISLPF7_LC_19_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISLPF7_LC_19_13_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISLPF7_LC_19_13_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISLPF7_LC_19_13_4  (
            .in0(N__40842),
            .in1(N__53689),
            .in2(_gnd_net_),
            .in3(N__40851),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_14_LC_19_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_14_LC_19_13_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_14_LC_19_13_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_14_LC_19_13_5  (
            .in0(_gnd_net_),
            .in1(N__41139),
            .in2(N__40836),
            .in3(N__55722),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net ),
            .ce(N__55539),
            .sr(N__62908));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIHOQL2_LC_19_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIHOQL2_LC_19_13_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIHOQL2_LC_19_13_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIHOQL2_LC_19_13_6  (
            .in0(N__55030),
            .in1(N__54821),
            .in2(N__41020),
            .in3(N__40823),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQKV43_LC_19_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQKV43_LC_19_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQKV43_LC_19_14_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQKV43_LC_19_14_0  (
            .in0(N__45871),
            .in1(N__46042),
            .in2(N__49255),
            .in3(N__49285),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISAK93_LC_19_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISAK93_LC_19_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISAK93_LC_19_14_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISAK93_LC_19_14_1  (
            .in0(N__46043),
            .in1(N__45872),
            .in2(N__49747),
            .in3(N__49948),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISO153_LC_19_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISO153_LC_19_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISO153_LC_19_14_2 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISO153_LC_19_14_2  (
            .in0(N__45873),
            .in1(N__46045),
            .in2(N__42445),
            .in3(N__40973),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUCK93_LC_19_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUCK93_LC_19_14_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUCK93_LC_19_14_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUCK93_LC_19_14_3  (
            .in0(N__46044),
            .in1(N__45874),
            .in2(N__49636),
            .in3(N__49693),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUOV43_LC_19_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUOV43_LC_19_14_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUOV43_LC_19_14_4 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUOV43_LC_19_14_4  (
            .in0(N__45875),
            .in1(N__46046),
            .in2(N__41197),
            .in3(N__46339),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_10_LC_19_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_10_LC_19_14_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_10_LC_19_14_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_10_LC_19_14_5  (
            .in0(_gnd_net_),
            .in1(N__59640),
            .in2(_gnd_net_),
            .in3(N__58788),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65588),
            .ce(N__58867),
            .sr(N__62898));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_2_LC_19_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_2_LC_19_14_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_2_LC_19_14_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_2_LC_19_14_6  (
            .in0(N__59642),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61737),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65588),
            .ce(N__58867),
            .sr(N__62898));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_20_LC_19_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_20_LC_19_14_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_20_LC_19_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_20_LC_19_14_7  (
            .in0(_gnd_net_),
            .in1(N__59641),
            .in2(_gnd_net_),
            .in3(N__61531),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65588),
            .ce(N__58867),
            .sr(N__62898));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKKQI1_LC_19_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKKQI1_LC_19_15_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKKQI1_LC_19_15_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKKQI1_LC_19_15_0  (
            .in0(N__55250),
            .in1(N__55409),
            .in2(N__42701),
            .in3(N__40957),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7Q5H2_LC_19_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7Q5H2_LC_19_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7Q5H2_LC_19_15_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7Q5H2_LC_19_15_1  (
            .in0(N__55029),
            .in1(N__54783),
            .in2(N__40962),
            .in3(N__42697),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_0_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI788D7_LC_19_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI788D7_LC_19_15_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI788D7_LC_19_15_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI788D7_LC_19_15_2  (
            .in0(N__54001),
            .in1(N__41221),
            .in2(N__40935),
            .in3(N__40932),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_0_i_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIBPF7_LC_19_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIBPF7_LC_19_15_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIBPF7_LC_19_15_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIBPF7_LC_19_15_3  (
            .in0(_gnd_net_),
            .in1(N__53712),
            .in2(N__40926),
            .in3(N__40923),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12_LC_19_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12_LC_19_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12_LC_19_15_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12_LC_19_15_4  (
            .in0(_gnd_net_),
            .in1(N__46101),
            .in2(N__40917),
            .in3(N__55695),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net ),
            .ce(N__55538),
            .sr(N__62887));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8D7_LC_19_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8D7_LC_19_15_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8D7_LC_19_15_5 .LUT_INIT=16'b0111010111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8D7_LC_19_15_5  (
            .in0(N__40914),
            .in1(N__54002),
            .in2(N__40892),
            .in3(N__42819),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINGPF7_LC_19_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINGPF7_LC_19_15_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINGPF7_LC_19_15_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINGPF7_LC_19_15_6  (
            .in0(N__53713),
            .in1(_gnd_net_),
            .in2(N__40860),
            .in3(N__40857),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_13_LC_19_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_13_LC_19_15_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_13_LC_19_15_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_13_LC_19_15_7  (
            .in0(N__55696),
            .in1(_gnd_net_),
            .in2(N__41148),
            .in3(N__41145),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net ),
            .ce(N__55538),
            .sr(N__62887));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_1_LC_19_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_1_LC_19_16_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_1_LC_19_16_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_1_LC_19_16_0  (
            .in0(N__59546),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61871),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_2_LC_19_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_2_LC_19_16_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_2_LC_19_16_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_2_LC_19_16_1  (
            .in0(N__61738),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59550),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_5_LC_19_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_5_LC_19_16_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_5_LC_19_16_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_5_LC_19_16_2  (
            .in0(N__59547),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63702),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_6_LC_19_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_6_LC_19_16_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_6_LC_19_16_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_6_LC_19_16_3  (
            .in0(N__63584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59551),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_7_LC_19_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_7_LC_19_16_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_7_LC_19_16_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_7_LC_19_16_4  (
            .in0(N__59548),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63471),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_8_LC_19_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_8_LC_19_16_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_8_LC_19_16_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_8_LC_19_16_5  (
            .in0(_gnd_net_),
            .in1(N__59552),
            .in2(_gnd_net_),
            .in3(N__63145),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_9_LC_19_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_9_LC_19_16_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_9_LC_19_16_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_9_LC_19_16_6  (
            .in0(N__59549),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46523),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_10_LC_19_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_10_LC_19_16_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_10_LC_19_16_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_10_LC_19_16_7  (
            .in0(_gnd_net_),
            .in1(N__58779),
            .in2(_gnd_net_),
            .in3(N__59545),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65608),
            .ce(N__45567),
            .sr(N__62880));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIE9AV5_LC_19_17_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIE9AV5_LC_19_17_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIE9AV5_LC_19_17_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIE9AV5_LC_19_17_0  (
            .in0(N__60345),
            .in1(N__41292),
            .in2(_gnd_net_),
            .in3(N__41154),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11_LC_19_17_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11_LC_19_17_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11_LC_19_17_1 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11_LC_19_17_1  (
            .in0(_gnd_net_),
            .in1(N__49857),
            .in2(N__41286),
            .in3(N__60164),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net ),
            .ce(N__59984),
            .sr(N__62871));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GH5_LC_19_17_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GH5_LC_19_17_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GH5_LC_19_17_2 .LUT_INIT=16'b0111111101011111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GH5_LC_19_17_2  (
            .in0(N__41283),
            .in1(N__60516),
            .in2(N__41169),
            .in3(N__46346),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJEAV5_LC_19_17_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJEAV5_LC_19_17_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJEAV5_LC_19_17_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJEAV5_LC_19_17_3  (
            .in0(_gnd_net_),
            .in1(N__60346),
            .in2(N__41274),
            .in3(N__41271),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_12_LC_19_17_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_12_LC_19_17_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_12_LC_19_17_4 .LUT_INIT=16'b1101100011011000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_12_LC_19_17_4  (
            .in0(N__60165),
            .in1(N__41265),
            .in2(N__41259),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net ),
            .ce(N__59984),
            .sr(N__62871));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISV392_17_LC_19_17_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISV392_17_LC_19_17_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISV392_17_LC_19_17_5 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISV392_17_LC_19_17_5  (
            .in0(N__58158),
            .in1(N__57980),
            .in2(N__41238),
            .in3(N__41201),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQT392_17_LC_19_17_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQT392_17_LC_19_17_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQT392_17_LC_19_17_6 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQT392_17_LC_19_17_6  (
            .in0(N__57979),
            .in1(N__58159),
            .in2(N__42528),
            .in3(N__42554),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFH5_LC_19_17_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFH5_LC_19_17_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFH5_LC_19_17_7 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFH5_LC_19_17_7  (
            .in0(N__60515),
            .in1(N__46376),
            .in2(N__41157),
            .in3(N__42921),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFHZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIR9FE1_9_LC_19_18_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIR9FE1_9_LC_19_18_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIR9FE1_9_LC_19_18_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIR9FE1_9_LC_19_18_0  (
            .in0(N__46938),
            .in1(N__47042),
            .in2(N__56440),
            .in3(N__47007),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_7_3_i_a2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_10_LC_19_18_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_10_LC_19_18_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_10_LC_19_18_2 .LUT_INIT=16'b1100000010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_10_LC_19_18_2  (
            .in0(N__43059),
            .in1(N__41304),
            .in2(N__64584),
            .in3(N__47380),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65634),
            .ce(N__50076),
            .sr(N__64995));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_4_LC_19_18_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_4_LC_19_18_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_4_LC_19_18_3 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_4_LC_19_18_3  (
            .in0(N__47378),
            .in1(N__64582),
            .in2(N__41328),
            .in3(N__42837),
            .lcout(s_paddr_I2C_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65634),
            .ce(N__50076),
            .sr(N__64995));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_11_LC_19_18_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_11_LC_19_18_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_11_LC_19_18_4 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_11_LC_19_18_4  (
            .in0(N__64581),
            .in1(N__41298),
            .in2(N__47403),
            .in3(N__43050),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65634),
            .ce(N__50076),
            .sr(N__64995));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_9_LC_19_18_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_9_LC_19_18_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_9_LC_19_18_5 .LUT_INIT=16'b1101010110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_9_LC_19_18_5  (
            .in0(N__47379),
            .in1(N__64583),
            .in2(N__41313),
            .in3(N__43068),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65634),
            .ce(N__50076),
            .sr(N__64995));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIIP1Q6_13_LC_19_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIIP1Q6_13_LC_19_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIIP1Q6_13_LC_19_18_6 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIIP1Q6_13_LC_19_18_6  (
            .in0(N__64713),
            .in1(N__55794),
            .in2(N__56250),
            .in3(N__55988),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_0_LC_19_18_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_0_LC_19_18_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_0_LC_19_18_7 .LUT_INIT=16'b1100010111001010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_0_LC_19_18_7  (
            .in0(N__55989),
            .in1(N__64485),
            .in2(N__41316),
            .in3(N__46756),
            .lcout(s_paddr_I2C_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65634),
            .ce(N__50076),
            .sr(N__64995));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_0_LC_19_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_0_LC_19_19_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_0_LC_19_19_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_0_LC_19_19_0  (
            .in0(N__48292),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.s_addr1_o_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_1_LC_19_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_1_LC_19_19_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_1_LC_19_19_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_1_LC_19_19_1  (
            .in0(N__48157),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.s_addr1_o_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_2_LC_19_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_2_LC_19_19_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_2_LC_19_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_2_LC_19_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48106),
            .lcout(\I2C_top_level_inst1.s_addr1_o_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_3_LC_19_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_3_LC_19_19_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_3_LC_19_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_3_LC_19_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48048),
            .lcout(\I2C_top_level_inst1.s_addr1_o_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_4_LC_19_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_4_LC_19_19_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_4_LC_19_19_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_4_LC_19_19_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41378),
            .lcout(\I2C_top_level_inst1.s_addr1_o_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_5_LC_19_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_5_LC_19_19_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_5_LC_19_19_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_5_LC_19_19_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41807),
            .lcout(\I2C_top_level_inst1.s_addr1_o_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_6_LC_19_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_6_LC_19_19_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_6_LC_19_19_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_6_LC_19_19_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41752),
            .lcout(\I2C_top_level_inst1.s_addr1_o_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_7_LC_19_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_7_LC_19_19_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr1_reg_inst.c_addr1_7_LC_19_19_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr1_reg_inst.c_addr1_7_LC_19_19_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41690),
            .lcout(\I2C_top_level_inst1.s_addr1_o_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47990),
            .ce(N__41420),
            .sr(N__62859));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_0_LC_19_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_0_LC_19_20_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_0_LC_19_20_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_0_LC_19_20_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48293),
            .lcout(\I2C_top_level_inst1.s_addr0_o_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_1_LC_19_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_1_LC_19_20_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_1_LC_19_20_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_1_LC_19_20_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48158),
            .lcout(\I2C_top_level_inst1.s_addr0_o_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_2_LC_19_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_2_LC_19_20_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_2_LC_19_20_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_2_LC_19_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48107),
            .lcout(\I2C_top_level_inst1.s_addr0_o_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_3_LC_19_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_3_LC_19_20_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_3_LC_19_20_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_3_LC_19_20_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48049),
            .lcout(\I2C_top_level_inst1.s_addr0_o_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_4_LC_19_20_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_4_LC_19_20_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_4_LC_19_20_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_4_LC_19_20_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41379),
            .lcout(\I2C_top_level_inst1.s_addr0_o_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_5_LC_19_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_5_LC_19_20_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_5_LC_19_20_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_5_LC_19_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41808),
            .lcout(\I2C_top_level_inst1.s_addr0_o_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_6_LC_19_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_6_LC_19_20_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_6_LC_19_20_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_6_LC_19_20_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41753),
            .lcout(\I2C_top_level_inst1.s_addr0_o_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_7_LC_19_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_7_LC_19_20_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.addr0_reg_inst.c_addr0_7_LC_19_20_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.addr0_reg_inst.c_addr0_7_LC_19_20_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41691),
            .lcout(\I2C_top_level_inst1.s_addr0_o_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47992),
            .ce(N__43739),
            .sr(N__62853));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_0_LC_19_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_0_LC_19_21_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_0_LC_19_21_0 .LUT_INIT=16'b0011000111110101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_0_LC_19_21_0  (
            .in0(N__44142),
            .in1(N__47055),
            .in2(N__48330),
            .in3(N__41619),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_304_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_2_LC_19_21_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_2_LC_19_21_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_2_LC_19_21_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_2_LC_19_21_2  (
            .in0(N__66769),
            .in1(N__56661),
            .in2(N__41598),
            .in3(N__56818),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_0_LC_19_21_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_0_LC_19_21_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_0_LC_19_21_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_0_LC_19_21_3  (
            .in0(N__64374),
            .in1(N__56376),
            .in2(N__41583),
            .in3(N__41541),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNOZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_LC_19_21_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_LC_19_21_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_LC_19_21_4 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_LC_19_21_4  (
            .in0(N__56181),
            .in1(N__41563),
            .in2(N__41580),
            .in3(N__56594),
            .lcout(\I2C_top_level_inst1.s_no_restart ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65676),
            .ce(),
            .sr(N__65007));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_1_LC_19_21_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_1_LC_19_21_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_1_LC_19_21_5 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_1_LC_19_21_5  (
            .in0(N__64794),
            .in1(N__48325),
            .in2(N__44151),
            .in3(N__44141),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_LC_19_22_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_LC_19_22_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_LC_19_22_4 .LUT_INIT=16'b0010000011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_LC_19_22_4  (
            .in0(N__66867),
            .in1(N__64803),
            .in2(N__41517),
            .in3(N__41535),
            .lcout(\I2C_top_level_inst1.s_ack ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65685),
            .ce(),
            .sr(N__65011));
    defparam \serializer_mod_inst.shift_reg_6_LC_19_23_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_6_LC_19_23_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_6_LC_19_23_1 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_6_LC_19_23_1  (
            .in0(N__45461),
            .in1(N__41838),
            .in2(_gnd_net_),
            .in3(N__45040),
            .lcout(\serializer_mod_inst.shift_regZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65700),
            .ce(),
            .sr(N__62836));
    defparam \serializer_mod_inst.shift_reg_64_LC_19_23_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_64_LC_19_23_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_64_LC_19_23_4 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_64_LC_19_23_4  (
            .in0(N__45039),
            .in1(N__44199),
            .in2(_gnd_net_),
            .in3(N__45460),
            .lcout(\serializer_mod_inst.shift_regZ0Z_64 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65700),
            .ce(),
            .sr(N__62836));
    defparam \serializer_mod_inst.shift_reg_5_LC_19_24_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_5_LC_19_24_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_5_LC_19_24_0 .LUT_INIT=16'b0010001011001100;
    LogicCell40 \serializer_mod_inst.shift_reg_5_LC_19_24_0  (
            .in0(N__41820),
            .in1(N__45045),
            .in2(_gnd_net_),
            .in3(N__45456),
            .lcout(\serializer_mod_inst.shift_regZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65718),
            .ce(),
            .sr(N__62833));
    defparam \serializer_mod_inst.shift_reg_3_LC_19_24_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_3_LC_19_24_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_3_LC_19_24_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_3_LC_19_24_1  (
            .in0(N__47730),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41832),
            .lcout(\serializer_mod_inst.shift_regZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65718),
            .ce(),
            .sr(N__62833));
    defparam \serializer_mod_inst.shift_reg_4_LC_19_24_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_4_LC_19_24_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_4_LC_19_24_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_4_LC_19_24_4  (
            .in0(_gnd_net_),
            .in1(N__41826),
            .in2(_gnd_net_),
            .in3(N__47731),
            .lcout(\serializer_mod_inst.shift_regZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65718),
            .ce(),
            .sr(N__62833));
    defparam \serializer_mod_inst.shift_reg_28_LC_19_24_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_28_LC_19_24_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_28_LC_19_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_28_LC_19_24_5  (
            .in0(N__47729),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41949),
            .lcout(\serializer_mod_inst.shift_regZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65718),
            .ce(),
            .sr(N__62833));
    defparam \serializer_mod_inst.shift_reg_126_LC_19_24_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_126_LC_19_24_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_126_LC_19_24_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_126_LC_19_24_6  (
            .in0(_gnd_net_),
            .in1(N__41886),
            .in2(_gnd_net_),
            .in3(N__47728),
            .lcout(\serializer_mod_inst.shift_regZ0Z_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65718),
            .ce(),
            .sr(N__62833));
    defparam \serializer_mod_inst.shift_reg_24_LC_19_25_1 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_24_LC_19_25_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_24_LC_19_25_1 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_24_LC_19_25_1  (
            .in0(N__45454),
            .in1(N__41937),
            .in2(_gnd_net_),
            .in3(N__45043),
            .lcout(\serializer_mod_inst.shift_regZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65727),
            .ce(),
            .sr(N__62826));
    defparam \serializer_mod_inst.shift_reg_21_LC_19_25_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_21_LC_19_25_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_21_LC_19_25_2 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_21_LC_19_25_2  (
            .in0(N__45041),
            .in1(N__41904),
            .in2(_gnd_net_),
            .in3(N__45452),
            .lcout(\serializer_mod_inst.shift_regZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65727),
            .ce(),
            .sr(N__62826));
    defparam \serializer_mod_inst.shift_reg_27_LC_19_25_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_27_LC_19_25_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_27_LC_19_25_3 .LUT_INIT=16'b0101010110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_27_LC_19_25_3  (
            .in0(N__45455),
            .in1(N__41853),
            .in2(_gnd_net_),
            .in3(N__45044),
            .lcout(\serializer_mod_inst.shift_regZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65727),
            .ce(),
            .sr(N__62826));
    defparam \serializer_mod_inst.shift_reg_23_LC_19_25_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_23_LC_19_25_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_23_LC_19_25_4 .LUT_INIT=16'b0100010010101010;
    LogicCell40 \serializer_mod_inst.shift_reg_23_LC_19_25_4  (
            .in0(N__45042),
            .in1(N__41943),
            .in2(_gnd_net_),
            .in3(N__45453),
            .lcout(\serializer_mod_inst.shift_regZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65727),
            .ce(),
            .sr(N__62826));
    defparam \serializer_mod_inst.shift_reg_109_LC_19_25_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_109_LC_19_25_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_109_LC_19_25_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_109_LC_19_25_5  (
            .in0(_gnd_net_),
            .in1(N__41931),
            .in2(_gnd_net_),
            .in3(N__47706),
            .lcout(\serializer_mod_inst.shift_regZ0Z_109 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65727),
            .ce(),
            .sr(N__62826));
    defparam \serializer_mod_inst.shift_reg_20_LC_19_25_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_20_LC_19_25_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_20_LC_19_25_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_20_LC_19_25_6  (
            .in0(N__47707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41913),
            .lcout(\serializer_mod_inst.shift_regZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65727),
            .ce(),
            .sr(N__62826));
    defparam \serializer_mod_inst.shift_reg_124_LC_19_26_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_124_LC_19_26_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_124_LC_19_26_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_124_LC_19_26_0  (
            .in0(_gnd_net_),
            .in1(N__41865),
            .in2(_gnd_net_),
            .in3(N__47646),
            .lcout(\serializer_mod_inst.shift_regZ0Z_124 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65737),
            .ce(),
            .sr(N__62821));
    defparam \serializer_mod_inst.shift_reg_25_LC_19_26_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_25_LC_19_26_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_25_LC_19_26_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_25_LC_19_26_4  (
            .in0(_gnd_net_),
            .in1(N__41898),
            .in2(_gnd_net_),
            .in3(N__47648),
            .lcout(\serializer_mod_inst.shift_regZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65737),
            .ce(),
            .sr(N__62821));
    defparam \serializer_mod_inst.shift_reg_125_LC_19_26_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_125_LC_19_26_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_125_LC_19_26_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_125_LC_19_26_5  (
            .in0(N__47647),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41892),
            .lcout(\serializer_mod_inst.shift_regZ0Z_125 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65737),
            .ce(),
            .sr(N__62821));
    defparam \serializer_mod_inst.shift_reg_123_LC_19_26_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_123_LC_19_26_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_123_LC_19_26_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_123_LC_19_26_6  (
            .in0(_gnd_net_),
            .in1(N__41877),
            .in2(_gnd_net_),
            .in3(N__47645),
            .lcout(\serializer_mod_inst.shift_regZ0Z_123 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65737),
            .ce(),
            .sr(N__62821));
    defparam \serializer_mod_inst.shift_reg_26_LC_19_26_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_26_LC_19_26_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_26_LC_19_26_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_26_LC_19_26_7  (
            .in0(N__47649),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__41859),
            .lcout(\serializer_mod_inst.shift_regZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65737),
            .ce(),
            .sr(N__62821));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_27_LC_20_8_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_27_LC_20_8_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_27_LC_20_8_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_27_LC_20_8_1  (
            .in0(N__42144),
            .in1(N__52771),
            .in2(N__42126),
            .in3(N__52526),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_27_LC_20_8_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_27_LC_20_8_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_27_LC_20_8_2 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_27_LC_20_8_2  (
            .in0(N__49143),
            .in1(_gnd_net_),
            .in2(N__42105),
            .in3(N__52231),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_27_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_27_LC_20_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_27_LC_20_8_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_27_LC_20_8_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_27_LC_20_8_3  (
            .in0(N__42102),
            .in1(N__42096),
            .in2(N__42084),
            .in3(N__42060),
            .lcout(I2C_top_level_inst1_s_data_oreg_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65534),
            .ce(N__54500),
            .sr(N__65023));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_27_LC_20_8_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_27_LC_20_8_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_27_LC_20_8_4 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_27_LC_20_8_4  (
            .in0(N__51921),
            .in1(N__42081),
            .in2(N__48504),
            .in3(N__42072),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_16_LC_20_9_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_16_LC_20_9_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_16_LC_20_9_7 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_16_LC_20_9_7  (
            .in0(N__52998),
            .in1(N__53524),
            .in2(N__53323),
            .in3(N__54207),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_16_LC_20_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_16_LC_20_10_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_16_LC_20_10_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_16_LC_20_10_0  (
            .in0(N__42054),
            .in1(N__52745),
            .in2(N__42036),
            .in3(N__52492),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_16_LC_20_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_16_LC_20_10_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_16_LC_20_10_1 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_16_LC_20_10_1  (
            .in0(_gnd_net_),
            .in1(N__52187),
            .in2(N__42015),
            .in3(N__42012),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_16_LC_20_10_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_16_LC_20_10_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_16_LC_20_10_2 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_16_LC_20_10_2  (
            .in0(N__44432),
            .in1(N__41988),
            .in2(N__63134),
            .in3(N__44658),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_16_LC_20_10_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_16_LC_20_10_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_16_LC_20_10_3 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_16_LC_20_10_3  (
            .in0(N__41970),
            .in1(N__51922),
            .in2(N__41952),
            .in3(N__51657),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_16_LC_20_10_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_16_LC_20_10_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_16_LC_20_10_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_16_LC_20_10_4  (
            .in0(N__42336),
            .in1(N__42327),
            .in2(N__42321),
            .in3(N__42318),
            .lcout(I2C_top_level_inst1_s_data_oreg_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65554),
            .ce(N__54497),
            .sr(N__65018));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_24_LC_20_10_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_24_LC_20_10_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_24_LC_20_10_5 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_24_LC_20_10_5  (
            .in0(N__42312),
            .in1(N__44657),
            .in2(N__57608),
            .in3(N__44431),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_22_LC_20_11_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_22_LC_20_11_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_22_LC_20_11_0 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_22_LC_20_11_0  (
            .in0(N__59587),
            .in1(N__61348),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_3_LC_20_11_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_3_LC_20_11_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_3_LC_20_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_3_LC_20_11_1  (
            .in0(_gnd_net_),
            .in1(N__59589),
            .in2(_gnd_net_),
            .in3(N__63940),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_4_LC_20_11_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_4_LC_20_11_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_4_LC_20_11_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_4_LC_20_11_2  (
            .in0(_gnd_net_),
            .in1(N__59727),
            .in2(_gnd_net_),
            .in3(N__63827),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_5_LC_20_11_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_5_LC_20_11_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_5_LC_20_11_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_5_LC_20_11_3  (
            .in0(_gnd_net_),
            .in1(N__59590),
            .in2(_gnd_net_),
            .in3(N__63687),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_6_LC_20_11_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_6_LC_20_11_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_6_LC_20_11_4 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_6_LC_20_11_4  (
            .in0(N__59588),
            .in1(N__63581),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_7_LC_20_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_7_LC_20_11_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_7_LC_20_11_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_7_LC_20_11_5  (
            .in0(_gnd_net_),
            .in1(N__59591),
            .in2(_gnd_net_),
            .in3(N__63483),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_17_LC_20_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_17_LC_20_11_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_17_LC_20_11_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_17_LC_20_11_6  (
            .in0(_gnd_net_),
            .in1(N__59726),
            .in2(_gnd_net_),
            .in3(N__57392),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_9_LC_20_11_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_9_LC_20_11_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_9_LC_20_11_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_9_LC_20_11_7  (
            .in0(_gnd_net_),
            .in1(N__59592),
            .in2(_gnd_net_),
            .in3(N__46500),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65566),
            .ce(N__58880),
            .sr(N__62934));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQQQI1_LC_20_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQQQI1_LC_20_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQQQI1_LC_20_12_0 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQQQI1_LC_20_12_0  (
            .in0(N__46597),
            .in1(N__55249),
            .in2(N__42608),
            .in3(N__55449),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNID06H2_LC_20_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNID06H2_LC_20_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNID06H2_LC_20_12_1 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNID06H2_LC_20_12_1  (
            .in0(N__55056),
            .in1(N__46598),
            .in2(N__54835),
            .in3(N__42604),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8D7_LC_20_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8D7_LC_20_12_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8D7_LC_20_12_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8D7_LC_20_12_2  (
            .in0(N__53993),
            .in1(N__53371),
            .in2(N__42387),
            .in3(N__45546),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1RPF7_LC_20_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1RPF7_LC_20_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1RPF7_LC_20_12_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1RPF7_LC_20_12_3  (
            .in0(_gnd_net_),
            .in1(N__53714),
            .in2(N__42384),
            .in3(N__42381),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15_LC_20_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15_LC_20_12_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15_LC_20_12_4 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15_LC_20_12_4  (
            .in0(N__42375),
            .in1(_gnd_net_),
            .in2(N__42369),
            .in3(N__55724),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net ),
            .ce(N__55570),
            .sr(N__62925));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8D7_LC_20_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8D7_LC_20_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8D7_LC_20_12_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8D7_LC_20_12_5  (
            .in0(N__53960),
            .in1(N__54206),
            .in2(N__42366),
            .in3(N__45540),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI60QF7_LC_20_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI60QF7_LC_20_12_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI60QF7_LC_20_12_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI60QF7_LC_20_12_6  (
            .in0(N__53715),
            .in1(_gnd_net_),
            .in2(N__42357),
            .in3(N__42354),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_16_LC_20_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_16_LC_20_12_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_16_LC_20_12_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_16_LC_20_12_7  (
            .in0(N__55725),
            .in1(_gnd_net_),
            .in2(N__42348),
            .in3(N__42345),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net ),
            .ce(N__55570),
            .sr(N__62925));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_1_LC_20_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_1_LC_20_13_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_1_LC_20_13_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_1_LC_20_13_0  (
            .in0(N__59514),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61860),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_2_LC_20_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_2_LC_20_13_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_2_LC_20_13_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_2_LC_20_13_1  (
            .in0(_gnd_net_),
            .in1(N__61745),
            .in2(_gnd_net_),
            .in3(N__59511),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_3_LC_20_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_3_LC_20_13_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_3_LC_20_13_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_3_LC_20_13_2  (
            .in0(N__59515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__63945),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_4_LC_20_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_4_LC_20_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_4_LC_20_13_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_4_LC_20_13_3  (
            .in0(N__63789),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59512),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_9_LC_20_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_9_LC_20_13_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_9_LC_20_13_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_9_LC_20_13_4  (
            .in0(N__59516),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__46530),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_10_LC_20_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_10_LC_20_13_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_10_LC_20_13_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_10_LC_20_13_5  (
            .in0(_gnd_net_),
            .in1(N__58796),
            .in2(_gnd_net_),
            .in3(N__59509),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_11_LC_20_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_11_LC_20_13_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_11_LC_20_13_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_11_LC_20_13_6  (
            .in0(N__59513),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58691),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_20_LC_20_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_20_LC_20_13_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_20_LC_20_13_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_20_LC_20_13_7  (
            .in0(_gnd_net_),
            .in1(N__59510),
            .in2(_gnd_net_),
            .in3(N__61546),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65589),
            .ce(N__48724),
            .sr(N__62917));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_20_LC_20_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_20_LC_20_14_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_20_LC_20_14_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_20_LC_20_14_0  (
            .in0(N__59428),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61547),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_12_LC_20_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_12_LC_20_14_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_12_LC_20_14_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_12_LC_20_14_1  (
            .in0(N__58590),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59430),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_21_LC_20_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_21_LC_20_14_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_21_LC_20_14_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_21_LC_20_14_2  (
            .in0(N__59429),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61437),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_22_LC_20_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_22_LC_20_14_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_22_LC_20_14_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_22_LC_20_14_3  (
            .in0(_gnd_net_),
            .in1(N__61356),
            .in2(_gnd_net_),
            .in3(N__59424),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_14_LC_20_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_14_LC_20_14_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_14_LC_20_14_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_14_LC_20_14_4  (
            .in0(N__59426),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58499),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_23_LC_20_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_23_LC_20_14_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_23_LC_20_14_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_23_LC_20_14_5  (
            .in0(_gnd_net_),
            .in1(N__61248),
            .in2(_gnd_net_),
            .in3(N__59425),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_15_LC_20_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_15_LC_20_14_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_15_LC_20_14_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_15_LC_20_14_6  (
            .in0(N__59427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57535),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_16_LC_20_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_16_LC_20_14_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_16_LC_20_14_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_16_LC_20_14_7  (
            .in0(_gnd_net_),
            .in1(N__57618),
            .in2(_gnd_net_),
            .in3(N__59423),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65601),
            .ce(N__45571),
            .sr(N__62909));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISMV43_LC_20_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISMV43_LC_20_15_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISMV43_LC_20_15_0 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISMV43_LC_20_15_0  (
            .in0(N__46064),
            .in1(N__46369),
            .in2(N__45921),
            .in3(N__42550),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238D7_LC_20_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238D7_LC_20_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238D7_LC_20_15_1 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238D7_LC_20_15_1  (
            .in0(N__42514),
            .in1(N__54003),
            .in2(N__42489),
            .in3(N__42825),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID6PF7_LC_20_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID6PF7_LC_20_15_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID6PF7_LC_20_15_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID6PF7_LC_20_15_2  (
            .in0(N__46115),
            .in1(_gnd_net_),
            .in2(N__42828),
            .in3(N__53673),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5O5H2_LC_20_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5O5H2_LC_20_15_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5O5H2_LC_20_15_3 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5O5H2_LC_20_15_3  (
            .in0(N__54781),
            .in1(N__42940),
            .in2(N__55052),
            .in3(N__42905),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_11_LC_20_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_11_LC_20_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_11_LC_20_15_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_11_LC_20_15_4  (
            .in0(N__58701),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59431),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65609),
            .ce(N__45569),
            .sr(N__62899));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9S5H2_LC_20_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9S5H2_LC_20_15_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9S5H2_LC_20_15_5 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9S5H2_LC_20_15_5  (
            .in0(N__55022),
            .in1(N__54782),
            .in2(N__46159),
            .in3(N__42793),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_13_LC_20_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_13_LC_20_15_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_13_LC_20_15_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_13_LC_20_15_6  (
            .in0(_gnd_net_),
            .in1(N__58376),
            .in2(_gnd_net_),
            .in3(N__59432),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65609),
            .ce(N__45569),
            .sr(N__62899));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIB08H2_LC_20_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIB08H2_LC_20_15_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIB08H2_LC_20_15_7 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIB08H2_LC_20_15_7  (
            .in0(N__54780),
            .in1(N__49480),
            .in2(N__55053),
            .in3(N__49453),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIGGQI1_LC_20_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIGGQI1_LC_20_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIGGQI1_LC_20_16_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIGGQI1_LC_20_16_0  (
            .in0(N__55231),
            .in1(N__55427),
            .in2(N__42728),
            .in3(N__42751),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3M5H2_LC_20_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3M5H2_LC_20_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3M5H2_LC_20_16_1 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3M5H2_LC_20_16_1  (
            .in0(N__42724),
            .in1(N__55020),
            .in2(N__42758),
            .in3(N__54818),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_10_LC_20_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_10_LC_20_16_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_10_LC_20_16_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_10_LC_20_16_2  (
            .in0(N__59422),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58797),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65622),
            .ce(N__49063),
            .sr(N__62888));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNII6FN1_LC_20_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNII6FN1_LC_20_16_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNII6FN1_LC_20_16_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNII6FN1_LC_20_16_3  (
            .in0(N__55429),
            .in1(N__55232),
            .in2(N__43004),
            .in3(N__42964),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_2_LC_20_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_2_LC_20_16_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_2_LC_20_16_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_2_LC_20_16_4  (
            .in0(N__59421),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61719),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65622),
            .ce(N__49063),
            .sr(N__62888));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5CQL2_LC_20_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5CQL2_LC_20_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5CQL2_LC_20_16_5 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5CQL2_LC_20_16_5  (
            .in0(N__55021),
            .in1(N__54817),
            .in2(N__43003),
            .in3(N__42965),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIIQI1_LC_20_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIIQI1_LC_20_16_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIIQI1_LC_20_16_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIIQI1_LC_20_16_6  (
            .in0(N__55230),
            .in1(N__55428),
            .in2(N__42944),
            .in3(N__42904),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_11_LC_20_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_11_LC_20_16_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_11_LC_20_16_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_11_LC_20_16_7  (
            .in0(_gnd_net_),
            .in1(N__59420),
            .in2(_gnd_net_),
            .in3(N__58700),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65622),
            .ce(N__49063),
            .sr(N__62888));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_c_0_LC_20_17_0 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_c_0_LC_20_17_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_c_0_LC_20_17_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_c_0_LC_20_17_0  (
            .in0(_gnd_net_),
            .in1(N__55982),
            .in2(N__46763),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_20_17_0_),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_1_LC_20_17_1 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_1_LC_20_17_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_1_LC_20_17_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_1_LC_20_17_1  (
            .in0(_gnd_net_),
            .in1(N__46824),
            .in2(_gnd_net_),
            .in3(N__42873),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_1 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_2_LC_20_17_2 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_2_LC_20_17_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_2_LC_20_17_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_2_LC_20_17_2  (
            .in0(_gnd_net_),
            .in1(N__46907),
            .in2(_gnd_net_),
            .in3(N__42855),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_2 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_LUT4_0_LC_20_17_3 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_LUT4_0_LC_20_17_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_LUT4_0_LC_20_17_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_LUT4_0_LC_20_17_3  (
            .in0(_gnd_net_),
            .in1(N__54338),
            .in2(_gnd_net_),
            .in3(N__42840),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_4_LC_20_17_4 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_4_LC_20_17_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_4_LC_20_17_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_4_LC_20_17_4  (
            .in0(_gnd_net_),
            .in1(N__47197),
            .in2(_gnd_net_),
            .in3(N__42831),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_4 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_5_LC_20_17_5 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_5_LC_20_17_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_5_LC_20_17_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_5_LC_20_17_5  (
            .in0(_gnd_net_),
            .in1(N__47247),
            .in2(_gnd_net_),
            .in3(N__43104),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_5 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_6_LC_20_17_6 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_6_LC_20_17_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_6_LC_20_17_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_6_LC_20_17_6  (
            .in0(_gnd_net_),
            .in1(N__47170),
            .in2(_gnd_net_),
            .in3(N__43089),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_6 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_7_LC_20_17_7 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_7_LC_20_17_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_7_LC_20_17_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_7_LC_20_17_7  (
            .in0(_gnd_net_),
            .in1(N__47118),
            .in2(_gnd_net_),
            .in3(N__43074),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_7 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_LUT4_0_LC_20_18_0 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_LUT4_0_LC_20_18_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_LUT4_0_LC_20_18_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_LUT4_0_LC_20_18_0  (
            .in0(_gnd_net_),
            .in1(N__56122),
            .in2(_gnd_net_),
            .in3(N__43071),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_20_18_0_),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_9_LC_20_18_1 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_9_LC_20_18_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_9_LC_20_18_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_9_LC_20_18_1  (
            .in0(_gnd_net_),
            .in1(N__47008),
            .in2(_gnd_net_),
            .in3(N__43062),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_9 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_10_LC_20_18_2 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_10_LC_20_18_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_10_LC_20_18_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_10_LC_20_18_2  (
            .in0(_gnd_net_),
            .in1(N__47037),
            .in2(_gnd_net_),
            .in3(N__43053),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_10 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_11_LC_20_18_3 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_11_LC_20_18_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_11_LC_20_18_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_11_LC_20_18_3  (
            .in0(_gnd_net_),
            .in1(N__46942),
            .in2(_gnd_net_),
            .in3(N__43044),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_11 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_12_LC_20_18_4 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_12_LC_20_18_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_12_LC_20_18_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_12_LC_20_18_4  (
            .in0(_gnd_net_),
            .in1(N__43041),
            .in2(_gnd_net_),
            .in3(N__43008),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_12 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_13_LC_20_18_5 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_13_LC_20_18_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_13_LC_20_18_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_13_LC_20_18_5  (
            .in0(_gnd_net_),
            .in1(N__43275),
            .in2(_gnd_net_),
            .in3(N__43245),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_13 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_14_LC_20_18_6 .C_ON=1'b1;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_14_LC_20_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_14_LC_20_18_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_14_LC_20_18_6  (
            .in0(_gnd_net_),
            .in1(N__43242),
            .in2(_gnd_net_),
            .in3(N__43212),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_14 ),
            .ltout(),
            .carryin(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13 ),
            .carryout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_15_LC_20_18_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_15_LC_20_18_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_15_LC_20_18_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_15_LC_20_18_7  (
            .in0(_gnd_net_),
            .in1(N__43209),
            .in2(_gnd_net_),
            .in3(N__43188),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_13_LC_20_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_13_LC_20_19_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_13_LC_20_19_0 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_13_LC_20_19_0  (
            .in0(N__56621),
            .in1(N__66264),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_103_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_2_LC_20_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_2_LC_20_19_1 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_2_LC_20_19_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_2_LC_20_19_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43158),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65661),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_1_LC_20_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_1_LC_20_19_2 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_1_LC_20_19_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_1_LC_20_19_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43152),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65661),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_0_LC_20_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_0_LC_20_19_3 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_0_LC_20_19_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_0_LC_20_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43746),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65661),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIABID_21_LC_20_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIABID_21_LC_20_19_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIABID_21_LC_20_19_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIABID_21_LC_20_19_4  (
            .in0(N__56232),
            .in1(N__43619),
            .in2(_gnd_net_),
            .in3(N__43146),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_291 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_291_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_0_LC_20_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_0_LC_20_19_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_0_LC_20_19_5 .LUT_INIT=16'b0100000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_0_LC_20_19_5  (
            .in0(N__66794),
            .in1(N__56620),
            .in2(N__43119),
            .in3(N__57237),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_RNO_0_LC_20_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_RNO_0_LC_20_19_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_RNO_0_LC_20_19_6 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_RNO_0_LC_20_19_6  (
            .in0(N__43747),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43669),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_6_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_0_LC_20_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_0_LC_20_19_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_0_LC_20_19_7 .LUT_INIT=16'b1000100011011101;
    LogicCell40 \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_0_LC_20_19_7  (
            .in0(N__43670),
            .in1(N__50886),
            .in2(_gnd_net_),
            .in3(N__43836),
            .lcout(\I2C_top_level_inst1.I2C_FSM_inst.N_1378 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI5MGJ_2_LC_20_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI5MGJ_2_LC_20_20_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI5MGJ_2_LC_20_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI5MGJ_2_LC_20_20_0  (
            .in0(N__65871),
            .in1(N__56361),
            .in2(N__64789),
            .in3(N__56816),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m24_i_a3_LC_20_20_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m24_i_a3_LC_20_20_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m24_i_a3_LC_20_20_1 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m24_i_a3_LC_20_20_1  (
            .in0(N__56817),
            .in1(N__66273),
            .in2(N__65986),
            .in3(N__65872),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_1676_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_2_LC_20_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_2_LC_20_20_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_2_LC_20_20_2 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_2_LC_20_20_2  (
            .in0(N__66165),
            .in1(N__64343),
            .in2(N__43626),
            .in3(N__62455),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65677),
            .ce(),
            .sr(N__65008));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_22_LC_20_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_22_LC_20_20_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_22_LC_20_20_3 .LUT_INIT=16'b0010001000100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_22_LC_20_20_3  (
            .in0(N__43623),
            .in1(N__66164),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65677),
            .ce(),
            .sr(N__65008));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIEVJ7_22_LC_20_20_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIEVJ7_22_LC_20_20_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIEVJ7_22_LC_20_20_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIEVJ7_22_LC_20_20_4  (
            .in0(_gnd_net_),
            .in1(N__65974),
            .in2(_gnd_net_),
            .in3(N__56815),
            .lcout(c_state_RNIEVJ7_22),
            .ltout(c_state_RNIEVJ7_22_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASSA_22_LC_20_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASSA_22_LC_20_20_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASSA_22_LC_20_20_5 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASSA_22_LC_20_20_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__43587),
            .in3(N__43513),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_77_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_14_LC_20_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_14_LC_20_20_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_14_LC_20_20_6 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_14_LC_20_20_6  (
            .in0(N__57123),
            .in1(N__57089),
            .in2(N__43299),
            .in3(N__64432),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_0_LC_20_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_0_LC_20_21_0 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_0_LC_20_21_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_0_LC_20_21_0  (
            .in0(N__43955),
            .in1(N__43905),
            .in2(_gnd_net_),
            .in3(N__48290),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65686),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_2_1_4_LC_20_21_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_2_1_4_LC_20_21_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_2_1_4_LC_20_21_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_2_1_4_LC_20_21_1  (
            .in0(_gnd_net_),
            .in1(N__48195),
            .in2(_gnd_net_),
            .in3(N__50112),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1606_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_2_LC_20_21_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_2_LC_20_21_2 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_2_LC_20_21_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_2_LC_20_21_2  (
            .in0(N__43767),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65686),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_0_LC_20_21_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_0_LC_20_21_3 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_0_LC_20_21_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_0_LC_20_21_3  (
            .in0(N__43857),
            .in1(N__43829),
            .in2(_gnd_net_),
            .in3(N__43794),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65686),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_2_LC_20_21_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_2_LC_20_21_4 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_2_LC_20_21_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_2_LC_20_21_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43755),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65686),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_1_LC_20_21_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_1_LC_20_21_5 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_1_LC_20_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_1_LC_20_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43773),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65686),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_15_LC_20_21_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_15_LC_20_21_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_15_LC_20_21_6 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_15_LC_20_21_6  (
            .in0(N__66150),
            .in1(N__48310),
            .in2(_gnd_net_),
            .in3(N__44140),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_607 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_1_LC_20_21_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_1_LC_20_21_7 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_1_LC_20_21_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_1_LC_20_21_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43761),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65686),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI1I79_18_LC_20_22_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI1I79_18_LC_20_22_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI1I79_18_LC_20_22_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI1I79_18_LC_20_22_2  (
            .in0(N__47563),
            .in1(N__50536),
            .in2(_gnd_net_),
            .in3(N__56584),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_294 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_4_LC_20_22_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_4_LC_20_22_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_4_LC_20_22_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_4_LC_20_22_3  (
            .in0(_gnd_net_),
            .in1(N__47562),
            .in2(_gnd_net_),
            .in3(N__56729),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_0_1_LC_20_22_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_0_1_LC_20_22_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_0_1_LC_20_22_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_0_1_LC_20_22_4  (
            .in0(_gnd_net_),
            .in1(N__56583),
            .in2(_gnd_net_),
            .in3(N__50113),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_RNISHA8_2_LC_20_22_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_RNISHA8_2_LC_20_22_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_RNISHA8_2_LC_20_22_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_RNISHA8_2_LC_20_22_5  (
            .in0(N__50537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50933),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_0_LC_20_22_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_0_LC_20_22_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_0_LC_20_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_0_LC_20_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48291),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65701),
            .ce(N__44061),
            .sr(N__65019));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_1_LC_20_22_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_1_LC_20_22_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_1_LC_20_22_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_1_LC_20_22_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48156),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65701),
            .ce(N__44061),
            .sr(N__65019));
    defparam \serializer_mod_inst.shift_reg_65_LC_20_23_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_65_LC_20_23_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_65_LC_20_23_3 .LUT_INIT=16'b0011001110001000;
    LogicCell40 \serializer_mod_inst.shift_reg_65_LC_20_23_3  (
            .in0(N__44025),
            .in1(N__45446),
            .in2(_gnd_net_),
            .in3(N__45046),
            .lcout(\serializer_mod_inst.shift_regZ0Z_65 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65719),
            .ce(),
            .sr(N__62842));
    defparam \serializer_mod_inst.shift_reg_128_LC_20_23_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_128_LC_20_23_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_128_LC_20_23_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_128_LC_20_23_4  (
            .in0(N__47814),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__43968),
            .lcout(\serializer_mod_inst.shift_regZ0Z_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65719),
            .ce(),
            .sr(N__62842));
    defparam \serializer_mod_inst.shift_reg_127_LC_20_23_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_127_LC_20_23_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_127_LC_20_23_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_127_LC_20_23_5  (
            .in0(_gnd_net_),
            .in1(N__43974),
            .in2(_gnd_net_),
            .in3(N__47813),
            .lcout(\serializer_mod_inst.shift_regZ0Z_127 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65719),
            .ce(),
            .sr(N__62842));
    defparam \serializer_mod_inst.shift_reg_29_LC_20_24_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_29_LC_20_24_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_29_LC_20_24_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_29_LC_20_24_2  (
            .in0(_gnd_net_),
            .in1(N__43962),
            .in2(_gnd_net_),
            .in3(N__47724),
            .lcout(\serializer_mod_inst.shift_regZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65728),
            .ce(),
            .sr(N__62837));
    defparam \serializer_mod_inst.shift_reg_62_LC_20_24_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_62_LC_20_24_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_62_LC_20_24_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_62_LC_20_24_3  (
            .in0(N__47726),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44175),
            .lcout(\serializer_mod_inst.shift_regZ0Z_62 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65728),
            .ce(),
            .sr(N__62837));
    defparam \serializer_mod_inst.shift_reg_30_LC_20_24_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_30_LC_20_24_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_30_LC_20_24_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_30_LC_20_24_5  (
            .in0(N__47725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44220),
            .lcout(\serializer_mod_inst.shift_regZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65728),
            .ce(),
            .sr(N__62837));
    defparam \serializer_mod_inst.shift_reg_63_LC_20_24_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_63_LC_20_24_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_63_LC_20_24_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_63_LC_20_24_7  (
            .in0(N__47727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44205),
            .lcout(\serializer_mod_inst.shift_regZ0Z_63 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65728),
            .ce(),
            .sr(N__62837));
    defparam \serializer_mod_inst.shift_reg_58_LC_20_25_2 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_58_LC_20_25_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_58_LC_20_25_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_58_LC_20_25_2  (
            .in0(_gnd_net_),
            .in1(N__44157),
            .in2(_gnd_net_),
            .in3(N__47651),
            .lcout(\serializer_mod_inst.shift_regZ0Z_58 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65738),
            .ce(),
            .sr(N__62834));
    defparam \serializer_mod_inst.shift_reg_59_LC_20_25_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_59_LC_20_25_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_59_LC_20_25_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_59_LC_20_25_3  (
            .in0(N__47652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44193),
            .lcout(\serializer_mod_inst.shift_regZ0Z_59 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65738),
            .ce(),
            .sr(N__62834));
    defparam \serializer_mod_inst.shift_reg_60_LC_20_25_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_60_LC_20_25_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_60_LC_20_25_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_60_LC_20_25_4  (
            .in0(_gnd_net_),
            .in1(N__44187),
            .in2(_gnd_net_),
            .in3(N__47653),
            .lcout(\serializer_mod_inst.shift_regZ0Z_60 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65738),
            .ce(),
            .sr(N__62834));
    defparam \serializer_mod_inst.shift_reg_61_LC_20_25_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_61_LC_20_25_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_61_LC_20_25_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_61_LC_20_25_5  (
            .in0(N__47654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__44181),
            .lcout(\serializer_mod_inst.shift_regZ0Z_61 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65738),
            .ce(),
            .sr(N__62834));
    defparam \serializer_mod_inst.shift_reg_57_LC_20_25_6 .C_ON=1'b0;
    defparam \serializer_mod_inst.shift_reg_57_LC_20_25_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.shift_reg_57_LC_20_25_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \serializer_mod_inst.shift_reg_57_LC_20_25_6  (
            .in0(_gnd_net_),
            .in1(N__44169),
            .in2(_gnd_net_),
            .in3(N__47650),
            .lcout(\serializer_mod_inst.shift_regZ0Z_57 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65738),
            .ce(),
            .sr(N__62834));
    defparam \serializer_mod_inst.current_state_RNIVDDK_0_0_LC_20_26_0 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_RNIVDDK_0_0_LC_20_26_0 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.current_state_RNIVDDK_0_0_LC_20_26_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \serializer_mod_inst.current_state_RNIVDDK_0_0_LC_20_26_0  (
            .in0(N__45201),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__45035),
            .lcout(\serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.current_state_RNO_1_0_LC_20_26_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_RNO_1_0_LC_20_26_3 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.current_state_RNO_1_0_LC_20_26_3 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \serializer_mod_inst.current_state_RNO_1_0_LC_20_26_3  (
            .in0(_gnd_net_),
            .in1(N__48430),
            .in2(_gnd_net_),
            .in3(N__48478),
            .lcout(),
            .ltout(\serializer_mod_inst.un22_next_state_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.current_state_RNO_0_0_LC_20_26_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_RNO_0_0_LC_20_26_4 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.current_state_RNO_0_0_LC_20_26_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \serializer_mod_inst.current_state_RNO_0_0_LC_20_26_4  (
            .in0(N__48616),
            .in1(N__48458),
            .in2(N__45501),
            .in3(N__48489),
            .lcout(\serializer_mod_inst.un22_next_state ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.current_state_RNIVDDK_0_LC_20_27_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_RNIVDDK_0_LC_20_27_5 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.current_state_RNIVDDK_0_LC_20_27_5 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \serializer_mod_inst.current_state_RNIVDDK_0_LC_20_27_5  (
            .in0(_gnd_net_),
            .in1(N__45402),
            .in2(_gnd_net_),
            .in3(N__45088),
            .lcout(\serializer_mod_inst.next_state32_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_0_LC_21_7_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_0_LC_21_7_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_0_LC_21_7_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_0_LC_21_7_3  (
            .in0(N__44244),
            .in1(N__44250),
            .in2(N__44721),
            .in3(N__44706),
            .lcout(I2C_top_level_inst1_s_data_oreg_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65535),
            .ce(N__54501),
            .sr(N__65028));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_0_LC_21_8_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_0_LC_21_8_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_0_LC_21_8_0 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_0_LC_21_8_0  (
            .in0(N__44691),
            .in1(N__44676),
            .in2(N__44454),
            .in3(N__44433),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_0_LC_21_8_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_0_LC_21_8_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_0_LC_21_8_1 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_0_LC_21_8_1  (
            .in0(N__44274),
            .in1(N__51920),
            .in2(N__44253),
            .in3(N__58256),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_0_LC_21_8_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_0_LC_21_8_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_0_LC_21_8_3 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_0_LC_21_8_3  (
            .in0(N__58227),
            .in1(N__53014),
            .in2(N__53310),
            .in3(N__60645),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_25_LC_21_10_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_25_LC_21_10_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_25_LC_21_10_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_25_LC_21_10_0  (
            .in0(N__61018),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59717),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65567),
            .ce(N__45573),
            .sr(N__62946));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_17_LC_21_10_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_17_LC_21_10_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_17_LC_21_10_1 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_17_LC_21_10_1  (
            .in0(N__57412),
            .in1(_gnd_net_),
            .in2(N__59729),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65567),
            .ce(N__45573),
            .sr(N__62946));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_26_LC_21_10_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_26_LC_21_10_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_26_LC_21_10_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_26_LC_21_10_2  (
            .in0(_gnd_net_),
            .in1(N__59718),
            .in2(_gnd_net_),
            .in3(N__60905),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_3Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65567),
            .ce(N__45573),
            .sr(N__62946));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_18_LC_21_10_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_18_LC_21_10_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_18_LC_21_10_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_18_LC_21_10_3  (
            .in0(N__59844),
            .in1(_gnd_net_),
            .in2(N__59730),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65567),
            .ce(N__45573),
            .sr(N__62946));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_19_LC_21_10_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_19_LC_21_10_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_19_LC_21_10_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_19_LC_21_10_4  (
            .in0(_gnd_net_),
            .in1(N__59716),
            .in2(_gnd_net_),
            .in3(N__61644),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65567),
            .ce(N__45573),
            .sr(N__62946));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_0_LC_21_10_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_0_LC_21_10_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_0_LC_21_10_5 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_0_LC_21_10_5  (
            .in0(N__59719),
            .in1(N__61930),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkstopmask_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65567),
            .ce(N__45573),
            .sr(N__62946));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4VV43_LC_21_11_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4VV43_LC_21_11_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4VV43_LC_21_11_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4VV43_LC_21_11_0  (
            .in0(N__45903),
            .in1(N__46056),
            .in2(N__48565),
            .in3(N__46198),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI61053_LC_21_11_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI61053_LC_21_11_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI61053_LC_21_11_1 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI61053_LC_21_11_1  (
            .in0(N__46054),
            .in1(N__45904),
            .in2(N__53525),
            .in3(N__51652),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI6LK93_LC_21_11_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI6LK93_LC_21_11_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI6LK93_LC_21_11_2 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI6LK93_LC_21_11_2  (
            .in0(N__46057),
            .in1(N__45530),
            .in2(N__45919),
            .in3(N__48745),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIA5053_LC_21_11_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIA5053_LC_21_11_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIA5053_LC_21_11_3 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIA5053_LC_21_11_3  (
            .in0(N__46055),
            .in1(N__45905),
            .in2(N__51434),
            .in3(N__51364),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIAPK93_LC_21_11_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIAPK93_LC_21_11_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIAPK93_LC_21_11_4 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIAPK93_LC_21_11_4  (
            .in0(N__45906),
            .in1(N__46052),
            .in2(N__49382),
            .in3(N__49819),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIC7053_LC_21_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIC7053_LC_21_11_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIC7053_LC_21_11_5 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIC7053_LC_21_11_5  (
            .in0(N__46053),
            .in1(N__45907),
            .in2(N__51505),
            .in3(N__57323),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIO6K93_LC_21_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIO6K93_LC_21_11_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIO6K93_LC_21_11_6 .LUT_INIT=16'b1010001011110011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIO6K93_LC_21_11_6  (
            .in0(N__46058),
            .in1(N__60641),
            .in2(N__45920),
            .in3(N__58246),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQ8K93_LC_21_11_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQ8K93_LC_21_11_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQ8K93_LC_21_11_7 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQ8K93_LC_21_11_7  (
            .in0(N__46051),
            .in1(N__45908),
            .in2(N__60709),
            .in3(N__57826),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUUQI1_LC_21_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUUQI1_LC_21_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUUQI1_LC_21_12_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUUQI1_LC_21_12_0  (
            .in0(N__55262),
            .in1(N__55450),
            .in2(N__46556),
            .in3(N__45613),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI83053_LC_21_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI83053_LC_21_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI83053_LC_21_12_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI83053_LC_21_12_1  (
            .in0(N__45902),
            .in1(N__46059),
            .in2(N__51588),
            .in3(N__51610),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029D7_LC_21_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029D7_LC_21_12_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029D7_LC_21_12_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029D7_LC_21_12_2  (
            .in0(N__53961),
            .in1(N__54152),
            .in2(N__45645),
            .in3(N__45594),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB5QF7_LC_21_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB5QF7_LC_21_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB5QF7_LC_21_12_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB5QF7_LC_21_12_3  (
            .in0(_gnd_net_),
            .in1(N__53721),
            .in2(N__45642),
            .in3(N__45639),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17_LC_21_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17_LC_21_12_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17_LC_21_12_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17_LC_21_12_4  (
            .in0(N__55744),
            .in1(_gnd_net_),
            .in2(N__45633),
            .in3(N__45630),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net ),
            .ce(N__55558),
            .sr(N__62935));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIH46H2_LC_21_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIH46H2_LC_21_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIH46H2_LC_21_12_5 .LUT_INIT=16'b1010111100100011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIH46H2_LC_21_12_5  (
            .in0(N__54816),
            .in1(N__46552),
            .in2(N__45618),
            .in3(N__55055),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_0_LC_21_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_0_LC_21_12_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_0_LC_21_12_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_0_LC_21_12_6  (
            .in0(N__55742),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48878),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net ),
            .ce(N__55558),
            .sr(N__62935));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_11_LC_21_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_11_LC_21_12_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_11_LC_21_12_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_11_LC_21_12_7  (
            .in0(N__46686),
            .in1(N__55743),
            .in2(_gnd_net_),
            .in3(N__46116),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net ),
            .ce(N__55558),
            .sr(N__62935));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIS1692_17_LC_21_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIS1692_17_LC_21_13_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIS1692_17_LC_21_13_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIS1692_17_LC_21_13_0  (
            .in0(N__57981),
            .in1(N__58179),
            .in2(N__45743),
            .in3(N__45763),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LH5_LC_21_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LH5_LC_21_13_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LH5_LC_21_13_1 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LH5_LC_21_13_1  (
            .in0(N__60597),
            .in1(N__46306),
            .in2(N__46089),
            .in3(N__46074),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LHZ0Z5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKMSI1_LC_21_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKMSI1_LC_21_13_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKMSI1_LC_21_13_2 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKMSI1_LC_21_13_2  (
            .in0(N__55254),
            .in1(N__55444),
            .in2(N__45674),
            .in3(N__45691),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_21_LC_21_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_21_LC_21_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_21_LC_21_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_21_LC_21_13_3  (
            .in0(N__59508),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61435),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65602),
            .ce(N__49093),
            .sr(N__62926));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUQ153_LC_21_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUQ153_LC_21_13_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUQ153_LC_21_13_4 .LUT_INIT=16'b1100010011110101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUQ153_LC_21_13_4  (
            .in0(N__46307),
            .in1(N__46060),
            .in2(N__45870),
            .in3(N__45764),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_21_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDD7_LC_21_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDD7_LC_21_13_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDD7_LC_21_13_5 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDD7_LC_21_13_5  (
            .in0(N__45742),
            .in1(N__53966),
            .in2(N__45711),
            .in3(N__45651),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDDZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7S7H2_LC_21_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7S7H2_LC_21_13_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7S7H2_LC_21_13_6 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7S7H2_LC_21_13_6  (
            .in0(N__54806),
            .in1(N__45692),
            .in2(N__55019),
            .in3(N__45670),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_11_LC_21_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_11_LC_21_14_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_11_LC_21_14_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_11_LC_21_14_0  (
            .in0(_gnd_net_),
            .in1(N__58696),
            .in2(_gnd_net_),
            .in3(N__59416),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_12_LC_21_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_12_LC_21_14_1 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_12_LC_21_14_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_12_LC_21_14_1  (
            .in0(N__59412),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58591),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_21_LC_21_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_21_LC_21_14_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_21_LC_21_14_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_21_LC_21_14_2  (
            .in0(_gnd_net_),
            .in1(N__61434),
            .in2(_gnd_net_),
            .in3(N__59418),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_21),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_30_LC_21_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_30_LC_21_14_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_30_LC_21_14_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_30_LC_21_14_3  (
            .in0(N__59415),
            .in1(_gnd_net_),
            .in2(N__62183),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_13_LC_21_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_13_LC_21_14_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_13_LC_21_14_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_13_LC_21_14_4  (
            .in0(N__58364),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59417),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_25_LC_21_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_25_LC_21_14_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_25_LC_21_14_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_25_LC_21_14_5  (
            .in0(N__59414),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61019),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_31_LC_21_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_31_LC_21_14_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_31_LC_21_14_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_31_LC_21_14_6  (
            .in0(_gnd_net_),
            .in1(N__62072),
            .in2(_gnd_net_),
            .in3(N__59419),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_15_LC_21_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_15_LC_21_14_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_15_LC_21_14_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_15_LC_21_14_7  (
            .in0(N__59413),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57536),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65610),
            .ce(N__58868),
            .sr(N__62918));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_13_LC_21_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_13_LC_21_15_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_13_LC_21_15_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_13_LC_21_15_0  (
            .in0(N__59433),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58377),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_31_LC_21_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_31_LC_21_15_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_31_LC_21_15_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_31_LC_21_15_1  (
            .in0(_gnd_net_),
            .in1(N__59439),
            .in2(_gnd_net_),
            .in3(N__62073),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_23_LC_21_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_23_LC_21_15_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_23_LC_21_15_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_23_LC_21_15_2  (
            .in0(N__59435),
            .in1(N__61254),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_15_LC_21_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_15_LC_21_15_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_15_LC_21_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_15_LC_21_15_3  (
            .in0(_gnd_net_),
            .in1(N__59437),
            .in2(_gnd_net_),
            .in3(N__57540),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_24_LC_21_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_24_LC_21_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_24_LC_21_15_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_24_LC_21_15_4  (
            .in0(N__59436),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61117),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_25_LC_21_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_25_LC_21_15_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_25_LC_21_15_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_25_LC_21_15_5  (
            .in0(_gnd_net_),
            .in1(N__59438),
            .in2(_gnd_net_),
            .in3(N__61013),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_17_LC_21_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_17_LC_21_15_6 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_17_LC_21_15_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_17_LC_21_15_6  (
            .in0(N__59434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57414),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_9_LC_21_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_9_LC_21_15_7 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_9_LC_21_15_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_9_LC_21_15_7  (
            .in0(_gnd_net_),
            .in1(N__59440),
            .in2(_gnd_net_),
            .in3(N__46526),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65623),
            .ce(N__49071),
            .sr(N__62910));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSL7_LC_21_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSL7_LC_21_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSL7_LC_21_16_0 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSL7_LC_21_16_0  (
            .in0(N__53967),
            .in1(N__49427),
            .in2(N__46419),
            .in3(N__46614),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI0FDO7_LC_21_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI0FDO7_LC_21_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI0FDO7_LC_21_16_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI0FDO7_LC_21_16_1  (
            .in0(_gnd_net_),
            .in1(N__53674),
            .in2(N__46404),
            .in3(N__46401),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9_LC_21_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9_LC_21_16_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9_LC_21_16_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9_LC_21_16_2  (
            .in0(N__55727),
            .in1(_gnd_net_),
            .in2(N__46395),
            .in3(N__46392),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net ),
            .ce(N__55571),
            .sr(N__62900));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7D7_LC_21_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7D7_LC_21_16_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7D7_LC_21_16_3 .LUT_INIT=16'b0111010111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7D7_LC_21_16_3  (
            .in0(N__46725),
            .in1(N__53968),
            .in2(N__49344),
            .in3(N__46710),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI81PF7_LC_21_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI81PF7_LC_21_16_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI81PF7_LC_21_16_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI81PF7_LC_21_16_4  (
            .in0(N__53675),
            .in1(_gnd_net_),
            .in2(N__46704),
            .in3(N__46701),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_10_LC_21_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_10_LC_21_16_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_10_LC_21_16_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_10_LC_21_16_5  (
            .in0(N__46695),
            .in1(_gnd_net_),
            .in2(N__46689),
            .in3(N__55726),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net ),
            .ce(N__55571),
            .sr(N__62900));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI0LFN1_LC_21_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI0LFN1_LC_21_16_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI0LFN1_LC_21_16_6 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI0LFN1_LC_21_16_6  (
            .in0(N__55255),
            .in1(N__55430),
            .in2(N__46667),
            .in3(N__46627),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJQQL2_LC_21_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJQQL2_LC_21_16_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJQQL2_LC_21_16_7 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJQQL2_LC_21_16_7  (
            .in0(N__46660),
            .in1(N__55036),
            .in2(N__46634),
            .in3(N__54834),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_0_4_LC_21_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_0_4_LC_21_17_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_0_4_LC_21_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_0_4_LC_21_17_0  (
            .in0(N__47168),
            .in1(N__47244),
            .in2(N__47122),
            .in3(N__47207),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_3_LC_21_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_3_LC_21_17_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_3_LC_21_17_1 .LUT_INIT=16'b1101010111110101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_3_LC_21_17_1  (
            .in0(N__56127),
            .in1(N__56057),
            .in2(N__46608),
            .in3(N__54335),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_2_LC_21_17_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_2_LC_21_17_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_2_LC_21_17_2 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_2_LC_21_17_2  (
            .in0(N__50545),
            .in1(N__56128),
            .in2(_gnd_net_),
            .in3(N__55916),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_1_LC_21_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_1_LC_21_17_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_1_LC_21_17_3 .LUT_INIT=16'b0101111101001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_1_LC_21_17_3  (
            .in0(N__54402),
            .in1(N__55868),
            .in2(N__46965),
            .in3(N__55796),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_4_LC_21_17_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_4_LC_21_17_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_4_LC_21_17_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_4_LC_21_17_6  (
            .in0(N__47169),
            .in1(N__47245),
            .in2(N__47123),
            .in3(N__47208),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_1_LC_21_18_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_1_LC_21_18_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_1_LC_21_18_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_1_LC_21_18_0  (
            .in0(N__47171),
            .in1(N__46980),
            .in2(N__47124),
            .in3(N__47061),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIOFAP_9_LC_21_18_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIOFAP_9_LC_21_18_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIOFAP_9_LC_21_18_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIOFAP_9_LC_21_18_1  (
            .in0(_gnd_net_),
            .in1(N__47041),
            .in2(_gnd_net_),
            .in3(N__47012),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_3_LC_21_18_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_3_LC_21_18_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_3_LC_21_18_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_3_LC_21_18_2  (
            .in0(N__46813),
            .in1(N__46762),
            .in2(N__46908),
            .in3(N__54337),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_LC_21_18_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_LC_21_18_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_LC_21_18_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_LC_21_18_3  (
            .in0(N__46761),
            .in1(N__46892),
            .in2(_gnd_net_),
            .in3(N__46812),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_0_3_LC_21_18_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_0_3_LC_21_18_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_0_3_LC_21_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_0_3_LC_21_18_4  (
            .in0(N__46974),
            .in1(N__56129),
            .in2(N__46968),
            .in3(N__54336),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_11_LC_21_18_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_11_LC_21_18_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_11_LC_21_18_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_11_LC_21_18_5  (
            .in0(N__46956),
            .in1(N__46946),
            .in2(N__46914),
            .in3(N__47468),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_0_LC_21_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_0_LC_21_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_0_LC_21_18_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_0_LC_21_18_6  (
            .in0(N__46891),
            .in1(N__46811),
            .in2(_gnd_net_),
            .in3(N__46760),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIKPI66_9_LC_21_18_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIKPI66_9_LC_21_18_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIKPI66_9_LC_21_18_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIKPI66_9_LC_21_18_7  (
            .in0(N__47478),
            .in1(N__50192),
            .in2(_gnd_net_),
            .in3(N__47469),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_394 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIGUM51_1_LC_21_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIGUM51_1_LC_21_19_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIGUM51_1_LC_21_19_0 .LUT_INIT=16'b0001010101010101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIGUM51_1_LC_21_19_0  (
            .in0(N__64679),
            .in1(N__56574),
            .in2(N__48222),
            .in3(N__55857),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_1_LC_21_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_1_LC_21_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_1_LC_21_19_1 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_1_LC_21_19_1  (
            .in0(N__55853),
            .in1(_gnd_net_),
            .in2(N__56591),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_8_LC_21_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_8_LC_21_19_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_8_LC_21_19_2 .LUT_INIT=16'b1010000010101111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_8_LC_21_19_2  (
            .in0(N__47445),
            .in1(_gnd_net_),
            .in2(N__47436),
            .in3(N__47426),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_8_LC_21_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_8_LC_21_19_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_8_LC_21_19_3 .LUT_INIT=16'b1101000111100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_8_LC_21_19_3  (
            .in0(N__56123),
            .in1(N__47413),
            .in2(N__47328),
            .in3(N__47325),
            .lcout(s_paddr_I2C_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65678),
            .ce(N__50052),
            .sr(N__65009));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_1_LC_21_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_1_LC_21_19_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_1_LC_21_19_4 .LUT_INIT=16'b0000111110101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_1_LC_21_19_4  (
            .in0(N__47319),
            .in1(_gnd_net_),
            .in2(N__48220),
            .in3(N__55855),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1651 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_2_LC_21_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_2_LC_21_19_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_2_LC_21_19_5 .LUT_INIT=16'b0111011100100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_2_LC_21_19_5  (
            .in0(N__55854),
            .in1(N__48209),
            .in2(_gnd_net_),
            .in3(N__47286),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1652 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_4_LC_21_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_4_LC_21_19_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_4_LC_21_19_6 .LUT_INIT=16'b1010000010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_4_LC_21_19_6  (
            .in0(N__64472),
            .in1(_gnd_net_),
            .in2(N__48221),
            .in3(N__55856),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_4_LC_21_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_4_LC_21_19_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_4_LC_21_19_7 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_4_LC_21_19_7  (
            .in0(N__56489),
            .in1(N__50681),
            .in2(N__47250),
            .in3(N__56469),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_14_LC_21_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_14_LC_21_20_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_14_LC_21_20_0 .LUT_INIT=16'b0111111101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_14_LC_21_20_0  (
            .in0(N__47493),
            .in1(N__56027),
            .in2(N__66609),
            .in3(N__48205),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_14_LC_21_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_14_LC_21_20_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_14_LC_21_20_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_14_LC_21_20_1  (
            .in0(N__66125),
            .in1(N__64696),
            .in2(_gnd_net_),
            .in3(N__50137),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_0_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_17_LC_21_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_17_LC_21_20_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_17_LC_21_20_2 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_17_LC_21_20_2  (
            .in0(N__64697),
            .in1(N__66324),
            .in2(_gnd_net_),
            .in3(N__65914),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_279_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_17_LC_21_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_17_LC_21_20_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_17_LC_21_20_3 .LUT_INIT=16'b0000010000000101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_17_LC_21_20_3  (
            .in0(N__66129),
            .in1(N__66325),
            .in2(N__47487),
            .in3(N__66607),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65687),
            .ce(),
            .sr(N__65012));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_7_LC_21_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_7_LC_21_20_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_7_LC_21_20_5 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_7_LC_21_20_5  (
            .in0(N__66375),
            .in1(N__62406),
            .in2(N__66156),
            .in3(N__50138),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_0_1_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_7_LC_21_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_7_LC_21_20_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_7_LC_21_20_6 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_7_LC_21_20_6  (
            .in0(N__55862),
            .in1(N__56028),
            .in2(N__47484),
            .in3(N__66376),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65687),
            .ce(),
            .sr(N__65012));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_20_LC_21_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_20_LC_21_20_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_20_LC_21_20_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_20_LC_21_20_7  (
            .in0(N__55861),
            .in1(N__50682),
            .in2(N__48219),
            .in3(N__64473),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65687),
            .ce(),
            .sr(N__65012));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_9_LC_21_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_9_LC_21_21_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_9_LC_21_21_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_9_LC_21_21_0  (
            .in0(N__50544),
            .in1(N__50930),
            .in2(N__56520),
            .in3(N__57287),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_268_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_9_LC_21_21_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_9_LC_21_21_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_9_LC_21_21_1 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_9_LC_21_21_1  (
            .in0(N__66603),
            .in1(N__50643),
            .in2(N__47481),
            .in3(N__50166),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65702),
            .ce(),
            .sr(N__65020));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_10_LC_21_21_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_10_LC_21_21_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_10_LC_21_21_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_10_LC_21_21_3  (
            .in0(_gnd_net_),
            .in1(N__50642),
            .in2(_gnd_net_),
            .in3(N__66602),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_10_LC_21_21_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_10_LC_21_21_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_10_LC_21_21_4 .LUT_INIT=16'b0111010100110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_10_LC_21_21_4  (
            .in0(N__66109),
            .in1(N__47510),
            .in2(N__47571),
            .in3(N__66755),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65702),
            .ce(),
            .sr(N__65020));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_18_LC_21_21_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_18_LC_21_21_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_18_LC_21_21_5 .LUT_INIT=16'b0101010111001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_18_LC_21_21_5  (
            .in0(N__50721),
            .in1(N__47564),
            .in2(_gnd_net_),
            .in3(N__50543),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_18_LC_21_21_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_18_LC_21_21_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_18_LC_21_21_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_18_LC_21_21_6  (
            .in0(N__66110),
            .in1(_gnd_net_),
            .in2(N__47568),
            .in3(N__50932),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65702),
            .ce(),
            .sr(N__65020));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_8_LC_21_21_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_8_LC_21_21_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_8_LC_21_21_7 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_8_LC_21_21_7  (
            .in0(N__50931),
            .in1(N__66111),
            .in2(_gnd_net_),
            .in3(N__47565),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65702),
            .ce(),
            .sr(N__65020));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_o2_26_LC_21_22_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_o2_26_LC_21_22_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_o2_26_LC_21_22_0 .LUT_INIT=16'b0000011000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_o2_26_LC_21_22_0  (
            .in0(N__51078),
            .in1(N__51052),
            .in2(N__51023),
            .in3(N__51121),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1605_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_0_0_LC_21_22_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_0_0_LC_21_22_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_0_0_LC_21_22_1 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_0_0_LC_21_22_1  (
            .in0(N__48181),
            .in1(N__51076),
            .in2(_gnd_net_),
            .in3(N__47526),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_0_o2_LC_21_22_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_0_o2_LC_21_22_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_0_o2_LC_21_22_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_0_o2_LC_21_22_2  (
            .in0(N__51013),
            .in1(N__51048),
            .in2(_gnd_net_),
            .in3(N__51118),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_14_LC_21_22_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_14_LC_21_22_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_14_LC_21_22_3 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_14_LC_21_22_3  (
            .in0(N__48183),
            .in1(N__64433),
            .in2(N__47520),
            .in3(N__51079),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_a3_1_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI68137_11_LC_21_22_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI68137_11_LC_21_22_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI68137_11_LC_21_22_4 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI68137_11_LC_21_22_4  (
            .in0(N__56173),
            .in1(N__50004),
            .in2(_gnd_net_),
            .in3(N__48182),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.un1_command_1_i_i_o2_LC_21_22_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.un1_command_1_i_i_o2_LC_21_22_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.un1_command_1_i_i_o2_LC_21_22_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.un1_command_1_i_i_o2_LC_21_22_5  (
            .in0(N__51119),
            .in1(N__51014),
            .in2(N__51054),
            .in3(N__51075),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_o4_1_1_a3_0_o2_4_LC_21_22_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_o4_1_1_a3_0_o2_4_LC_21_22_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_o4_1_1_a3_0_o2_4_LC_21_22_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_o4_1_1_a3_0_o2_4_LC_21_22_7  (
            .in0(N__51120),
            .in1(N__51015),
            .in2(_gnd_net_),
            .in3(N__51077),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_0_LC_21_23_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_0_LC_21_23_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_0_LC_21_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_0_LC_21_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48294),
            .lcout(\I2C_top_level_inst1.s_command_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47996),
            .ce(N__47931),
            .sr(N__62848));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_1_LC_21_23_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_1_LC_21_23_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_1_LC_21_23_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_1_LC_21_23_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48162),
            .lcout(\I2C_top_level_inst1.s_command_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47996),
            .ce(N__47931),
            .sr(N__62848));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_2_LC_21_23_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_2_LC_21_23_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_2_LC_21_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_2_LC_21_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48111),
            .lcout(\I2C_top_level_inst1.s_command_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47996),
            .ce(N__47931),
            .sr(N__62848));
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_3_LC_21_23_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_3_LC_21_23_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.command_reg_inst.c_command_3_LC_21_23_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.command_reg_inst.c_command_3_LC_21_23_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__48056),
            .lcout(\I2C_top_level_inst1.s_command_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__47996),
            .ce(N__47931),
            .sr(N__62848));
    defparam \serializer_mod_inst.counter_sr_RNIO9BB_0_LC_21_25_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.counter_sr_RNIO9BB_0_LC_21_25_3 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.counter_sr_RNIO9BB_0_LC_21_25_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \serializer_mod_inst.counter_sr_RNIO9BB_0_LC_21_25_3  (
            .in0(N__48357),
            .in1(N__48435),
            .in2(_gnd_net_),
            .in3(N__48483),
            .lcout(\serializer_mod_inst.un1_counter_srlto6_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.counter_sr_RNIDF4F_1_LC_21_26_3 .C_ON=1'b0;
    defparam \serializer_mod_inst.counter_sr_RNIDF4F_1_LC_21_26_3 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.counter_sr_RNIDF4F_1_LC_21_26_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \serializer_mod_inst.counter_sr_RNIDF4F_1_LC_21_26_3  (
            .in0(N__48374),
            .in1(N__48392),
            .in2(N__48459),
            .in3(N__48410),
            .lcout(),
            .ltout(\serializer_mod_inst.un1_counter_srlto6_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.counter_sr_RNIREMI1_7_LC_21_26_4 .C_ON=1'b0;
    defparam \serializer_mod_inst.counter_sr_RNIREMI1_7_LC_21_26_4 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.counter_sr_RNIREMI1_7_LC_21_26_4 .LUT_INIT=16'b1101010111111111;
    LogicCell40 \serializer_mod_inst.counter_sr_RNIREMI1_7_LC_21_26_4  (
            .in0(N__48617),
            .in1(N__47892),
            .in2(N__47886),
            .in3(N__47644),
            .lcout(\serializer_mod_inst.counter_sre_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.current_state_RNO_2_0_LC_21_26_5 .C_ON=1'b0;
    defparam \serializer_mod_inst.current_state_RNO_2_0_LC_21_26_5 .SEQ_MODE=4'b0000;
    defparam \serializer_mod_inst.current_state_RNO_2_0_LC_21_26_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \serializer_mod_inst.current_state_RNO_2_0_LC_21_26_5  (
            .in0(N__48373),
            .in1(N__48391),
            .in2(N__48356),
            .in3(N__48409),
            .lcout(\serializer_mod_inst.un22_next_state_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \serializer_mod_inst.counter_sr_0_LC_21_27_0 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_0_LC_21_27_0 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_0_LC_21_27_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_0_LC_21_27_0  (
            .in0(N__48651),
            .in1(N__48482),
            .in2(_gnd_net_),
            .in3(N__48462),
            .lcout(\serializer_mod_inst.counter_srZ0Z_0 ),
            .ltout(),
            .carryin(bfn_21_27_0_),
            .carryout(\serializer_mod_inst.counter_sr_cry_0 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_1_LC_21_27_1 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_1_LC_21_27_1 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_1_LC_21_27_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_1_LC_21_27_1  (
            .in0(N__48638),
            .in1(N__48457),
            .in2(_gnd_net_),
            .in3(N__48438),
            .lcout(\serializer_mod_inst.counter_srZ0Z_1 ),
            .ltout(),
            .carryin(\serializer_mod_inst.counter_sr_cry_0 ),
            .carryout(\serializer_mod_inst.counter_sr_cry_1 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_2_LC_21_27_2 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_2_LC_21_27_2 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_2_LC_21_27_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_2_LC_21_27_2  (
            .in0(N__48652),
            .in1(N__48434),
            .in2(_gnd_net_),
            .in3(N__48414),
            .lcout(\serializer_mod_inst.counter_srZ0Z_2 ),
            .ltout(),
            .carryin(\serializer_mod_inst.counter_sr_cry_1 ),
            .carryout(\serializer_mod_inst.counter_sr_cry_2 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_3_LC_21_27_3 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_3_LC_21_27_3 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_3_LC_21_27_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_3_LC_21_27_3  (
            .in0(N__48639),
            .in1(N__48411),
            .in2(_gnd_net_),
            .in3(N__48396),
            .lcout(\serializer_mod_inst.counter_srZ0Z_3 ),
            .ltout(),
            .carryin(\serializer_mod_inst.counter_sr_cry_2 ),
            .carryout(\serializer_mod_inst.counter_sr_cry_3 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_4_LC_21_27_4 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_4_LC_21_27_4 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_4_LC_21_27_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_4_LC_21_27_4  (
            .in0(N__48653),
            .in1(N__48393),
            .in2(_gnd_net_),
            .in3(N__48378),
            .lcout(\serializer_mod_inst.counter_srZ0Z_4 ),
            .ltout(),
            .carryin(\serializer_mod_inst.counter_sr_cry_3 ),
            .carryout(\serializer_mod_inst.counter_sr_cry_4 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_5_LC_21_27_5 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_5_LC_21_27_5 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_5_LC_21_27_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_5_LC_21_27_5  (
            .in0(N__48640),
            .in1(N__48375),
            .in2(_gnd_net_),
            .in3(N__48360),
            .lcout(\serializer_mod_inst.counter_srZ0Z_5 ),
            .ltout(),
            .carryin(\serializer_mod_inst.counter_sr_cry_4 ),
            .carryout(\serializer_mod_inst.counter_sr_cry_5 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_6_LC_21_27_6 .C_ON=1'b1;
    defparam \serializer_mod_inst.counter_sr_6_LC_21_27_6 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_6_LC_21_27_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_6_LC_21_27_6  (
            .in0(N__48654),
            .in1(N__48355),
            .in2(_gnd_net_),
            .in3(N__48333),
            .lcout(\serializer_mod_inst.counter_srZ0Z_6 ),
            .ltout(),
            .carryin(\serializer_mod_inst.counter_sr_cry_5 ),
            .carryout(\serializer_mod_inst.counter_sr_cry_6 ),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \serializer_mod_inst.counter_sr_7_LC_21_27_7 .C_ON=1'b0;
    defparam \serializer_mod_inst.counter_sr_7_LC_21_27_7 .SEQ_MODE=4'b1010;
    defparam \serializer_mod_inst.counter_sr_7_LC_21_27_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \serializer_mod_inst.counter_sr_7_LC_21_27_7  (
            .in0(N__48641),
            .in1(N__48618),
            .in2(_gnd_net_),
            .in3(N__48621),
            .lcout(\serializer_mod_inst.counter_srZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65754),
            .ce(N__48600),
            .sr(N__62827));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_15_LC_22_9_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_15_LC_22_9_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_15_LC_22_9_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_15_LC_22_9_0  (
            .in0(_gnd_net_),
            .in1(N__57524),
            .in2(_gnd_net_),
            .in3(N__59708),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_24_LC_22_9_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_24_LC_22_9_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_24_LC_22_9_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_24_LC_22_9_1  (
            .in0(N__59712),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61113),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_16_LC_22_9_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_16_LC_22_9_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_16_LC_22_9_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_16_LC_22_9_2  (
            .in0(_gnd_net_),
            .in1(N__59709),
            .in2(_gnd_net_),
            .in3(N__57627),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_25_LC_22_9_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_25_LC_22_9_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_25_LC_22_9_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_25_LC_22_9_3  (
            .in0(N__59713),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60981),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_17_LC_22_9_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_17_LC_22_9_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_17_LC_22_9_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_17_LC_22_9_4  (
            .in0(_gnd_net_),
            .in1(N__59710),
            .in2(_gnd_net_),
            .in3(N__57413),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_26_LC_22_9_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_26_LC_22_9_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_26_LC_22_9_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_26_LC_22_9_5  (
            .in0(N__59714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60897),
            .lcout(\cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_2Z0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_18_LC_22_9_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_18_LC_22_9_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_18_LC_22_9_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_18_LC_22_9_6  (
            .in0(_gnd_net_),
            .in1(N__59711),
            .in2(_gnd_net_),
            .in3(N__59865),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_27_LC_22_9_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_27_LC_22_9_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_27_LC_22_9_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_27_LC_22_9_7  (
            .in0(N__59715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__60786),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65568),
            .ce(N__48726),
            .sr(N__62955));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_19_LC_22_10_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_19_LC_22_10_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_19_LC_22_10_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_19_LC_22_10_0  (
            .in0(_gnd_net_),
            .in1(N__61645),
            .in2(_gnd_net_),
            .in3(N__59593),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65580),
            .ce(N__48725),
            .sr(N__62952));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_28_LC_22_10_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_28_LC_22_10_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_28_LC_22_10_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_28_LC_22_10_1  (
            .in0(N__59596),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62367),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65580),
            .ce(N__48725),
            .sr(N__62952));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_29_LC_22_10_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_29_LC_22_10_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_29_LC_22_10_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_29_LC_22_10_2  (
            .in0(N__62262),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59597),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65580),
            .ce(N__48725),
            .sr(N__62952));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_0_LC_22_10_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_0_LC_22_10_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_0_LC_22_10_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_0_LC_22_10_3  (
            .in0(N__59595),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61943),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65580),
            .ce(N__48725),
            .sr(N__62952));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_7_LC_22_10_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_7_LC_22_10_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_7_LC_22_10_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_7_LC_22_10_4  (
            .in0(_gnd_net_),
            .in1(N__63482),
            .in2(_gnd_net_),
            .in3(N__59594),
            .lcout(cemf_module_64ch_ctrl_inst1_data_interrupts_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65580),
            .ce(N__48725),
            .sr(N__62952));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI23RI1_LC_22_11_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI23RI1_LC_22_11_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI23RI1_LC_22_11_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI23RI1_LC_22_11_0  (
            .in0(N__55228),
            .in1(N__55455),
            .in2(N__48677),
            .in3(N__48694),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIL86H2_LC_22_11_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIL86H2_LC_22_11_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIL86H2_LC_22_11_1 .LUT_INIT=16'b1101110100001101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIL86H2_LC_22_11_1  (
            .in0(N__48670),
            .in1(N__55057),
            .in2(N__48701),
            .in3(N__54832),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_19_LC_22_11_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_19_LC_22_11_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_19_LC_22_11_2 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_19_LC_22_11_2  (
            .in0(_gnd_net_),
            .in1(N__61646),
            .in2(_gnd_net_),
            .in3(N__59599),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65591),
            .ce(N__49095),
            .sr(N__62947));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIE2FN1_LC_22_11_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIE2FN1_LC_22_11_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIE2FN1_LC_22_11_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIE2FN1_LC_22_11_3  (
            .in0(N__55454),
            .in1(N__55229),
            .in2(N__48914),
            .in3(N__48934),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_0_LC_22_11_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_0_LC_22_11_4 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_0_LC_22_11_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_0_LC_22_11_4  (
            .in0(_gnd_net_),
            .in1(N__61969),
            .in2(_gnd_net_),
            .in3(N__59598),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65591),
            .ce(N__49095),
            .sr(N__62947));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI18QL2_LC_22_11_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI18QL2_LC_22_11_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI18QL2_LC_22_11_5 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI18QL2_LC_22_11_5  (
            .in0(N__54833),
            .in1(N__48935),
            .in2(N__55062),
            .in3(N__48910),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQL7_LC_22_11_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQL7_LC_22_11_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQL7_LC_22_11_6 .LUT_INIT=16'b0111111100111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQL7_LC_22_11_6  (
            .in0(N__54006),
            .in1(N__48891),
            .in2(N__48885),
            .in3(N__58223),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIJ0CO7_LC_22_11_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIJ0CO7_LC_22_11_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIJ0CO7_LC_22_11_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIJ0CO7_LC_22_11_7  (
            .in0(N__53718),
            .in1(_gnd_net_),
            .in2(N__48882),
            .in3(N__48879),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI01RI1_LC_22_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI01RI1_LC_22_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI01RI1_LC_22_12_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI01RI1_LC_22_12_0  (
            .in0(N__55263),
            .in1(N__55445),
            .in2(N__48867),
            .in3(N__49156),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJ66H2_LC_22_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJ66H2_LC_22_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJ66H2_LC_22_12_1 .LUT_INIT=16'b1100111101000101;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJ66H2_LC_22_12_1  (
            .in0(N__48866),
            .in1(N__55058),
            .in2(N__49163),
            .in3(N__54837),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579D7_LC_22_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579D7_LC_22_12_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579D7_LC_22_12_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579D7_LC_22_12_2  (
            .in0(N__53962),
            .in1(N__51395),
            .in2(N__48837),
            .in3(N__48834),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIGAQF7_LC_22_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIGAQF7_LC_22_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIGAQF7_LC_22_12_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIGAQF7_LC_22_12_3  (
            .in0(_gnd_net_),
            .in1(N__53716),
            .in2(N__48828),
            .in3(N__48825),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18_LC_22_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18_LC_22_12_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18_LC_22_12_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18_LC_22_12_4  (
            .in0(_gnd_net_),
            .in1(N__48819),
            .in2(N__48813),
            .in3(N__55745),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net ),
            .ce(N__55559),
            .sr(N__62941));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9D7_LC_22_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9D7_LC_22_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9D7_LC_22_12_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9D7_LC_22_12_5  (
            .in0(N__53948),
            .in1(N__51476),
            .in2(N__48810),
            .in3(N__48801),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9DZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILFQF7_LC_22_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILFQF7_LC_22_12_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILFQF7_LC_22_12_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILFQF7_LC_22_12_6  (
            .in0(N__53717),
            .in1(_gnd_net_),
            .in2(N__49209),
            .in3(N__49206),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_19_LC_22_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_19_LC_22_12_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_19_LC_22_12_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_19_LC_22_12_7  (
            .in0(N__55746),
            .in1(_gnd_net_),
            .in2(N__49200),
            .in3(N__49197),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net ),
            .ce(N__55559),
            .sr(N__62941));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_18_LC_22_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_18_LC_22_13_0 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_18_LC_22_13_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_18_LC_22_13_0  (
            .in0(N__59505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59853),
            .lcout(cemf_module_64ch_ctrl_inst1_data_clkctrovf_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65611),
            .ce(N__49094),
            .sr(N__62936));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_27_LC_22_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_27_LC_22_13_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_27_LC_22_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_27_LC_22_13_1  (
            .in0(_gnd_net_),
            .in1(N__59504),
            .in2(_gnd_net_),
            .in3(N__60806),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65611),
            .ce(N__49094),
            .sr(N__62936));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_28_LC_22_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_28_LC_22_13_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_28_LC_22_13_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_28_LC_22_13_2  (
            .in0(N__59506),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62356),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65611),
            .ce(N__49094),
            .sr(N__62936));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_29_LC_22_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_29_LC_22_13_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_29_LC_22_13_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_29_LC_22_13_3  (
            .in0(N__62263),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59507),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65611),
            .ce(N__49094),
            .sr(N__62936));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI06692_17_LC_22_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI06692_17_LC_22_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI06692_17_LC_22_14_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI06692_17_LC_22_14_0  (
            .in0(N__57926),
            .in1(N__58184),
            .in2(N__49008),
            .in3(N__51241),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLH5_LC_22_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLH5_LC_22_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLH5_LC_22_14_1 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLH5_LC_22_14_1  (
            .in0(N__60598),
            .in1(N__48975),
            .in2(N__48945),
            .in3(N__49437),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITTFV5_LC_22_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITTFV5_LC_22_14_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITTFV5_LC_22_14_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITTFV5_LC_22_14_2  (
            .in0(N__60379),
            .in1(_gnd_net_),
            .in2(N__49572),
            .in3(N__49569),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23_LC_22_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23_LC_22_14_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23_LC_22_14_3 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23_LC_22_14_3  (
            .in0(_gnd_net_),
            .in1(N__49503),
            .in2(N__49563),
            .in3(N__60196),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.dout_conf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net ),
            .ce(N__60023),
            .sr(N__62927));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOOFV5_LC_22_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOOFV5_LC_22_14_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOOFV5_LC_22_14_4 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOOFV5_LC_22_14_4  (
            .in0(N__60378),
            .in1(N__49527),
            .in2(N__49539),
            .in3(_gnd_net_),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_22_LC_22_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_22_LC_22_14_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_22_LC_22_14_5 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_22_LC_22_14_5  (
            .in0(_gnd_net_),
            .in1(N__49521),
            .in2(N__49506),
            .in3(N__60195),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net ),
            .ce(N__60023),
            .sr(N__62927));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOQSI1_LC_22_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOQSI1_LC_22_14_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOQSI1_LC_22_14_6 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOQSI1_LC_22_14_6  (
            .in0(N__55453),
            .in1(N__55156),
            .in2(N__49493),
            .in3(N__49454),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI81C92_17_LC_22_15_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI81C92_17_LC_22_15_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI81C92_17_LC_22_15_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI81C92_17_LC_22_15_0  (
            .in0(N__58182),
            .in1(N__57989),
            .in2(N__49431),
            .in3(N__49378),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOR392_17_LC_22_15_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOR392_17_LC_22_15_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOR392_17_LC_22_15_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOR392_17_LC_22_15_1  (
            .in0(N__57990),
            .in1(N__58183),
            .in2(N__49339),
            .in3(N__49308),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFH5_LC_22_15_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFH5_LC_22_15_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFH5_LC_22_15_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFH5_LC_22_15_2  (
            .in0(N__60618),
            .in1(N__49268),
            .in2(N__49233),
            .in3(N__49230),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI94AV5_LC_22_15_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI94AV5_LC_22_15_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI94AV5_LC_22_15_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI94AV5_LC_22_15_3  (
            .in0(N__60377),
            .in1(_gnd_net_),
            .in2(N__49218),
            .in3(N__49215),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10_LC_22_15_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10_LC_22_15_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10_LC_22_15_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10_LC_22_15_4  (
            .in0(N__60193),
            .in1(_gnd_net_),
            .in2(N__49860),
            .in3(N__49758),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net ),
            .ce(N__60022),
            .sr(N__62919));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044Q5_LC_22_15_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044Q5_LC_22_15_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044Q5_LC_22_15_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044Q5_LC_22_15_5  (
            .in0(N__60617),
            .in1(N__49832),
            .in2(N__49803),
            .in3(N__49791),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1IU76_LC_22_15_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1IU76_LC_22_15_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1IU76_LC_22_15_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1IU76_LC_22_15_6  (
            .in0(_gnd_net_),
            .in1(N__60376),
            .in2(N__49785),
            .in3(N__49782),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_9_LC_22_15_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_9_LC_22_15_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_9_LC_22_15_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_9_LC_22_15_7  (
            .in0(_gnd_net_),
            .in1(N__49776),
            .in2(N__49761),
            .in3(N__60194),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net ),
            .ce(N__60022),
            .sr(N__62919));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQIB92_17_LC_22_16_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQIB92_17_LC_22_16_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQIB92_17_LC_22_16_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQIB92_17_LC_22_16_0  (
            .in0(N__58013),
            .in1(N__58110),
            .in2(N__53793),
            .in3(N__49751),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISKB92_17_LC_22_16_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISKB92_17_LC_22_16_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISKB92_17_LC_22_16_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISKB92_17_LC_22_16_1  (
            .in0(N__58111),
            .in1(N__58014),
            .in2(N__49718),
            .in3(N__49677),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253Q5_LC_22_16_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253Q5_LC_22_16_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253Q5_LC_22_16_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253Q5_LC_22_16_2  (
            .in0(N__60605),
            .in1(N__49637),
            .in2(N__49599),
            .in3(N__49596),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI3JT76_LC_22_16_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI3JT76_LC_22_16_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI3JT76_LC_22_16_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI3JT76_LC_22_16_3  (
            .in0(_gnd_net_),
            .in1(N__60374),
            .in2(N__49581),
            .in3(N__49578),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3_LC_22_16_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3_LC_22_16_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3_LC_22_16_4 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3_LC_22_16_4  (
            .in0(_gnd_net_),
            .in1(N__49905),
            .in2(N__49986),
            .in3(N__60167),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net ),
            .ce(N__60018),
            .sr(N__62911));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2Q5_LC_22_16_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2Q5_LC_22_16_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2Q5_LC_22_16_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2Q5_LC_22_16_5  (
            .in0(N__60612),
            .in1(N__49961),
            .in2(N__49935),
            .in3(N__49926),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIUDT76_LC_22_16_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIUDT76_LC_22_16_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIUDT76_LC_22_16_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIUDT76_LC_22_16_6  (
            .in0(N__60375),
            .in1(_gnd_net_),
            .in2(N__49917),
            .in3(N__49914),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_2_LC_22_16_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_2_LC_22_16_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_2_LC_22_16_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_2_LC_22_16_7  (
            .in0(N__60166),
            .in1(_gnd_net_),
            .in2(N__49908),
            .in3(N__60657),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net ),
            .ce(N__60018),
            .sr(N__62911));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_2_LC_22_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_2_LC_22_17_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_2_LC_22_17_0 .LUT_INIT=16'b1111111101001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_2_LC_22_17_0  (
            .in0(N__54403),
            .in1(N__56726),
            .in2(N__50196),
            .in3(N__56447),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_2_LC_22_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_2_LC_22_17_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_2_LC_22_17_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_2_LC_22_17_1  (
            .in0(N__50218),
            .in1(N__50611),
            .in2(N__49893),
            .in3(N__50050),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65662),
            .ce(),
            .sr(N__65004));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_3_LC_22_17_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_3_LC_22_17_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_3_LC_22_17_2 .LUT_INIT=16'b1111011110000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_3_LC_22_17_2  (
            .in0(N__50051),
            .in1(N__50219),
            .in2(N__54231),
            .in3(N__55943),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65662),
            .ce(),
            .sr(N__65004));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_15_LC_22_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_15_LC_22_17_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_15_LC_22_17_3 .LUT_INIT=16'b0000000001110101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_15_LC_22_17_3  (
            .in0(N__56725),
            .in1(N__50015),
            .in2(N__54405),
            .in3(N__49890),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_15_LC_22_17_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_15_LC_22_17_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_15_LC_22_17_4 .LUT_INIT=16'b1101000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_15_LC_22_17_4  (
            .in0(N__50140),
            .in1(N__50175),
            .in2(N__49878),
            .in3(N__56446),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_1_LC_22_17_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_1_LC_22_17_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_1_LC_22_17_5 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_1_LC_22_17_5  (
            .in0(N__54237),
            .in1(N__55964),
            .in2(N__50220),
            .in3(N__50049),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65662),
            .ce(),
            .sr(N__65004));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_3_LC_22_17_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_3_LC_22_17_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_3_LC_22_17_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_3_LC_22_17_6  (
            .in0(_gnd_net_),
            .in1(N__50191),
            .in2(_gnd_net_),
            .in3(N__54398),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIMJR28_26_LC_22_17_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIMJR28_26_LC_22_17_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIMJR28_26_LC_22_17_7 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIMJR28_26_LC_22_17_7  (
            .in0(N__55864),
            .in1(N__56448),
            .in2(N__50169),
            .in3(N__50139),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIJU6F7_23_LC_22_18_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIJU6F7_23_LC_22_18_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIJU6F7_23_LC_22_18_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIJU6F7_23_LC_22_18_1  (
            .in0(N__50016),
            .in1(N__54404),
            .in2(_gnd_net_),
            .in3(N__56718),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_267 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_267_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAOTPE_26_LC_22_18_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAOTPE_26_LC_22_18_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAOTPE_26_LC_22_18_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAOTPE_26_LC_22_18_2  (
            .in0(N__50154),
            .in1(N__56439),
            .in2(N__50148),
            .in3(N__50141),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIC372_3_LC_22_18_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIC372_3_LC_22_18_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIC372_3_LC_22_18_3 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIC372_3_LC_22_18_3  (
            .in0(N__54251),
            .in1(N__56056),
            .in2(_gnd_net_),
            .in3(N__54342),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_1_1_i_m2_1_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIDH244_3_LC_22_18_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIDH244_3_LC_22_18_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIDH244_3_LC_22_18_4 .LUT_INIT=16'b1011001100000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIDH244_3_LC_22_18_4  (
            .in0(N__54343),
            .in1(N__54419),
            .in2(N__50019),
            .in3(N__56130),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_101 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_2_LC_22_18_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_2_LC_22_18_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_2_LC_22_18_7 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_2_LC_22_18_7  (
            .in0(N__49997),
            .in1(N__56360),
            .in2(N__64737),
            .in3(N__55929),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1802 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_0_2_LC_22_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_0_2_LC_22_19_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_0_2_LC_22_19_0 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_0_2_LC_22_19_0  (
            .in0(N__50714),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66118),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_904 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_0_LC_22_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_0_LC_22_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_0_LC_22_19_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_0_LC_22_19_1  (
            .in0(N__56358),
            .in1(_gnd_net_),
            .in2(N__66155),
            .in3(N__64420),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_1_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_0_LC_22_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_0_LC_22_19_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_0_LC_22_19_2 .LUT_INIT=16'b1111111101000101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_0_LC_22_19_2  (
            .in0(N__56512),
            .in1(N__50551),
            .in2(N__50469),
            .in3(N__57209),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3TI11_2_LC_22_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3TI11_2_LC_22_19_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3TI11_2_LC_22_19_3 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3TI11_2_LC_22_19_3  (
            .in0(N__56357),
            .in1(_gnd_net_),
            .in2(N__66154),
            .in3(N__50715),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_7_14_LC_22_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_7_14_LC_22_19_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_7_14_LC_22_19_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_7_14_LC_22_19_4  (
            .in0(_gnd_net_),
            .in1(N__64316),
            .in2(N__50466),
            .in3(N__64265),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_14_LC_22_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_14_LC_22_19_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_14_LC_22_19_5 .LUT_INIT=16'b0000010000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_14_LC_22_19_5  (
            .in0(N__50581),
            .in1(N__50226),
            .in2(N__50463),
            .in3(N__50460),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_412_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_14_LC_22_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_14_LC_22_19_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_14_LC_22_19_6 .LUT_INIT=16'b1010101110111011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_14_LC_22_19_6  (
            .in0(N__50766),
            .in1(N__50427),
            .in2(N__50418),
            .in3(N__50415),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65688),
            .ce(),
            .sr(N__65013));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_14_LC_22_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_14_LC_22_19_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_14_LC_22_19_7 .LUT_INIT=16'b0011001101111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_14_LC_22_19_7  (
            .in0(N__56359),
            .in1(N__56511),
            .in2(N__50386),
            .in3(N__64421),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_1_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_25_LC_22_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_25_LC_22_20_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_25_LC_22_20_0 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_25_LC_22_20_0  (
            .in0(N__50923),
            .in1(N__50631),
            .in2(N__57014),
            .in3(N__66453),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65703),
            .ce(),
            .sr(N__65021));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_RNISQP11_2_LC_22_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_RNISQP11_2_LC_22_20_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_RNISQP11_2_LC_22_20_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_RNISQP11_2_LC_22_20_1  (
            .in0(N__65852),
            .in1(N__50666),
            .in2(N__65932),
            .in3(N__66020),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9FLC_24_LC_22_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9FLC_24_LC_22_20_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9FLC_24_LC_22_20_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9FLC_24_LC_22_20_3  (
            .in0(_gnd_net_),
            .in1(N__50921),
            .in2(_gnd_net_),
            .in3(N__57029),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_25_LC_22_20_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_25_LC_22_20_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_25_LC_22_20_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_25_LC_22_20_4  (
            .in0(N__66560),
            .in1(N__57002),
            .in2(N__50634),
            .in3(N__66691),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_24_LC_22_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_24_LC_22_20_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_24_LC_22_20_5 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_24_LC_22_20_5  (
            .in0(N__66608),
            .in1(N__50922),
            .in2(N__57013),
            .in3(N__57030),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_24_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_24_LC_22_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_24_LC_22_20_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_24_LC_22_20_6 .LUT_INIT=16'b0100111100001111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_24_LC_22_20_6  (
            .in0(N__50621),
            .in1(N__50585),
            .in2(N__50565),
            .in3(N__55920),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65703),
            .ce(),
            .sr(N__65021));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_14_LC_22_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_14_LC_22_20_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_14_LC_22_20_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_14_LC_22_20_7  (
            .in0(N__65926),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__66021),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_86_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_11_LC_22_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_11_LC_22_21_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_11_LC_22_21_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_11_LC_22_21_0  (
            .in0(_gnd_net_),
            .in1(N__66093),
            .in2(_gnd_net_),
            .in3(N__66554),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_11_LC_22_21_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_11_LC_22_21_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_11_LC_22_21_1 .LUT_INIT=16'b0111000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_11_LC_22_21_1  (
            .in0(N__50717),
            .in1(N__50538),
            .in2(N__50562),
            .in3(N__64788),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_11_LC_22_21_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_11_LC_22_21_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_11_LC_22_21_2 .LUT_INIT=16'b0101000001100000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_11_LC_22_21_2  (
            .in0(N__50539),
            .in1(N__66680),
            .in2(N__50493),
            .in3(N__66503),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_1_LC_22_21_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_1_LC_22_21_3 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_1_LC_22_21_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_1_LC_22_21_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50727),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65720),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_14_LC_22_21_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_14_LC_22_21_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_14_LC_22_21_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_14_LC_22_21_4  (
            .in0(N__66105),
            .in1(N__65848),
            .in2(N__50775),
            .in3(N__50667),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_95_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_0_LC_22_21_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_0_LC_22_21_5 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_0_LC_22_21_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_0_LC_22_21_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50757),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65720),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_2_LC_22_21_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_2_LC_22_21_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_2_LC_22_21_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_2_LC_22_21_6  (
            .in0(_gnd_net_),
            .in1(N__50716),
            .in2(_gnd_net_),
            .in3(N__66094),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_844_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_2_LC_22_21_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_2_LC_22_21_7 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_2_LC_22_21_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_2_LC_22_21_7  (
            .in0(N__50655),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65720),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_i_o2_LC_22_22_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_i_o2_LC_22_22_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_i_o2_LC_22_22_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_i_o2_LC_22_22_0  (
            .in0(N__51080),
            .in1(N__51044),
            .in2(N__51024),
            .in3(N__51122),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_1_LC_22_22_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_1_LC_22_22_1 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_1_LC_22_22_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_1_LC_22_22_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57642),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65729),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_2_LC_22_22_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_2_LC_22_22_2 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_2_LC_22_22_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_2_LC_22_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50649),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65729),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_1_LC_22_22_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_1_LC_22_22_3 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_1_LC_22_22_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_1_LC_22_22_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51129),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65729),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQUIH_10_LC_22_22_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQUIH_10_LC_22_22_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQUIH_10_LC_22_22_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQUIH_10_LC_22_22_4  (
            .in0(_gnd_net_),
            .in1(N__66095),
            .in2(_gnd_net_),
            .in3(N__64787),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1754_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_2_LC_22_22_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_2_LC_22_22_5 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_2_LC_22_22_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_2_LC_22_22_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51213),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65729),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_0_LC_22_22_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_0_LC_22_22_6 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_0_LC_22_22_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_0_LC_22_22_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51206),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65729),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6_0_a2_LC_22_22_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6_0_a2_LC_22_22_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6_0_a2_LC_22_22_7 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6_0_a2_LC_22_22_7  (
            .in0(N__51123),
            .in1(N__51081),
            .in2(N__51053),
            .in3(N__51022),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_0_LC_22_23_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_0_LC_22_23_0 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_0_LC_22_23_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_0_LC_22_23_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50993),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65739),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_1_LC_22_23_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_1_LC_22_23_1 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_1_LC_22_23_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_1_LC_22_23_1  (
            .in0(N__50955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65739),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_2_LC_22_23_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_2_LC_22_23_2 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_2_LC_22_23_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_2_LC_22_23_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50949),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65739),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_1_LC_22_23_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_1_LC_22_23_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_1_LC_22_23_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_1_LC_22_23_4  (
            .in0(N__66383),
            .in1(N__66789),
            .in2(N__66693),
            .in3(N__66412),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1666 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_2_LC_22_23_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_2_LC_22_23_5 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_2_LC_22_23_5 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_2_LC_22_23_5  (
            .in0(_gnd_net_),
            .in1(N__51309),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65739),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_0_LC_22_23_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_0_LC_22_23_6 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_0_LC_22_23_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_0_LC_22_23_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__50882),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65739),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_6_0_LC_22_23_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_6_0_LC_22_23_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_6_0_LC_22_23_7 .LUT_INIT=16'b1111111000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_6_0_LC_22_23_7  (
            .in0(N__66790),
            .in1(N__66382),
            .in2(N__66419),
            .in3(N__66504),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_122_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_1_LC_22_24_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_1_LC_22_24_0 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_1_LC_22_24_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_1_LC_22_24_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51285),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65747),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_0_LC_22_24_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_0_LC_22_24_1 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_0_LC_22_24_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_0_LC_22_24_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__51303),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65747),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_18_LC_23_9_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_18_LC_23_9_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_18_LC_23_9_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_18_LC_23_9_0  (
            .in0(N__59672),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59864),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_18),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65581),
            .ce(N__54123),
            .sr(N__62958));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_27_LC_23_9_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_27_LC_23_9_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_27_LC_23_9_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_27_LC_23_9_1  (
            .in0(_gnd_net_),
            .in1(N__59675),
            .in2(_gnd_net_),
            .in3(N__60787),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_27),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65581),
            .ce(N__54123),
            .sr(N__62958));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_19_LC_23_9_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_19_LC_23_9_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_19_LC_23_9_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_19_LC_23_9_2  (
            .in0(N__59673),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61631),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65581),
            .ce(N__54123),
            .sr(N__62958));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_25_LC_23_9_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_25_LC_23_9_3 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_25_LC_23_9_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_25_LC_23_9_3  (
            .in0(N__60980),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__59676),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65581),
            .ce(N__54123),
            .sr(N__62958));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_29_LC_23_9_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_29_LC_23_9_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_29_LC_23_9_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_29_LC_23_9_4  (
            .in0(N__59674),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__62246),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65581),
            .ce(N__54123),
            .sr(N__62958));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_23_LC_23_9_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_23_LC_23_9_5 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_23_LC_23_9_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_23_LC_23_9_5  (
            .in0(_gnd_net_),
            .in1(N__59671),
            .in2(_gnd_net_),
            .in3(N__61242),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_23),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65581),
            .ce(N__54123),
            .sr(N__62958));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HH5_LC_23_10_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HH5_LC_23_10_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HH5_LC_23_10_0 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HH5_LC_23_10_0  (
            .in0(N__57319),
            .in1(N__60614),
            .in2(N__51447),
            .in3(N__51543),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIMIBV5_LC_23_10_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIMIBV5_LC_23_10_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIMIBV5_LC_23_10_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIMIBV5_LC_23_10_1  (
            .in0(N__60385),
            .in1(_gnd_net_),
            .in2(N__51537),
            .in3(N__51534),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19_LC_23_10_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19_LC_23_10_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19_LC_23_10_2 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19_LC_23_10_2  (
            .in0(N__60207),
            .in1(_gnd_net_),
            .in2(N__51528),
            .in3(N__51315),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net ),
            .ce(N__60017),
            .sr(N__62956));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIAE492_17_LC_23_10_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIAE492_17_LC_23_10_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIAE492_17_LC_23_10_3 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIAE492_17_LC_23_10_3  (
            .in0(N__58006),
            .in1(N__58199),
            .in2(N__51506),
            .in3(N__51463),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI8C492_17_LC_23_10_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI8C492_17_LC_23_10_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI8C492_17_LC_23_10_4 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI8C492_17_LC_23_10_4  (
            .in0(N__58200),
            .in1(N__58007),
            .in2(N__51430),
            .in3(N__51382),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGH5_LC_23_10_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGH5_LC_23_10_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGH5_LC_23_10_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGH5_LC_23_10_5  (
            .in0(N__60613),
            .in1(N__51369),
            .in2(N__51342),
            .in3(N__51339),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIHDBV5_LC_23_10_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIHDBV5_LC_23_10_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIHDBV5_LC_23_10_6 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIHDBV5_LC_23_10_6  (
            .in0(_gnd_net_),
            .in1(N__60384),
            .in2(N__51327),
            .in3(N__51324),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_18_LC_23_10_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_18_LC_23_10_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_18_LC_23_10_7 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_18_LC_23_10_7  (
            .in0(_gnd_net_),
            .in1(N__53535),
            .in2(N__51318),
            .in3(N__60206),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net ),
            .ce(N__60017),
            .sr(N__62956));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_25_LC_23_11_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_25_LC_23_11_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_25_LC_23_11_0 .LUT_INIT=16'b0000011101110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_25_LC_23_11_0  (
            .in0(N__53340),
            .in1(N__53266),
            .in2(N__53034),
            .in3(N__53009),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_25_LC_23_11_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_25_LC_23_11_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_25_LC_23_11_1 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_25_LC_23_11_1  (
            .in0(N__52803),
            .in1(N__52782),
            .in2(N__52548),
            .in3(N__52525),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_25_LC_23_11_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_25_LC_23_11_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_25_LC_23_11_2 .LUT_INIT=16'b0011000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_25_LC_23_11_2  (
            .in0(_gnd_net_),
            .in1(N__52254),
            .in2(N__52239),
            .in3(N__52235),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_25_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_25_LC_23_11_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_25_LC_23_11_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_25_LC_23_11_3 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_25_LC_23_11_3  (
            .in0(N__51984),
            .in1(N__51975),
            .in2(N__51969),
            .in3(N__51663),
            .lcout(I2C_top_level_inst1_s_data_oreg_25),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65604),
            .ce(N__54495),
            .sr(N__65024));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_25_LC_23_11_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_25_LC_23_11_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_25_LC_23_11_4 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_25_LC_23_11_4  (
            .in0(N__51966),
            .in1(N__51923),
            .in2(N__51684),
            .in3(N__51672),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI48492_17_LC_23_12_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI48492_17_LC_23_12_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI48492_17_LC_23_12_0 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI48492_17_LC_23_12_0  (
            .in0(N__58196),
            .in1(N__57991),
            .in2(N__51656),
            .in3(N__54193),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6A492_17_LC_23_12_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6A492_17_LC_23_12_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6A492_17_LC_23_12_1 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6A492_17_LC_23_12_1  (
            .in0(N__57992),
            .in1(N__58197),
            .in2(N__51620),
            .in3(N__54142),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGH5_LC_23_12_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGH5_LC_23_12_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGH5_LC_23_12_2 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGH5_LC_23_12_2  (
            .in0(N__51587),
            .in1(N__60590),
            .in2(N__51555),
            .in3(N__51552),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIC8BV5_LC_23_12_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIC8BV5_LC_23_12_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIC8BV5_LC_23_12_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIC8BV5_LC_23_12_3  (
            .in0(_gnd_net_),
            .in1(N__60383),
            .in2(N__53547),
            .in3(N__53544),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17_LC_23_12_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17_LC_23_12_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17_LC_23_12_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17_LC_23_12_4  (
            .in0(N__60163),
            .in1(_gnd_net_),
            .in2(N__53538),
            .in3(N__53454),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net ),
            .ce(N__60016),
            .sr(N__62948));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGH5_LC_23_12_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGH5_LC_23_12_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGH5_LC_23_12_5 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGH5_LC_23_12_5  (
            .in0(N__60589),
            .in1(N__53526),
            .in2(N__53496),
            .in3(N__53481),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGHZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI73BV5_LC_23_12_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI73BV5_LC_23_12_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI73BV5_LC_23_12_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI73BV5_LC_23_12_6  (
            .in0(N__60382),
            .in1(_gnd_net_),
            .in2(N__53475),
            .in3(N__53472),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_16_LC_23_12_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_16_LC_23_12_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_16_LC_23_12_7 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_16_LC_23_12_7  (
            .in0(N__53466),
            .in1(_gnd_net_),
            .in2(N__53457),
            .in3(N__60162),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net ),
            .ce(N__60016),
            .sr(N__62948));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_31_LC_23_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_31_LC_23_13_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_31_LC_23_13_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_31_LC_23_13_0  (
            .in0(_gnd_net_),
            .in1(N__62059),
            .in2(_gnd_net_),
            .in3(N__59602),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_31),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_14_LC_23_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_14_LC_23_13_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_14_LC_23_13_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_14_LC_23_13_1  (
            .in0(N__59603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__58489),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_0_LC_23_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_0_LC_23_13_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_0_LC_23_13_2 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_0_LC_23_13_2  (
            .in0(_gnd_net_),
            .in1(N__59607),
            .in2(_gnd_net_),
            .in3(N__61968),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_15_LC_23_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_15_LC_23_13_3 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_15_LC_23_13_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_15_LC_23_13_3  (
            .in0(N__59604),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57534),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_15),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_24_LC_23_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_24_LC_23_13_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_24_LC_23_13_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_24_LC_23_13_4  (
            .in0(_gnd_net_),
            .in1(N__59600),
            .in2(_gnd_net_),
            .in3(N__61124),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_24),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_16_LC_23_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_16_LC_23_13_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_16_LC_23_13_5 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_16_LC_23_13_5  (
            .in0(N__59605),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57628),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_16),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_28_LC_23_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_28_LC_23_13_6 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_28_LC_23_13_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_28_LC_23_13_6  (
            .in0(_gnd_net_),
            .in1(N__59601),
            .in2(_gnd_net_),
            .in3(N__62357),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_28),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_17_LC_23_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_17_LC_23_13_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_17_LC_23_13_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_17_LC_23_13_7  (
            .in0(N__59606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__57418),
            .lcout(cemf_module_64ch_ctrl_inst1_data_config_17),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65625),
            .ce(N__54118),
            .sr(N__62942));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RL7_LC_23_14_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RL7_LC_23_14_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RL7_LC_23_14_0 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RL7_LC_23_14_0  (
            .in0(N__53992),
            .in1(N__57801),
            .in2(N__54048),
            .in3(N__54576),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIO5CO7_LC_23_14_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIO5CO7_LC_23_14_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIO5CO7_LC_23_14_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIO5CO7_LC_23_14_1  (
            .in0(_gnd_net_),
            .in1(N__53719),
            .in2(N__54030),
            .in3(N__54027),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1_LC_23_14_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1_LC_23_14_2 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1_LC_23_14_2 .LUT_INIT=16'b1100110011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1_LC_23_14_2  (
            .in0(_gnd_net_),
            .in1(N__54021),
            .in2(N__54009),
            .in3(N__55740),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net ),
            .ce(N__55572),
            .sr(N__62937));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RL7_LC_23_14_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RL7_LC_23_14_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RL7_LC_23_14_3 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RL7_LC_23_14_3  (
            .in0(N__53991),
            .in1(N__53788),
            .in2(N__53745),
            .in3(N__53730),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RLZ0Z7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITACO7_LC_23_14_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITACO7_LC_23_14_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITACO7_LC_23_14_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITACO7_LC_23_14_4  (
            .in0(N__53720),
            .in1(_gnd_net_),
            .in2(N__55755),
            .in3(N__55752),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_2_LC_23_14_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_2_LC_23_14_5 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_2_LC_23_14_5 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_2_LC_23_14_5  (
            .in0(N__55741),
            .in1(_gnd_net_),
            .in2(N__55596),
            .in3(N__55593),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net ),
            .ce(N__55572),
            .sr(N__62937));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIG4FN1_LC_23_14_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIG4FN1_LC_23_14_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIG4FN1_LC_23_14_6 .LUT_INIT=16'b1011000010111011;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIG4FN1_LC_23_14_6  (
            .in0(N__55452),
            .in1(N__54634),
            .in2(N__55192),
            .in3(N__54598),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3AQL2_LC_23_14_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3AQL2_LC_23_14_7 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3AQL2_LC_23_14_7 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3AQL2_LC_23_14_7  (
            .in0(N__55054),
            .in1(N__54825),
            .in2(N__54638),
            .in3(N__54599),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_26_LC_23_15_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_26_LC_23_15_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_26_LC_23_15_7 .LUT_INIT=16'b0001000000110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_26_LC_23_15_7  (
            .in0(N__54570),
            .in1(N__54558),
            .in2(N__54546),
            .in3(N__64266),
            .lcout(I2C_top_level_inst1_s_data_oreg_26),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65651),
            .ce(N__54494),
            .sr(N__65010));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIBPUN4_3_LC_23_16_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIBPUN4_3_LC_23_16_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIBPUN4_3_LC_23_16_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIBPUN4_3_LC_23_16_1  (
            .in0(N__54423),
            .in1(N__54380),
            .in2(_gnd_net_),
            .in3(N__54344),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_230 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_230_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_1_LC_23_16_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_1_LC_23_16_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_1_LC_23_16_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_1_LC_23_16_2  (
            .in0(N__56145),
            .in1(N__54258),
            .in2(N__54240),
            .in3(N__56727),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_3_LC_23_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_3_LC_23_16_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_3_LC_23_16_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_3_LC_23_16_3  (
            .in0(N__56728),
            .in1(N__56146),
            .in2(N__56040),
            .in3(N__56070),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_2_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_8_LC_23_16_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_8_LC_23_16_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_8_LC_23_16_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_8_LC_23_16_4  (
            .in0(N__56144),
            .in1(N__56069),
            .in2(_gnd_net_),
            .in3(N__56036),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_4_LC_23_16_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_4_LC_23_16_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_4_LC_23_16_5 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_4_LC_23_16_5  (
            .in0(_gnd_net_),
            .in1(N__62402),
            .in2(N__56013),
            .in3(N__66174),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_365_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_4_LC_23_16_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_4_LC_23_16_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_4_LC_23_16_6 .LUT_INIT=16'b1111010111010101;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_4_LC_23_16_6  (
            .in0(N__56010),
            .in1(N__55869),
            .in2(N__55998),
            .in3(N__55800),
            .lcout(I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65663),
            .ce(),
            .sr(N__65001));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQQ5F_13_LC_23_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQQ5F_13_LC_23_17_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQQ5F_13_LC_23_17_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQQ5F_13_LC_23_17_0  (
            .in0(N__56248),
            .in1(N__64705),
            .in2(N__56353),
            .in3(N__56560),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_4_0_a2_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI4NN21_13_LC_23_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI4NN21_13_LC_23_17_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI4NN21_13_LC_23_17_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI4NN21_13_LC_23_17_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__55995),
            .in3(N__64496),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_676_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIFO0G5_7_LC_23_17_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIFO0G5_7_LC_23_17_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIFO0G5_7_LC_23_17_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIFO0G5_7_LC_23_17_2  (
            .in0(N__55761),
            .in1(N__55767),
            .in2(N__55992),
            .in3(N__55875),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_address ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNISM8F1_3_LC_23_17_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNISM8F1_3_LC_23_17_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNISM8F1_3_LC_23_17_3 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNISM8F1_3_LC_23_17_3  (
            .in0(N__55960),
            .in1(N__56336),
            .in2(N__55944),
            .in3(N__55928),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI05EA2_7_LC_23_17_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI05EA2_7_LC_23_17_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI05EA2_7_LC_23_17_5 .LUT_INIT=16'b0000101000101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI05EA2_7_LC_23_17_5  (
            .in0(N__64704),
            .in1(N__55863),
            .in2(N__57291),
            .in3(N__55795),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1565_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF5IJ_13_LC_23_17_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF5IJ_13_LC_23_17_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF5IJ_13_LC_23_17_6 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF5IJ_13_LC_23_17_6  (
            .in0(_gnd_net_),
            .in1(N__56247),
            .in2(_gnd_net_),
            .in3(N__66244),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_16_LC_23_17_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_16_LC_23_17_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_16_LC_23_17_7 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_16_LC_23_17_7  (
            .in0(_gnd_net_),
            .in1(N__56660),
            .in2(N__56364),
            .in3(N__57208),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_7_0_LC_23_18_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_7_0_LC_23_18_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_7_0_LC_23_18_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_7_0_LC_23_18_0  (
            .in0(N__65897),
            .in1(N__64706),
            .in2(N__57015),
            .in3(N__56350),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_0_LC_23_18_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_0_LC_23_18_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_0_LC_23_18_1 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_0_LC_23_18_1  (
            .in0(N__64707),
            .in1(N__62472),
            .in2(_gnd_net_),
            .in3(N__56351),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_0_LC_23_18_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_0_LC_23_18_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_0_LC_23_18_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_0_LC_23_18_3  (
            .in0(N__66290),
            .in1(N__64802),
            .in2(_gnd_net_),
            .in3(N__64407),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_0_LC_23_18_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_0_LC_23_18_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_0_LC_23_18_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_0_LC_23_18_4  (
            .in0(N__56748),
            .in1(N__56853),
            .in2(N__56283),
            .in3(N__56280),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_11_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_0_LC_23_18_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_0_LC_23_18_5 .SEQ_MODE=4'b1011;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_0_LC_23_18_5 .LUT_INIT=16'b0100110011001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_0_LC_23_18_5  (
            .in0(N__56274),
            .in1(N__56262),
            .in2(N__56253),
            .in3(N__57132),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65689),
            .ce(),
            .sr(N__65014));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASHJ_14_LC_23_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASHJ_14_LC_23_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASHJ_14_LC_23_18_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASHJ_14_LC_23_18_6  (
            .in0(N__64406),
            .in1(N__56700),
            .in2(N__57216),
            .in3(N__56441),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_691 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_23_LC_23_19_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_23_LC_23_19_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_23_LC_23_19_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_23_LC_23_19_0  (
            .in0(N__66251),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__56249),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_23_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_23_LC_23_19_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_23_LC_23_19_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_23_LC_23_19_1 .LUT_INIT=16'b1010101110101111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_23_LC_23_19_1  (
            .in0(N__66166),
            .in1(N__56180),
            .in2(N__56154),
            .in3(N__56559),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAAHD_16_LC_23_19_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAAHD_16_LC_23_19_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAAHD_16_LC_23_19_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAAHD_16_LC_23_19_2  (
            .in0(N__56649),
            .in1(N__64457),
            .in2(_gnd_net_),
            .in3(N__57736),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_288 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_288_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9QGJ_23_LC_23_19_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9QGJ_23_LC_23_19_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9QGJ_23_LC_23_19_3 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9QGJ_23_LC_23_19_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__56742),
            .in3(N__56701),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_231 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_23_LC_23_19_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_23_LC_23_19_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_23_LC_23_19_4 .LUT_INIT=16'b0011001110110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_23_LC_23_19_4  (
            .in0(N__57012),
            .in1(N__56739),
            .in2(N__66449),
            .in3(N__66692),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65704),
            .ce(),
            .sr(N__65022));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_16_LC_23_19_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_16_LC_23_19_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_16_LC_23_19_5 .LUT_INIT=16'b0011000100000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_16_LC_23_19_5  (
            .in0(N__66167),
            .in1(N__56670),
            .in2(N__57227),
            .in3(N__56627),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65704),
            .ce(),
            .sr(N__65022));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_1_LC_23_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_1_LC_23_19_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_1_LC_23_19_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_1_LC_23_19_6  (
            .in0(N__56650),
            .in1(_gnd_net_),
            .in2(N__56631),
            .in3(N__66168),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65704),
            .ce(),
            .sr(N__65022));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_3_LC_23_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_3_LC_23_19_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_3_LC_23_19_7 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_3_LC_23_19_7  (
            .in0(N__64458),
            .in1(N__56516),
            .in2(N__56493),
            .in3(N__56468),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65704),
            .ce(),
            .sr(N__65022));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI046R_4_LC_23_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI046R_4_LC_23_20_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI046R_4_LC_23_20_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI046R_4_LC_23_20_0  (
            .in0(N__56442),
            .in1(N__56908),
            .in2(N__56844),
            .in3(N__56946),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.un30_i_a2_9_a2_4_a2_0_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISICG1_25_LC_23_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISICG1_25_LC_23_20_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISICG1_25_LC_23_20_1 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISICG1_25_LC_23_20_1  (
            .in0(N__56994),
            .in1(N__57056),
            .in2(N__56379),
            .in3(N__64686),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1446 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1446_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPVAM1_12_LC_23_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPVAM1_12_LC_23_20_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPVAM1_12_LC_23_20_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPVAM1_12_LC_23_20_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57060),
            .in3(N__56885),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_245 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI59N81_25_LC_23_20_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI59N81_25_LC_23_20_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI59N81_25_LC_23_20_3 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI59N81_25_LC_23_20_3  (
            .in0(N__56993),
            .in1(N__56770),
            .in2(N__57057),
            .in3(N__64685),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIKLID_24_LC_23_20_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIKLID_24_LC_23_20_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIKLID_24_LC_23_20_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIKLID_24_LC_23_20_4  (
            .in0(N__57028),
            .in1(N__66019),
            .in2(_gnd_net_),
            .in3(N__65978),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_232 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_232_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBFN81_25_LC_23_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBFN81_25_LC_23_20_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBFN81_25_LC_23_20_5 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBFN81_25_LC_23_20_5  (
            .in0(N__56995),
            .in1(N__56964),
            .in2(N__56955),
            .in3(N__64687),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ47E3_25_LC_23_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ47E3_25_LC_23_20_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ47E3_25_LC_23_20_6 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ47E3_25_LC_23_20_6  (
            .in0(N__56771),
            .in1(N__57124),
            .in2(N__56952),
            .in3(N__57082),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_0_LC_23_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_0_LC_23_20_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_0_LC_23_20_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_0_LC_23_20_7  (
            .in0(N__56947),
            .in1(N__56909),
            .in2(N__66333),
            .in3(N__56886),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_0_LC_23_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_0_LC_23_21_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_0_LC_23_21_0 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_0_LC_23_21_0  (
            .in0(N__57255),
            .in1(N__57066),
            .in2(N__56757),
            .in3(N__57300),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65730),
            .ce(),
            .sr(N__65025));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_8_0_LC_23_21_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_8_0_LC_23_21_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_8_0_LC_23_21_1 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_8_0_LC_23_21_1  (
            .in0(N__66779),
            .in1(N__56843),
            .in2(N__64801),
            .in3(N__56829),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_0_LC_23_21_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_0_LC_23_21_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_0_LC_23_21_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_0_LC_23_21_2  (
            .in0(N__56787),
            .in1(N__57146),
            .in2(N__56778),
            .in3(N__56775),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_212 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_0_LC_23_21_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_0_LC_23_21_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_0_LC_23_21_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_0_LC_23_21_3  (
            .in0(N__66780),
            .in1(_gnd_net_),
            .in2(N__57147),
            .in3(N__65800),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_211 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_2_LC_23_21_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_2_LC_23_21_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_2_LC_23_21_4 .LUT_INIT=16'b1100010011110111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_2_LC_23_21_4  (
            .in0(N__65819),
            .in1(N__66493),
            .in2(N__65807),
            .in3(N__57744),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1653_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_2_LC_23_21_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_2_LC_23_21_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_2_LC_23_21_5 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_2_LC_23_21_5  (
            .in0(N__57753),
            .in1(N__66675),
            .in2(N__57294),
            .in3(N__66699),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65730),
            .ce(),
            .sr(N__65025));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_0_LC_23_21_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_0_LC_23_21_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_0_LC_23_21_6 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_0_LC_23_21_6  (
            .in0(N__66548),
            .in1(N__66653),
            .in2(_gnd_net_),
            .in3(N__66492),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_0_LC_23_22_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_0_LC_23_22_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_0_LC_23_22_0 .LUT_INIT=16'b0000100000001010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_0_LC_23_22_0  (
            .in0(N__66851),
            .in1(N__66674),
            .in2(N__57267),
            .in3(N__66559),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9PI7_14_LC_23_22_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9PI7_14_LC_23_22_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9PI7_14_LC_23_22_1 .LUT_INIT=16'b0001000100010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9PI7_14_LC_23_22_1  (
            .in0(N__57223),
            .in1(N__64425),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNI6FAA_0_LC_23_22_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNI6FAA_0_LC_23_22_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNI6FAA_0_LC_23_22_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNI6FAA_0_LC_23_22_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__57150),
            .in3(N__66497),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_239 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_239_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_0_LC_23_22_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_0_LC_23_22_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_0_LC_23_22_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_0_LC_23_22_3  (
            .in0(N__66788),
            .in1(N__66411),
            .in2(N__57135),
            .in3(N__66378),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_0_LC_23_22_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_0_LC_23_22_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_0_LC_23_22_4 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_0_LC_23_22_4  (
            .in0(N__57131),
            .in1(N__57705),
            .in2(N__57093),
            .in3(N__57090),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_2_LC_23_22_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_2_LC_23_22_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_2_LC_23_22_5 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_2_LC_23_22_5  (
            .in0(N__66673),
            .in1(N__66431),
            .in2(_gnd_net_),
            .in3(N__65783),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1776 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNINS3G1_8_LC_23_22_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNINS3G1_8_LC_23_22_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNINS3G1_8_LC_23_22_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNINS3G1_8_LC_23_22_6  (
            .in0(N__66410),
            .in1(N__66377),
            .in2(_gnd_net_),
            .in3(N__66787),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_5_0_LC_23_22_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_5_0_LC_23_22_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_5_0_LC_23_22_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_5_0_LC_23_22_7  (
            .in0(N__66498),
            .in1(N__66850),
            .in2(N__57747),
            .in3(N__57743),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_209 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_0_LC_23_23_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_0_LC_23_23_0 .SEQ_MODE=4'b1000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_0_LC_23_23_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_0_LC_23_23_0  (
            .in0(N__57686),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65748),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16_LC_24_10_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16_LC_24_10_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16_LC_24_10_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16_LC_24_10_0  (
            .in0(N__63341),
            .in1(N__57435),
            .in2(_gnd_net_),
            .in3(N__57620),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net ),
            .ce(N__63030),
            .sr(N__62959));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_15_LC_24_10_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_15_LC_24_10_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_15_LC_24_10_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_15_LC_24_10_1  (
            .in0(N__58386),
            .in1(N__63342),
            .in2(_gnd_net_),
            .in3(N__57496),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net ),
            .ce(N__63030),
            .sr(N__62959));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_17_LC_24_10_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_17_LC_24_10_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_17_LC_24_10_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_17_LC_24_10_7  (
            .in0(N__57429),
            .in1(N__63343),
            .in2(_gnd_net_),
            .in3(N__57419),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net ),
            .ce(N__63030),
            .sr(N__62959));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_19_LC_24_11_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_19_LC_24_11_0 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_19_LC_24_11_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_19_LC_24_11_0  (
            .in0(N__59652),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61640),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_19),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65613),
            .ce(N__58884),
            .sr(N__62957));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_29_LC_24_11_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_29_LC_24_11_1 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_29_LC_24_11_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_29_LC_24_11_1  (
            .in0(_gnd_net_),
            .in1(N__59651),
            .in2(_gnd_net_),
            .in3(N__62260),
            .lcout(cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_29),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65613),
            .ce(N__58884),
            .sr(N__62957));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_0_LC_24_11_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_0_LC_24_11_2 .SEQ_MODE=4'b1011;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_0_LC_24_11_2 .LUT_INIT=16'b0100010001000100;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_0_LC_24_11_2  (
            .in0(N__59653),
            .in1(N__61959),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(cemf_module_64ch_ctrl_inst1_data_coarseovf_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65613),
            .ce(N__58884),
            .sr(N__62957));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10_LC_24_12_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10_LC_24_12_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10_LC_24_12_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10_LC_24_12_0  (
            .in0(N__58818),
            .in1(N__63353),
            .in2(_gnd_net_),
            .in3(N__58795),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ),
            .ce(N__63025),
            .sr(N__62953));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_11_LC_24_12_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_11_LC_24_12_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_11_LC_24_12_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_11_LC_24_12_1  (
            .in0(N__63352),
            .in1(N__58707),
            .in2(_gnd_net_),
            .in3(N__58684),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ),
            .ce(N__63025),
            .sr(N__62953));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_12_LC_24_12_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_12_LC_24_12_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_12_LC_24_12_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_12_LC_24_12_2  (
            .in0(N__58602),
            .in1(N__63354),
            .in2(_gnd_net_),
            .in3(N__58592),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ),
            .ce(N__63025),
            .sr(N__62953));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_14_LC_24_12_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_14_LC_24_12_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_14_LC_24_12_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_14_LC_24_12_4  (
            .in0(N__58263),
            .in1(N__63355),
            .in2(_gnd_net_),
            .in3(N__58473),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ),
            .ce(N__63025),
            .sr(N__62953));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_13_LC_24_12_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_13_LC_24_12_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_13_LC_24_12_7 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_13_LC_24_12_7  (
            .in0(N__58348),
            .in1(_gnd_net_),
            .in2(N__63376),
            .in3(N__58269),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net ),
            .ce(N__63025),
            .sr(N__62953));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIMEB92_17_LC_24_13_0 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIMEB92_17_LC_24_13_0 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIMEB92_17_LC_24_13_0 .LUT_INIT=16'b1000101011001111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIMEB92_17_LC_24_13_0  (
            .in0(N__57987),
            .in1(N__58180),
            .in2(N__58257),
            .in3(N__58211),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOGB92_17_LC_24_13_1 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOGB92_17_LC_24_13_1 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOGB92_17_LC_24_13_1 .LUT_INIT=16'b1000110010101111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOGB92_17_LC_24_13_1  (
            .in0(N__58181),
            .in1(N__57988),
            .in2(N__57833),
            .in3(N__57799),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2Q5_LC_24_13_2 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2Q5_LC_24_13_2 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2Q5_LC_24_13_2 .LUT_INIT=16'b0100111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2Q5_LC_24_13_2  (
            .in0(N__60616),
            .in1(N__60714),
            .in2(N__60678),
            .in3(N__60675),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIP8T76_LC_24_13_3 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIP8T76_LC_24_13_3 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIP8T76_LC_24_13_3 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIP8T76_LC_24_13_3  (
            .in0(_gnd_net_),
            .in1(N__60387),
            .in2(N__60669),
            .in3(N__60666),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1_LC_24_13_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1_LC_24_13_4 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1_LC_24_13_4 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1_LC_24_13_4  (
            .in0(N__60205),
            .in1(_gnd_net_),
            .in2(N__60660),
            .in3(N__60030),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net ),
            .ce(N__60024),
            .sr(N__62949));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2Q5_LC_24_13_5 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2Q5_LC_24_13_5 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2Q5_LC_24_13_5 .LUT_INIT=16'b0010111111111111;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2Q5_LC_24_13_5  (
            .in0(N__60640),
            .in1(N__60615),
            .in2(N__60411),
            .in3(N__60393),
            .lcout(),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2QZ0Z5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIK3T76_LC_24_13_6 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIK3T76_LC_24_13_6 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIK3T76_LC_24_13_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIK3T76_LC_24_13_6  (
            .in0(N__60386),
            .in1(_gnd_net_),
            .in2(N__60219),
            .in3(N__60216),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0 ),
            .ltout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_0_LC_24_13_7 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_0_LC_24_13_7 .SEQ_MODE=4'b1010;
    defparam \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_0_LC_24_13_7 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_0_LC_24_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__60210),
            .in3(N__60204),
            .lcout(\cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net ),
            .ce(N__60024),
            .sr(N__62949));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18_LC_24_14_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18_LC_24_14_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18_LC_24_14_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18_LC_24_14_0  (
            .in0(N__59863),
            .in1(N__59763),
            .in2(_gnd_net_),
            .in3(N__63348),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_18 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_19_LC_24_14_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_19_LC_24_14_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_19_LC_24_14_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_19_LC_24_14_1  (
            .in0(N__63344),
            .in1(N__59754),
            .in2(_gnd_net_),
            .in3(N__61647),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_20_LC_24_14_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_20_LC_24_14_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_20_LC_24_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_20_LC_24_14_2  (
            .in0(N__61551),
            .in1(N__61461),
            .in2(_gnd_net_),
            .in3(N__63349),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_21_LC_24_14_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_21_LC_24_14_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_21_LC_24_14_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_21_LC_24_14_3  (
            .in0(N__63345),
            .in1(N__61455),
            .in2(_gnd_net_),
            .in3(N__61447),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_21 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_22_LC_24_14_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_22_LC_24_14_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_22_LC_24_14_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_22_LC_24_14_4  (
            .in0(N__61362),
            .in1(N__63350),
            .in2(_gnd_net_),
            .in3(N__61355),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_22 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_23_LC_24_14_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_23_LC_24_14_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_23_LC_24_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_23_LC_24_14_5  (
            .in0(N__63346),
            .in1(N__61260),
            .in2(_gnd_net_),
            .in3(N__61229),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_24_LC_24_14_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_24_LC_24_14_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_24_LC_24_14_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_24_LC_24_14_6  (
            .in0(N__61137),
            .in1(N__63351),
            .in2(_gnd_net_),
            .in3(N__61130),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_24 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_25_LC_24_14_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_25_LC_24_14_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_25_LC_24_14_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_25_LC_24_14_7  (
            .in0(N__63347),
            .in1(N__61026),
            .in2(_gnd_net_),
            .in3(N__61000),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_25 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net ),
            .ce(N__63003),
            .sr(N__62943));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26_LC_24_15_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26_LC_24_15_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26_LC_24_15_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26_LC_24_15_0  (
            .in0(N__60927),
            .in1(N__63298),
            .in2(_gnd_net_),
            .in3(N__60849),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_26 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_27_LC_24_15_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_27_LC_24_15_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_27_LC_24_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_27_LC_24_15_1  (
            .in0(N__63295),
            .in1(N__60822),
            .in2(_gnd_net_),
            .in3(N__60798),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_27 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_28_LC_24_15_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_28_LC_24_15_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_28_LC_24_15_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_28_LC_24_15_2  (
            .in0(N__62382),
            .in1(N__63299),
            .in2(_gnd_net_),
            .in3(N__62368),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_29_LC_24_15_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_29_LC_24_15_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_29_LC_24_15_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_29_LC_24_15_3  (
            .in0(N__63296),
            .in1(N__62271),
            .in2(_gnd_net_),
            .in3(N__62261),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_30_LC_24_15_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_30_LC_24_15_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_30_LC_24_15_4 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_30_LC_24_15_4  (
            .in0(N__63300),
            .in1(N__62190),
            .in2(_gnd_net_),
            .in3(N__62169),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_30 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_31_LC_24_15_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_31_LC_24_15_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_31_LC_24_15_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_31_LC_24_15_5  (
            .in0(N__63297),
            .in1(N__62079),
            .in2(_gnd_net_),
            .in3(N__62071),
            .lcout(\I2C_top_level_inst1.s_sda_o_reg ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_i_LC_24_15_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_i_LC_24_15_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_i_LC_24_15_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_i_LC_24_15_6  (
            .in0(_gnd_net_),
            .in1(N__63293),
            .in2(_gnd_net_),
            .in3(N__62421),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_0_LC_24_15_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_0_LC_24_15_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_0_LC_24_15_7 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_0_LC_24_15_7  (
            .in0(N__63294),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__61970),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net ),
            .ce(N__63002),
            .sr(N__62938));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1_LC_24_16_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1_LC_24_16_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1_LC_24_16_0 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1_LC_24_16_0  (
            .in0(N__61878),
            .in1(N__63381),
            .in2(_gnd_net_),
            .in3(N__61872),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_2_LC_24_16_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_2_LC_24_16_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_2_LC_24_16_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_2_LC_24_16_1  (
            .in0(N__63377),
            .in1(N__61752),
            .in2(_gnd_net_),
            .in3(N__61746),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_3_LC_24_16_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_3_LC_24_16_2 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_3_LC_24_16_2 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_3_LC_24_16_2  (
            .in0(N__63951),
            .in1(N__63382),
            .in2(_gnd_net_),
            .in3(N__63944),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_4_LC_24_16_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_4_LC_24_16_3 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_4_LC_24_16_3 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_4_LC_24_16_3  (
            .in0(N__63378),
            .in1(N__63837),
            .in2(_gnd_net_),
            .in3(N__63826),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_5_LC_24_16_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_5_LC_24_16_4 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_5_LC_24_16_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_5_LC_24_16_4  (
            .in0(N__63708),
            .in1(N__63383),
            .in2(_gnd_net_),
            .in3(N__63701),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_6_LC_24_16_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_6_LC_24_16_5 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_6_LC_24_16_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_6_LC_24_16_5  (
            .in0(N__63379),
            .in1(N__63591),
            .in2(_gnd_net_),
            .in3(N__63585),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_7_LC_24_16_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_7_LC_24_16_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_7_LC_24_16_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_7_LC_24_16_6  (
            .in0(N__63489),
            .in1(N__63384),
            .in2(_gnd_net_),
            .in3(N__63477),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_8_LC_24_16_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_8_LC_24_16_7 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_8_LC_24_16_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_8_LC_24_16_7  (
            .in0(N__63380),
            .in1(N__63156),
            .in2(_gnd_net_),
            .in3(N__63118),
            .lcout(\I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net ),
            .ce(N__63015),
            .sr(N__62928));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_LC_24_17_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_LC_24_17_0 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_LC_24_17_0 .LUT_INIT=16'b1000100011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_LC_24_17_0  (
            .in0(N__66866),
            .in1(N__66243),
            .in2(_gnd_net_),
            .in3(N__64605),
            .lcout(I2C_top_level_inst1_s_burst),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65690),
            .ce(),
            .sr(N__65015));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_load_rdata2_LC_24_17_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_load_rdata2_LC_24_17_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_load_rdata2_LC_24_17_1 .LUT_INIT=16'b0010001011111111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_load_rdata2_LC_24_17_1  (
            .in0(N__62420),
            .in1(N__64359),
            .in2(_gnd_net_),
            .in3(N__62480),
            .lcout(\I2C_top_level_inst1.s_load_rdata2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65690),
            .ce(),
            .sr(N__65015));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBMR9_7_LC_24_18_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBMR9_7_LC_24_18_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBMR9_7_LC_24_18_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBMR9_7_LC_24_18_2  (
            .in0(N__64712),
            .in1(N__66593),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_0_LC_24_18_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_0_LC_24_18_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_0_LC_24_18_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_0_LC_24_18_3  (
            .in0(N__64708),
            .in1(N__64629),
            .in2(N__64617),
            .in3(N__66561),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1609_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_0_LC_24_18_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_0_LC_24_18_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_0_LC_24_18_6 .LUT_INIT=16'b1101000111000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_0_LC_24_18_6  (
            .in0(N__64599),
            .in1(N__64551),
            .in2(N__64515),
            .in3(N__64497),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_address_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIG0J7_19_LC_24_19_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIG0J7_19_LC_24_19_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIG0J7_19_LC_24_19_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIG0J7_19_LC_24_19_6  (
            .in0(_gnd_net_),
            .in1(N__65892),
            .in2(_gnd_net_),
            .in3(N__66017),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_295 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_295_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_19_LC_24_19_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_19_LC_24_19_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_19_LC_24_19_7 .LUT_INIT=16'b0011001100100011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_19_LC_24_19_7  (
            .in0(N__65991),
            .in1(N__64323),
            .in2(N__64476),
            .in3(N__64355),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_3_LC_24_20_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_3_LC_24_20_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_3_LC_24_20_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_3_LC_24_20_0  (
            .in0(N__64465),
            .in1(N__65893),
            .in2(N__64437),
            .in3(N__66326),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_RNI63VI_2_LC_24_20_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_RNI63VI_2_LC_24_20_1 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_RNI63VI_2_LC_24_20_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_RNI63VI_2_LC_24_20_1  (
            .in0(N__66327),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__65933),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_19_LC_24_20_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_19_LC_24_20_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_19_LC_24_20_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_19_LC_24_20_2  (
            .in0(N__64344),
            .in1(N__66018),
            .in2(N__65987),
            .in3(N__66328),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_277 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_i2_i_i_o2_i_a2_LC_24_20_4 .C_ON=1'b0;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_i2_i_i_o2_i_a2_LC_24_20_4 .SEQ_MODE=4'b0000;
    defparam \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_i2_i_i_o2_i_a2_LC_24_20_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_i2_i_i_o2_i_a2_LC_24_20_4  (
            .in0(_gnd_net_),
            .in1(N__64299),
            .in2(_gnd_net_),
            .in3(N__64269),
            .lcout(),
            .ltout(N_73_i_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_19_LC_24_20_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_19_LC_24_20_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_19_LC_24_20_5 .LUT_INIT=16'b0100000001000100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_19_LC_24_20_5  (
            .in0(N__66329),
            .in1(N__66291),
            .in2(N__66279),
            .in3(N__66255),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_274_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_19_LC_24_20_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_19_LC_24_20_6 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_19_LC_24_20_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_19_LC_24_20_6  (
            .in0(N__66201),
            .in1(N__65829),
            .in2(N__66195),
            .in3(N__66163),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65731),
            .ce(),
            .sr(N__65026));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_19_LC_24_20_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_19_LC_24_20_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_19_LC_24_20_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_19_LC_24_20_7  (
            .in0(N__65985),
            .in1(N__65934),
            .in2(N__65898),
            .in3(N__65856),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_276 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_1_LC_24_21_0 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_1_LC_24_21_0 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_1_LC_24_21_0 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_1_LC_24_21_0  (
            .in0(N__66553),
            .in1(N__65820),
            .in2(N__65808),
            .in3(N__66687),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1669_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_1_LC_24_21_1 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_1_LC_24_21_1 .SEQ_MODE=4'b1010;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_1_LC_24_21_1 .LUT_INIT=16'b0000100000001100;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_1_LC_24_21_1  (
            .in0(N__65787),
            .in1(N__64809),
            .in2(N__65772),
            .in3(N__64722),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__65740),
            .ce(),
            .sr(N__65027));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_1_LC_24_21_2 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_1_LC_24_21_2 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_1_LC_24_21_2 .LUT_INIT=16'b0000101000001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_1_LC_24_21_2  (
            .in0(N__66853),
            .in1(N__66658),
            .in2(N__64824),
            .in3(N__66496),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_3_LC_24_21_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_3_LC_24_21_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_3_LC_24_21_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_3_LC_24_21_3  (
            .in0(N__64790),
            .in1(N__64721),
            .in2(_gnd_net_),
            .in3(N__66549),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIRCF5_0_LC_24_21_4 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIRCF5_0_LC_24_21_4 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIRCF5_0_LC_24_21_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIRCF5_0_LC_24_21_4  (
            .in0(_gnd_net_),
            .in1(N__66654),
            .in2(_gnd_net_),
            .in3(N__66494),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0 ),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_2_LC_24_21_5 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_2_LC_24_21_5 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_2_LC_24_21_5 .LUT_INIT=16'b1100110011000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_2_LC_24_21_5  (
            .in0(_gnd_net_),
            .in1(N__66852),
            .in2(N__66825),
            .in3(N__66551),
            .lcout(),
            .ltout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_2_LC_24_21_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_2_LC_24_21_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_2_LC_24_21_6 .LUT_INIT=16'b1111000010110000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_2_LC_24_21_6  (
            .in0(N__66552),
            .in1(N__66339),
            .in2(N__66822),
            .in3(N__66798),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_LC_24_21_7 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_LC_24_21_7 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_LC_24_21_7 .LUT_INIT=16'b1111101000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_LC_24_21_7  (
            .in0(N__66495),
            .in1(_gnd_net_),
            .in2(N__66676),
            .in3(N__66550),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNISDF5_0_LC_24_22_3 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNISDF5_0_LC_24_22_3 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNISDF5_0_LC_24_22_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNISDF5_0_LC_24_22_3  (
            .in0(_gnd_net_),
            .in1(N__66555),
            .in2(_gnd_net_),
            .in3(N__66502),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_2_LC_24_22_6 .C_ON=1'b0;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_2_LC_24_22_6 .SEQ_MODE=4'b0000;
    defparam \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_2_LC_24_22_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_2_LC_24_22_6  (
            .in0(_gnd_net_),
            .in1(N__66420),
            .in2(_gnd_net_),
            .in3(N__66384),
            .lcout(\I2C_top_level_inst1.I2C_Interpreter_inst.N_1666_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // cemf_module_64ch_main
