-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Mar 31 2025 15:38:38

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "cemf_module_64ch_main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of cemf_module_64ch_main
entity cemf_module_64ch_main is
port (
    clock : in std_logic;
    start0 : out std_logic;
    s0 : out std_logic;
    intb0 : in std_logic;
    dout1 : out std_logic;
    csb1 : out std_logic;
    sync_50hz : in std_logic;
    sdin1 : in std_logic;
    sda : inout std_logic;
    s1 : out std_logic;
    intb1 : in std_logic;
    dout0 : out std_logic;
    csb0 : out std_logic;
    serial_out_testing : out std_logic;
    sdin0 : in std_logic;
    scl : in std_logic;
    s2 : out std_logic;
    mcu_sclk : out std_logic;
    frame_sync : out std_logic;
    enable_config : out std_logic;
    elec_config_out : out std_logic;
    stop1 : out std_logic;
    s3 : out std_logic;
    rst_n : in std_logic;
    cemf_signal : in std_logic;
    trigger1 : in std_logic;
    stop0 : out std_logic;
    trigger0 : in std_logic;
    stop_fpga2 : out std_logic;
    sclk0 : out std_logic;
    next_sequence : out std_logic;
    start1 : out std_logic;
    sclk1 : out std_logic;
    mcu_data : out std_logic);
end cemf_module_64ch_main;

-- Architecture of cemf_module_64ch_main
-- View name is \INTERFACE\
architecture \INTERFACE\ of cemf_module_64ch_main is

signal \N__67138\ : std_logic;
signal \N__67137\ : std_logic;
signal \N__67136\ : std_logic;
signal \N__67129\ : std_logic;
signal \N__67128\ : std_logic;
signal \N__67127\ : std_logic;
signal \N__67120\ : std_logic;
signal \N__67119\ : std_logic;
signal \N__67118\ : std_logic;
signal \N__67111\ : std_logic;
signal \N__67110\ : std_logic;
signal \N__67109\ : std_logic;
signal \N__67102\ : std_logic;
signal \N__67101\ : std_logic;
signal \N__67100\ : std_logic;
signal \N__67093\ : std_logic;
signal \N__67092\ : std_logic;
signal \N__67091\ : std_logic;
signal \N__67084\ : std_logic;
signal \N__67083\ : std_logic;
signal \N__67082\ : std_logic;
signal \N__67075\ : std_logic;
signal \N__67074\ : std_logic;
signal \N__67073\ : std_logic;
signal \N__67066\ : std_logic;
signal \N__67065\ : std_logic;
signal \N__67064\ : std_logic;
signal \N__67057\ : std_logic;
signal \N__67056\ : std_logic;
signal \N__67055\ : std_logic;
signal \N__67048\ : std_logic;
signal \N__67047\ : std_logic;
signal \N__67046\ : std_logic;
signal \N__67039\ : std_logic;
signal \N__67038\ : std_logic;
signal \N__67037\ : std_logic;
signal \N__67030\ : std_logic;
signal \N__67029\ : std_logic;
signal \N__67028\ : std_logic;
signal \N__67021\ : std_logic;
signal \N__67020\ : std_logic;
signal \N__67019\ : std_logic;
signal \N__67012\ : std_logic;
signal \N__67011\ : std_logic;
signal \N__67010\ : std_logic;
signal \N__67003\ : std_logic;
signal \N__67002\ : std_logic;
signal \N__67001\ : std_logic;
signal \N__66994\ : std_logic;
signal \N__66993\ : std_logic;
signal \N__66992\ : std_logic;
signal \N__66985\ : std_logic;
signal \N__66984\ : std_logic;
signal \N__66983\ : std_logic;
signal \N__66976\ : std_logic;
signal \N__66975\ : std_logic;
signal \N__66974\ : std_logic;
signal \N__66967\ : std_logic;
signal \N__66966\ : std_logic;
signal \N__66965\ : std_logic;
signal \N__66958\ : std_logic;
signal \N__66957\ : std_logic;
signal \N__66956\ : std_logic;
signal \N__66949\ : std_logic;
signal \N__66948\ : std_logic;
signal \N__66947\ : std_logic;
signal \N__66940\ : std_logic;
signal \N__66939\ : std_logic;
signal \N__66938\ : std_logic;
signal \N__66931\ : std_logic;
signal \N__66930\ : std_logic;
signal \N__66929\ : std_logic;
signal \N__66922\ : std_logic;
signal \N__66921\ : std_logic;
signal \N__66920\ : std_logic;
signal \N__66913\ : std_logic;
signal \N__66912\ : std_logic;
signal \N__66911\ : std_logic;
signal \N__66904\ : std_logic;
signal \N__66903\ : std_logic;
signal \N__66902\ : std_logic;
signal \N__66895\ : std_logic;
signal \N__66894\ : std_logic;
signal \N__66893\ : std_logic;
signal \N__66886\ : std_logic;
signal \N__66885\ : std_logic;
signal \N__66884\ : std_logic;
signal \N__66867\ : std_logic;
signal \N__66866\ : std_logic;
signal \N__66863\ : std_logic;
signal \N__66860\ : std_logic;
signal \N__66857\ : std_logic;
signal \N__66854\ : std_logic;
signal \N__66853\ : std_logic;
signal \N__66852\ : std_logic;
signal \N__66851\ : std_logic;
signal \N__66850\ : std_logic;
signal \N__66847\ : std_logic;
signal \N__66844\ : std_logic;
signal \N__66839\ : std_logic;
signal \N__66834\ : std_logic;
signal \N__66825\ : std_logic;
signal \N__66822\ : std_logic;
signal \N__66819\ : std_logic;
signal \N__66816\ : std_logic;
signal \N__66815\ : std_logic;
signal \N__66814\ : std_logic;
signal \N__66813\ : std_logic;
signal \N__66806\ : std_logic;
signal \N__66803\ : std_logic;
signal \N__66800\ : std_logic;
signal \N__66799\ : std_logic;
signal \N__66798\ : std_logic;
signal \N__66795\ : std_logic;
signal \N__66794\ : std_logic;
signal \N__66791\ : std_logic;
signal \N__66790\ : std_logic;
signal \N__66789\ : std_logic;
signal \N__66788\ : std_logic;
signal \N__66787\ : std_logic;
signal \N__66784\ : std_logic;
signal \N__66781\ : std_logic;
signal \N__66780\ : std_logic;
signal \N__66779\ : std_logic;
signal \N__66776\ : std_logic;
signal \N__66773\ : std_logic;
signal \N__66770\ : std_logic;
signal \N__66769\ : std_logic;
signal \N__66764\ : std_logic;
signal \N__66759\ : std_logic;
signal \N__66756\ : std_logic;
signal \N__66755\ : std_logic;
signal \N__66752\ : std_logic;
signal \N__66747\ : std_logic;
signal \N__66744\ : std_logic;
signal \N__66739\ : std_logic;
signal \N__66736\ : std_logic;
signal \N__66731\ : std_logic;
signal \N__66728\ : std_logic;
signal \N__66725\ : std_logic;
signal \N__66720\ : std_logic;
signal \N__66715\ : std_logic;
signal \N__66708\ : std_logic;
signal \N__66699\ : std_logic;
signal \N__66696\ : std_logic;
signal \N__66693\ : std_logic;
signal \N__66692\ : std_logic;
signal \N__66691\ : std_logic;
signal \N__66688\ : std_logic;
signal \N__66687\ : std_logic;
signal \N__66684\ : std_logic;
signal \N__66681\ : std_logic;
signal \N__66680\ : std_logic;
signal \N__66677\ : std_logic;
signal \N__66676\ : std_logic;
signal \N__66675\ : std_logic;
signal \N__66674\ : std_logic;
signal \N__66673\ : std_logic;
signal \N__66670\ : std_logic;
signal \N__66665\ : std_logic;
signal \N__66662\ : std_logic;
signal \N__66659\ : std_logic;
signal \N__66658\ : std_logic;
signal \N__66655\ : std_logic;
signal \N__66654\ : std_logic;
signal \N__66653\ : std_logic;
signal \N__66650\ : std_logic;
signal \N__66645\ : std_logic;
signal \N__66640\ : std_logic;
signal \N__66637\ : std_logic;
signal \N__66634\ : std_logic;
signal \N__66627\ : std_logic;
signal \N__66624\ : std_logic;
signal \N__66609\ : std_logic;
signal \N__66608\ : std_logic;
signal \N__66607\ : std_logic;
signal \N__66604\ : std_logic;
signal \N__66603\ : std_logic;
signal \N__66602\ : std_logic;
signal \N__66599\ : std_logic;
signal \N__66594\ : std_logic;
signal \N__66593\ : std_logic;
signal \N__66590\ : std_logic;
signal \N__66587\ : std_logic;
signal \N__66582\ : std_logic;
signal \N__66579\ : std_logic;
signal \N__66574\ : std_logic;
signal \N__66571\ : std_logic;
signal \N__66568\ : std_logic;
signal \N__66561\ : std_logic;
signal \N__66560\ : std_logic;
signal \N__66559\ : std_logic;
signal \N__66556\ : std_logic;
signal \N__66555\ : std_logic;
signal \N__66554\ : std_logic;
signal \N__66553\ : std_logic;
signal \N__66552\ : std_logic;
signal \N__66551\ : std_logic;
signal \N__66550\ : std_logic;
signal \N__66549\ : std_logic;
signal \N__66548\ : std_logic;
signal \N__66545\ : std_logic;
signal \N__66542\ : std_logic;
signal \N__66539\ : std_logic;
signal \N__66536\ : std_logic;
signal \N__66533\ : std_logic;
signal \N__66522\ : std_logic;
signal \N__66519\ : std_logic;
signal \N__66504\ : std_logic;
signal \N__66503\ : std_logic;
signal \N__66502\ : std_logic;
signal \N__66499\ : std_logic;
signal \N__66498\ : std_logic;
signal \N__66497\ : std_logic;
signal \N__66496\ : std_logic;
signal \N__66495\ : std_logic;
signal \N__66494\ : std_logic;
signal \N__66493\ : std_logic;
signal \N__66492\ : std_logic;
signal \N__66489\ : std_logic;
signal \N__66486\ : std_logic;
signal \N__66483\ : std_logic;
signal \N__66478\ : std_logic;
signal \N__66471\ : std_logic;
signal \N__66466\ : std_logic;
signal \N__66453\ : std_logic;
signal \N__66450\ : std_logic;
signal \N__66449\ : std_logic;
signal \N__66446\ : std_logic;
signal \N__66443\ : std_logic;
signal \N__66440\ : std_logic;
signal \N__66437\ : std_logic;
signal \N__66432\ : std_logic;
signal \N__66431\ : std_logic;
signal \N__66428\ : std_logic;
signal \N__66425\ : std_logic;
signal \N__66420\ : std_logic;
signal \N__66419\ : std_logic;
signal \N__66416\ : std_logic;
signal \N__66413\ : std_logic;
signal \N__66412\ : std_logic;
signal \N__66411\ : std_logic;
signal \N__66410\ : std_logic;
signal \N__66407\ : std_logic;
signal \N__66402\ : std_logic;
signal \N__66397\ : std_logic;
signal \N__66394\ : std_logic;
signal \N__66389\ : std_logic;
signal \N__66384\ : std_logic;
signal \N__66383\ : std_logic;
signal \N__66382\ : std_logic;
signal \N__66379\ : std_logic;
signal \N__66378\ : std_logic;
signal \N__66377\ : std_logic;
signal \N__66376\ : std_logic;
signal \N__66375\ : std_logic;
signal \N__66370\ : std_logic;
signal \N__66367\ : std_logic;
signal \N__66364\ : std_logic;
signal \N__66361\ : std_logic;
signal \N__66356\ : std_logic;
signal \N__66353\ : std_logic;
signal \N__66346\ : std_logic;
signal \N__66339\ : std_logic;
signal \N__66336\ : std_logic;
signal \N__66333\ : std_logic;
signal \N__66330\ : std_logic;
signal \N__66329\ : std_logic;
signal \N__66328\ : std_logic;
signal \N__66327\ : std_logic;
signal \N__66326\ : std_logic;
signal \N__66325\ : std_logic;
signal \N__66324\ : std_logic;
signal \N__66321\ : std_logic;
signal \N__66312\ : std_logic;
signal \N__66309\ : std_logic;
signal \N__66306\ : std_logic;
signal \N__66303\ : std_logic;
signal \N__66300\ : std_logic;
signal \N__66291\ : std_logic;
signal \N__66290\ : std_logic;
signal \N__66287\ : std_logic;
signal \N__66284\ : std_logic;
signal \N__66279\ : std_logic;
signal \N__66276\ : std_logic;
signal \N__66275\ : std_logic;
signal \N__66274\ : std_logic;
signal \N__66273\ : std_logic;
signal \N__66268\ : std_logic;
signal \N__66265\ : std_logic;
signal \N__66264\ : std_logic;
signal \N__66261\ : std_logic;
signal \N__66256\ : std_logic;
signal \N__66255\ : std_logic;
signal \N__66252\ : std_logic;
signal \N__66251\ : std_logic;
signal \N__66248\ : std_logic;
signal \N__66245\ : std_logic;
signal \N__66244\ : std_logic;
signal \N__66243\ : std_logic;
signal \N__66240\ : std_logic;
signal \N__66237\ : std_logic;
signal \N__66234\ : std_logic;
signal \N__66229\ : std_logic;
signal \N__66226\ : std_logic;
signal \N__66223\ : std_logic;
signal \N__66220\ : std_logic;
signal \N__66215\ : std_logic;
signal \N__66210\ : std_logic;
signal \N__66201\ : std_logic;
signal \N__66198\ : std_logic;
signal \N__66195\ : std_logic;
signal \N__66192\ : std_logic;
signal \N__66191\ : std_logic;
signal \N__66188\ : std_logic;
signal \N__66187\ : std_logic;
signal \N__66186\ : std_logic;
signal \N__66185\ : std_logic;
signal \N__66184\ : std_logic;
signal \N__66175\ : std_logic;
signal \N__66174\ : std_logic;
signal \N__66169\ : std_logic;
signal \N__66168\ : std_logic;
signal \N__66167\ : std_logic;
signal \N__66166\ : std_logic;
signal \N__66165\ : std_logic;
signal \N__66164\ : std_logic;
signal \N__66163\ : std_logic;
signal \N__66160\ : std_logic;
signal \N__66157\ : std_logic;
signal \N__66156\ : std_logic;
signal \N__66155\ : std_logic;
signal \N__66154\ : std_logic;
signal \N__66151\ : std_logic;
signal \N__66150\ : std_logic;
signal \N__66143\ : std_logic;
signal \N__66138\ : std_logic;
signal \N__66135\ : std_logic;
signal \N__66130\ : std_logic;
signal \N__66129\ : std_logic;
signal \N__66126\ : std_logic;
signal \N__66125\ : std_logic;
signal \N__66122\ : std_logic;
signal \N__66119\ : std_logic;
signal \N__66118\ : std_logic;
signal \N__66115\ : std_logic;
signal \N__66112\ : std_logic;
signal \N__66111\ : std_logic;
signal \N__66110\ : std_logic;
signal \N__66109\ : std_logic;
signal \N__66106\ : std_logic;
signal \N__66105\ : std_logic;
signal \N__66102\ : std_logic;
signal \N__66099\ : std_logic;
signal \N__66096\ : std_logic;
signal \N__66095\ : std_logic;
signal \N__66094\ : std_logic;
signal \N__66093\ : std_logic;
signal \N__66086\ : std_logic;
signal \N__66079\ : std_logic;
signal \N__66074\ : std_logic;
signal \N__66067\ : std_logic;
signal \N__66064\ : std_logic;
signal \N__66061\ : std_logic;
signal \N__66054\ : std_logic;
signal \N__66051\ : std_logic;
signal \N__66046\ : std_logic;
signal \N__66041\ : std_logic;
signal \N__66038\ : std_logic;
signal \N__66021\ : std_logic;
signal \N__66020\ : std_logic;
signal \N__66019\ : std_logic;
signal \N__66018\ : std_logic;
signal \N__66017\ : std_logic;
signal \N__66012\ : std_logic;
signal \N__66009\ : std_logic;
signal \N__66006\ : std_logic;
signal \N__66003\ : std_logic;
signal \N__65998\ : std_logic;
signal \N__65991\ : std_logic;
signal \N__65988\ : std_logic;
signal \N__65987\ : std_logic;
signal \N__65986\ : std_logic;
signal \N__65985\ : std_logic;
signal \N__65982\ : std_logic;
signal \N__65979\ : std_logic;
signal \N__65978\ : std_logic;
signal \N__65975\ : std_logic;
signal \N__65974\ : std_logic;
signal \N__65971\ : std_logic;
signal \N__65968\ : std_logic;
signal \N__65965\ : std_logic;
signal \N__65962\ : std_logic;
signal \N__65957\ : std_logic;
signal \N__65946\ : std_logic;
signal \N__65945\ : std_logic;
signal \N__65942\ : std_logic;
signal \N__65939\ : std_logic;
signal \N__65934\ : std_logic;
signal \N__65933\ : std_logic;
signal \N__65932\ : std_logic;
signal \N__65927\ : std_logic;
signal \N__65926\ : std_logic;
signal \N__65923\ : std_logic;
signal \N__65920\ : std_logic;
signal \N__65915\ : std_logic;
signal \N__65914\ : std_logic;
signal \N__65909\ : std_logic;
signal \N__65906\ : std_logic;
signal \N__65903\ : std_logic;
signal \N__65898\ : std_logic;
signal \N__65897\ : std_logic;
signal \N__65894\ : std_logic;
signal \N__65893\ : std_logic;
signal \N__65892\ : std_logic;
signal \N__65889\ : std_logic;
signal \N__65884\ : std_logic;
signal \N__65881\ : std_logic;
signal \N__65878\ : std_logic;
signal \N__65873\ : std_logic;
signal \N__65872\ : std_logic;
signal \N__65871\ : std_logic;
signal \N__65866\ : std_logic;
signal \N__65861\ : std_logic;
signal \N__65856\ : std_logic;
signal \N__65853\ : std_logic;
signal \N__65852\ : std_logic;
signal \N__65849\ : std_logic;
signal \N__65848\ : std_logic;
signal \N__65845\ : std_logic;
signal \N__65842\ : std_logic;
signal \N__65839\ : std_logic;
signal \N__65836\ : std_logic;
signal \N__65829\ : std_logic;
signal \N__65826\ : std_logic;
signal \N__65823\ : std_logic;
signal \N__65820\ : std_logic;
signal \N__65819\ : std_logic;
signal \N__65816\ : std_logic;
signal \N__65813\ : std_logic;
signal \N__65808\ : std_logic;
signal \N__65807\ : std_logic;
signal \N__65804\ : std_logic;
signal \N__65801\ : std_logic;
signal \N__65800\ : std_logic;
signal \N__65797\ : std_logic;
signal \N__65792\ : std_logic;
signal \N__65787\ : std_logic;
signal \N__65784\ : std_logic;
signal \N__65783\ : std_logic;
signal \N__65780\ : std_logic;
signal \N__65777\ : std_logic;
signal \N__65772\ : std_logic;
signal \N__65769\ : std_logic;
signal \N__65768\ : std_logic;
signal \N__65767\ : std_logic;
signal \N__65764\ : std_logic;
signal \N__65761\ : std_logic;
signal \N__65758\ : std_logic;
signal \N__65755\ : std_logic;
signal \N__65754\ : std_logic;
signal \N__65753\ : std_logic;
signal \N__65752\ : std_logic;
signal \N__65751\ : std_logic;
signal \N__65750\ : std_logic;
signal \N__65749\ : std_logic;
signal \N__65748\ : std_logic;
signal \N__65747\ : std_logic;
signal \N__65746\ : std_logic;
signal \N__65745\ : std_logic;
signal \N__65744\ : std_logic;
signal \N__65743\ : std_logic;
signal \N__65742\ : std_logic;
signal \N__65741\ : std_logic;
signal \N__65740\ : std_logic;
signal \N__65739\ : std_logic;
signal \N__65738\ : std_logic;
signal \N__65737\ : std_logic;
signal \N__65736\ : std_logic;
signal \N__65735\ : std_logic;
signal \N__65734\ : std_logic;
signal \N__65733\ : std_logic;
signal \N__65732\ : std_logic;
signal \N__65731\ : std_logic;
signal \N__65730\ : std_logic;
signal \N__65729\ : std_logic;
signal \N__65728\ : std_logic;
signal \N__65727\ : std_logic;
signal \N__65726\ : std_logic;
signal \N__65725\ : std_logic;
signal \N__65724\ : std_logic;
signal \N__65723\ : std_logic;
signal \N__65722\ : std_logic;
signal \N__65721\ : std_logic;
signal \N__65720\ : std_logic;
signal \N__65719\ : std_logic;
signal \N__65718\ : std_logic;
signal \N__65717\ : std_logic;
signal \N__65716\ : std_logic;
signal \N__65715\ : std_logic;
signal \N__65714\ : std_logic;
signal \N__65713\ : std_logic;
signal \N__65710\ : std_logic;
signal \N__65707\ : std_logic;
signal \N__65706\ : std_logic;
signal \N__65705\ : std_logic;
signal \N__65704\ : std_logic;
signal \N__65703\ : std_logic;
signal \N__65702\ : std_logic;
signal \N__65701\ : std_logic;
signal \N__65700\ : std_logic;
signal \N__65699\ : std_logic;
signal \N__65698\ : std_logic;
signal \N__65697\ : std_logic;
signal \N__65696\ : std_logic;
signal \N__65695\ : std_logic;
signal \N__65694\ : std_logic;
signal \N__65693\ : std_logic;
signal \N__65692\ : std_logic;
signal \N__65691\ : std_logic;
signal \N__65690\ : std_logic;
signal \N__65689\ : std_logic;
signal \N__65688\ : std_logic;
signal \N__65687\ : std_logic;
signal \N__65686\ : std_logic;
signal \N__65685\ : std_logic;
signal \N__65684\ : std_logic;
signal \N__65683\ : std_logic;
signal \N__65682\ : std_logic;
signal \N__65681\ : std_logic;
signal \N__65680\ : std_logic;
signal \N__65679\ : std_logic;
signal \N__65678\ : std_logic;
signal \N__65677\ : std_logic;
signal \N__65676\ : std_logic;
signal \N__65675\ : std_logic;
signal \N__65674\ : std_logic;
signal \N__65673\ : std_logic;
signal \N__65672\ : std_logic;
signal \N__65671\ : std_logic;
signal \N__65670\ : std_logic;
signal \N__65669\ : std_logic;
signal \N__65668\ : std_logic;
signal \N__65667\ : std_logic;
signal \N__65666\ : std_logic;
signal \N__65665\ : std_logic;
signal \N__65664\ : std_logic;
signal \N__65663\ : std_logic;
signal \N__65662\ : std_logic;
signal \N__65661\ : std_logic;
signal \N__65660\ : std_logic;
signal \N__65659\ : std_logic;
signal \N__65658\ : std_logic;
signal \N__65657\ : std_logic;
signal \N__65656\ : std_logic;
signal \N__65655\ : std_logic;
signal \N__65654\ : std_logic;
signal \N__65653\ : std_logic;
signal \N__65652\ : std_logic;
signal \N__65651\ : std_logic;
signal \N__65650\ : std_logic;
signal \N__65649\ : std_logic;
signal \N__65648\ : std_logic;
signal \N__65647\ : std_logic;
signal \N__65646\ : std_logic;
signal \N__65645\ : std_logic;
signal \N__65644\ : std_logic;
signal \N__65643\ : std_logic;
signal \N__65642\ : std_logic;
signal \N__65641\ : std_logic;
signal \N__65640\ : std_logic;
signal \N__65639\ : std_logic;
signal \N__65638\ : std_logic;
signal \N__65637\ : std_logic;
signal \N__65636\ : std_logic;
signal \N__65635\ : std_logic;
signal \N__65634\ : std_logic;
signal \N__65633\ : std_logic;
signal \N__65632\ : std_logic;
signal \N__65631\ : std_logic;
signal \N__65630\ : std_logic;
signal \N__65629\ : std_logic;
signal \N__65628\ : std_logic;
signal \N__65627\ : std_logic;
signal \N__65626\ : std_logic;
signal \N__65625\ : std_logic;
signal \N__65624\ : std_logic;
signal \N__65623\ : std_logic;
signal \N__65622\ : std_logic;
signal \N__65621\ : std_logic;
signal \N__65620\ : std_logic;
signal \N__65619\ : std_logic;
signal \N__65618\ : std_logic;
signal \N__65617\ : std_logic;
signal \N__65616\ : std_logic;
signal \N__65615\ : std_logic;
signal \N__65614\ : std_logic;
signal \N__65613\ : std_logic;
signal \N__65612\ : std_logic;
signal \N__65611\ : std_logic;
signal \N__65610\ : std_logic;
signal \N__65609\ : std_logic;
signal \N__65608\ : std_logic;
signal \N__65607\ : std_logic;
signal \N__65606\ : std_logic;
signal \N__65605\ : std_logic;
signal \N__65604\ : std_logic;
signal \N__65603\ : std_logic;
signal \N__65602\ : std_logic;
signal \N__65601\ : std_logic;
signal \N__65600\ : std_logic;
signal \N__65599\ : std_logic;
signal \N__65598\ : std_logic;
signal \N__65597\ : std_logic;
signal \N__65596\ : std_logic;
signal \N__65595\ : std_logic;
signal \N__65594\ : std_logic;
signal \N__65593\ : std_logic;
signal \N__65592\ : std_logic;
signal \N__65591\ : std_logic;
signal \N__65590\ : std_logic;
signal \N__65589\ : std_logic;
signal \N__65588\ : std_logic;
signal \N__65587\ : std_logic;
signal \N__65586\ : std_logic;
signal \N__65585\ : std_logic;
signal \N__65584\ : std_logic;
signal \N__65583\ : std_logic;
signal \N__65582\ : std_logic;
signal \N__65581\ : std_logic;
signal \N__65580\ : std_logic;
signal \N__65579\ : std_logic;
signal \N__65578\ : std_logic;
signal \N__65577\ : std_logic;
signal \N__65576\ : std_logic;
signal \N__65575\ : std_logic;
signal \N__65574\ : std_logic;
signal \N__65573\ : std_logic;
signal \N__65572\ : std_logic;
signal \N__65571\ : std_logic;
signal \N__65570\ : std_logic;
signal \N__65569\ : std_logic;
signal \N__65568\ : std_logic;
signal \N__65567\ : std_logic;
signal \N__65566\ : std_logic;
signal \N__65565\ : std_logic;
signal \N__65564\ : std_logic;
signal \N__65563\ : std_logic;
signal \N__65562\ : std_logic;
signal \N__65561\ : std_logic;
signal \N__65560\ : std_logic;
signal \N__65559\ : std_logic;
signal \N__65558\ : std_logic;
signal \N__65557\ : std_logic;
signal \N__65556\ : std_logic;
signal \N__65555\ : std_logic;
signal \N__65554\ : std_logic;
signal \N__65553\ : std_logic;
signal \N__65552\ : std_logic;
signal \N__65551\ : std_logic;
signal \N__65550\ : std_logic;
signal \N__65549\ : std_logic;
signal \N__65548\ : std_logic;
signal \N__65547\ : std_logic;
signal \N__65546\ : std_logic;
signal \N__65545\ : std_logic;
signal \N__65544\ : std_logic;
signal \N__65543\ : std_logic;
signal \N__65542\ : std_logic;
signal \N__65541\ : std_logic;
signal \N__65540\ : std_logic;
signal \N__65539\ : std_logic;
signal \N__65538\ : std_logic;
signal \N__65537\ : std_logic;
signal \N__65536\ : std_logic;
signal \N__65535\ : std_logic;
signal \N__65534\ : std_logic;
signal \N__65533\ : std_logic;
signal \N__65532\ : std_logic;
signal \N__65531\ : std_logic;
signal \N__65530\ : std_logic;
signal \N__65529\ : std_logic;
signal \N__65528\ : std_logic;
signal \N__65527\ : std_logic;
signal \N__65526\ : std_logic;
signal \N__65525\ : std_logic;
signal \N__65524\ : std_logic;
signal \N__65523\ : std_logic;
signal \N__65522\ : std_logic;
signal \N__65521\ : std_logic;
signal \N__65520\ : std_logic;
signal \N__65519\ : std_logic;
signal \N__65518\ : std_logic;
signal \N__65517\ : std_logic;
signal \N__65516\ : std_logic;
signal \N__65515\ : std_logic;
signal \N__65514\ : std_logic;
signal \N__65513\ : std_logic;
signal \N__65034\ : std_logic;
signal \N__65031\ : std_logic;
signal \N__65028\ : std_logic;
signal \N__65027\ : std_logic;
signal \N__65026\ : std_logic;
signal \N__65025\ : std_logic;
signal \N__65024\ : std_logic;
signal \N__65023\ : std_logic;
signal \N__65022\ : std_logic;
signal \N__65021\ : std_logic;
signal \N__65020\ : std_logic;
signal \N__65019\ : std_logic;
signal \N__65018\ : std_logic;
signal \N__65017\ : std_logic;
signal \N__65016\ : std_logic;
signal \N__65015\ : std_logic;
signal \N__65014\ : std_logic;
signal \N__65013\ : std_logic;
signal \N__65012\ : std_logic;
signal \N__65011\ : std_logic;
signal \N__65010\ : std_logic;
signal \N__65009\ : std_logic;
signal \N__65008\ : std_logic;
signal \N__65007\ : std_logic;
signal \N__65006\ : std_logic;
signal \N__65005\ : std_logic;
signal \N__65004\ : std_logic;
signal \N__65003\ : std_logic;
signal \N__65002\ : std_logic;
signal \N__65001\ : std_logic;
signal \N__65000\ : std_logic;
signal \N__64999\ : std_logic;
signal \N__64998\ : std_logic;
signal \N__64997\ : std_logic;
signal \N__64996\ : std_logic;
signal \N__64995\ : std_logic;
signal \N__64994\ : std_logic;
signal \N__64993\ : std_logic;
signal \N__64992\ : std_logic;
signal \N__64991\ : std_logic;
signal \N__64990\ : std_logic;
signal \N__64989\ : std_logic;
signal \N__64988\ : std_logic;
signal \N__64987\ : std_logic;
signal \N__64986\ : std_logic;
signal \N__64985\ : std_logic;
signal \N__64984\ : std_logic;
signal \N__64983\ : std_logic;
signal \N__64982\ : std_logic;
signal \N__64981\ : std_logic;
signal \N__64980\ : std_logic;
signal \N__64979\ : std_logic;
signal \N__64978\ : std_logic;
signal \N__64977\ : std_logic;
signal \N__64976\ : std_logic;
signal \N__64975\ : std_logic;
signal \N__64974\ : std_logic;
signal \N__64973\ : std_logic;
signal \N__64972\ : std_logic;
signal \N__64971\ : std_logic;
signal \N__64970\ : std_logic;
signal \N__64969\ : std_logic;
signal \N__64968\ : std_logic;
signal \N__64967\ : std_logic;
signal \N__64966\ : std_logic;
signal \N__64965\ : std_logic;
signal \N__64964\ : std_logic;
signal \N__64963\ : std_logic;
signal \N__64830\ : std_logic;
signal \N__64827\ : std_logic;
signal \N__64824\ : std_logic;
signal \N__64821\ : std_logic;
signal \N__64818\ : std_logic;
signal \N__64815\ : std_logic;
signal \N__64812\ : std_logic;
signal \N__64809\ : std_logic;
signal \N__64806\ : std_logic;
signal \N__64803\ : std_logic;
signal \N__64802\ : std_logic;
signal \N__64801\ : std_logic;
signal \N__64798\ : std_logic;
signal \N__64795\ : std_logic;
signal \N__64794\ : std_logic;
signal \N__64791\ : std_logic;
signal \N__64790\ : std_logic;
signal \N__64789\ : std_logic;
signal \N__64788\ : std_logic;
signal \N__64787\ : std_logic;
signal \N__64784\ : std_logic;
signal \N__64781\ : std_logic;
signal \N__64778\ : std_logic;
signal \N__64775\ : std_logic;
signal \N__64772\ : std_logic;
signal \N__64769\ : std_logic;
signal \N__64766\ : std_logic;
signal \N__64763\ : std_logic;
signal \N__64756\ : std_logic;
signal \N__64751\ : std_logic;
signal \N__64748\ : std_logic;
signal \N__64737\ : std_logic;
signal \N__64734\ : std_logic;
signal \N__64731\ : std_logic;
signal \N__64728\ : std_logic;
signal \N__64725\ : std_logic;
signal \N__64722\ : std_logic;
signal \N__64721\ : std_logic;
signal \N__64716\ : std_logic;
signal \N__64713\ : std_logic;
signal \N__64712\ : std_logic;
signal \N__64709\ : std_logic;
signal \N__64708\ : std_logic;
signal \N__64707\ : std_logic;
signal \N__64706\ : std_logic;
signal \N__64705\ : std_logic;
signal \N__64704\ : std_logic;
signal \N__64701\ : std_logic;
signal \N__64698\ : std_logic;
signal \N__64697\ : std_logic;
signal \N__64696\ : std_logic;
signal \N__64693\ : std_logic;
signal \N__64688\ : std_logic;
signal \N__64687\ : std_logic;
signal \N__64686\ : std_logic;
signal \N__64685\ : std_logic;
signal \N__64680\ : std_logic;
signal \N__64679\ : std_logic;
signal \N__64674\ : std_logic;
signal \N__64669\ : std_logic;
signal \N__64664\ : std_logic;
signal \N__64657\ : std_logic;
signal \N__64654\ : std_logic;
signal \N__64651\ : std_logic;
signal \N__64648\ : std_logic;
signal \N__64641\ : std_logic;
signal \N__64638\ : std_logic;
signal \N__64629\ : std_logic;
signal \N__64626\ : std_logic;
signal \N__64623\ : std_logic;
signal \N__64620\ : std_logic;
signal \N__64617\ : std_logic;
signal \N__64614\ : std_logic;
signal \N__64611\ : std_logic;
signal \N__64608\ : std_logic;
signal \N__64605\ : std_logic;
signal \N__64602\ : std_logic;
signal \N__64599\ : std_logic;
signal \N__64596\ : std_logic;
signal \N__64593\ : std_logic;
signal \N__64590\ : std_logic;
signal \N__64587\ : std_logic;
signal \N__64584\ : std_logic;
signal \N__64583\ : std_logic;
signal \N__64582\ : std_logic;
signal \N__64581\ : std_logic;
signal \N__64578\ : std_logic;
signal \N__64577\ : std_logic;
signal \N__64576\ : std_logic;
signal \N__64575\ : std_logic;
signal \N__64574\ : std_logic;
signal \N__64573\ : std_logic;
signal \N__64572\ : std_logic;
signal \N__64571\ : std_logic;
signal \N__64570\ : std_logic;
signal \N__64561\ : std_logic;
signal \N__64552\ : std_logic;
signal \N__64551\ : std_logic;
signal \N__64542\ : std_logic;
signal \N__64539\ : std_logic;
signal \N__64536\ : std_logic;
signal \N__64533\ : std_logic;
signal \N__64526\ : std_logic;
signal \N__64523\ : std_logic;
signal \N__64518\ : std_logic;
signal \N__64515\ : std_logic;
signal \N__64512\ : std_logic;
signal \N__64509\ : std_logic;
signal \N__64506\ : std_logic;
signal \N__64503\ : std_logic;
signal \N__64500\ : std_logic;
signal \N__64497\ : std_logic;
signal \N__64496\ : std_logic;
signal \N__64493\ : std_logic;
signal \N__64490\ : std_logic;
signal \N__64485\ : std_logic;
signal \N__64482\ : std_logic;
signal \N__64479\ : std_logic;
signal \N__64476\ : std_logic;
signal \N__64473\ : std_logic;
signal \N__64472\ : std_logic;
signal \N__64469\ : std_logic;
signal \N__64466\ : std_logic;
signal \N__64465\ : std_logic;
signal \N__64462\ : std_logic;
signal \N__64459\ : std_logic;
signal \N__64458\ : std_logic;
signal \N__64457\ : std_logic;
signal \N__64454\ : std_logic;
signal \N__64449\ : std_logic;
signal \N__64444\ : std_logic;
signal \N__64437\ : std_logic;
signal \N__64434\ : std_logic;
signal \N__64433\ : std_logic;
signal \N__64432\ : std_logic;
signal \N__64429\ : std_logic;
signal \N__64426\ : std_logic;
signal \N__64425\ : std_logic;
signal \N__64422\ : std_logic;
signal \N__64421\ : std_logic;
signal \N__64420\ : std_logic;
signal \N__64417\ : std_logic;
signal \N__64414\ : std_logic;
signal \N__64411\ : std_logic;
signal \N__64408\ : std_logic;
signal \N__64407\ : std_logic;
signal \N__64406\ : std_logic;
signal \N__64401\ : std_logic;
signal \N__64398\ : std_logic;
signal \N__64393\ : std_logic;
signal \N__64390\ : std_logic;
signal \N__64385\ : std_logic;
signal \N__64374\ : std_logic;
signal \N__64371\ : std_logic;
signal \N__64368\ : std_logic;
signal \N__64365\ : std_logic;
signal \N__64362\ : std_logic;
signal \N__64359\ : std_logic;
signal \N__64356\ : std_logic;
signal \N__64355\ : std_logic;
signal \N__64352\ : std_logic;
signal \N__64349\ : std_logic;
signal \N__64344\ : std_logic;
signal \N__64343\ : std_logic;
signal \N__64340\ : std_logic;
signal \N__64337\ : std_logic;
signal \N__64334\ : std_logic;
signal \N__64331\ : std_logic;
signal \N__64328\ : std_logic;
signal \N__64323\ : std_logic;
signal \N__64320\ : std_logic;
signal \N__64317\ : std_logic;
signal \N__64316\ : std_logic;
signal \N__64313\ : std_logic;
signal \N__64312\ : std_logic;
signal \N__64309\ : std_logic;
signal \N__64306\ : std_logic;
signal \N__64303\ : std_logic;
signal \N__64300\ : std_logic;
signal \N__64299\ : std_logic;
signal \N__64296\ : std_logic;
signal \N__64293\ : std_logic;
signal \N__64290\ : std_logic;
signal \N__64287\ : std_logic;
signal \N__64284\ : std_logic;
signal \N__64281\ : std_logic;
signal \N__64274\ : std_logic;
signal \N__64269\ : std_logic;
signal \N__64268\ : std_logic;
signal \N__64267\ : std_logic;
signal \N__64266\ : std_logic;
signal \N__64265\ : std_logic;
signal \N__64262\ : std_logic;
signal \N__64261\ : std_logic;
signal \N__64260\ : std_logic;
signal \N__64259\ : std_logic;
signal \N__64256\ : std_logic;
signal \N__64253\ : std_logic;
signal \N__64252\ : std_logic;
signal \N__64251\ : std_logic;
signal \N__64250\ : std_logic;
signal \N__64249\ : std_logic;
signal \N__64248\ : std_logic;
signal \N__64247\ : std_logic;
signal \N__64246\ : std_logic;
signal \N__64245\ : std_logic;
signal \N__64244\ : std_logic;
signal \N__64243\ : std_logic;
signal \N__64240\ : std_logic;
signal \N__64237\ : std_logic;
signal \N__64236\ : std_logic;
signal \N__64235\ : std_logic;
signal \N__64234\ : std_logic;
signal \N__64231\ : std_logic;
signal \N__64230\ : std_logic;
signal \N__64229\ : std_logic;
signal \N__64228\ : std_logic;
signal \N__64225\ : std_logic;
signal \N__64220\ : std_logic;
signal \N__64219\ : std_logic;
signal \N__64218\ : std_logic;
signal \N__64217\ : std_logic;
signal \N__64216\ : std_logic;
signal \N__64215\ : std_logic;
signal \N__64214\ : std_logic;
signal \N__64213\ : std_logic;
signal \N__64210\ : std_logic;
signal \N__64209\ : std_logic;
signal \N__64208\ : std_logic;
signal \N__64207\ : std_logic;
signal \N__64206\ : std_logic;
signal \N__64205\ : std_logic;
signal \N__64204\ : std_logic;
signal \N__64203\ : std_logic;
signal \N__64202\ : std_logic;
signal \N__64201\ : std_logic;
signal \N__64198\ : std_logic;
signal \N__64193\ : std_logic;
signal \N__64190\ : std_logic;
signal \N__64175\ : std_logic;
signal \N__64174\ : std_logic;
signal \N__64173\ : std_logic;
signal \N__64172\ : std_logic;
signal \N__64169\ : std_logic;
signal \N__64166\ : std_logic;
signal \N__64161\ : std_logic;
signal \N__64158\ : std_logic;
signal \N__64157\ : std_logic;
signal \N__64154\ : std_logic;
signal \N__64153\ : std_logic;
signal \N__64152\ : std_logic;
signal \N__64149\ : std_logic;
signal \N__64144\ : std_logic;
signal \N__64139\ : std_logic;
signal \N__64124\ : std_logic;
signal \N__64121\ : std_logic;
signal \N__64118\ : std_logic;
signal \N__64117\ : std_logic;
signal \N__64100\ : std_logic;
signal \N__64095\ : std_logic;
signal \N__64092\ : std_logic;
signal \N__64089\ : std_logic;
signal \N__64082\ : std_logic;
signal \N__64081\ : std_logic;
signal \N__64078\ : std_logic;
signal \N__64075\ : std_logic;
signal \N__64074\ : std_logic;
signal \N__64073\ : std_logic;
signal \N__64072\ : std_logic;
signal \N__64071\ : std_logic;
signal \N__64070\ : std_logic;
signal \N__64069\ : std_logic;
signal \N__64068\ : std_logic;
signal \N__64067\ : std_logic;
signal \N__64066\ : std_logic;
signal \N__64061\ : std_logic;
signal \N__64058\ : std_logic;
signal \N__64055\ : std_logic;
signal \N__64050\ : std_logic;
signal \N__64043\ : std_logic;
signal \N__64038\ : std_logic;
signal \N__64033\ : std_logic;
signal \N__64028\ : std_logic;
signal \N__64021\ : std_logic;
signal \N__64018\ : std_logic;
signal \N__64013\ : std_logic;
signal \N__64010\ : std_logic;
signal \N__64007\ : std_logic;
signal \N__64000\ : std_logic;
signal \N__63991\ : std_logic;
signal \N__63988\ : std_logic;
signal \N__63977\ : std_logic;
signal \N__63970\ : std_logic;
signal \N__63951\ : std_logic;
signal \N__63948\ : std_logic;
signal \N__63945\ : std_logic;
signal \N__63944\ : std_logic;
signal \N__63941\ : std_logic;
signal \N__63940\ : std_logic;
signal \N__63939\ : std_logic;
signal \N__63936\ : std_logic;
signal \N__63933\ : std_logic;
signal \N__63930\ : std_logic;
signal \N__63927\ : std_logic;
signal \N__63924\ : std_logic;
signal \N__63923\ : std_logic;
signal \N__63918\ : std_logic;
signal \N__63915\ : std_logic;
signal \N__63914\ : std_logic;
signal \N__63911\ : std_logic;
signal \N__63910\ : std_logic;
signal \N__63909\ : std_logic;
signal \N__63906\ : std_logic;
signal \N__63905\ : std_logic;
signal \N__63902\ : std_logic;
signal \N__63899\ : std_logic;
signal \N__63896\ : std_logic;
signal \N__63893\ : std_logic;
signal \N__63890\ : std_logic;
signal \N__63887\ : std_logic;
signal \N__63884\ : std_logic;
signal \N__63881\ : std_logic;
signal \N__63878\ : std_logic;
signal \N__63873\ : std_logic;
signal \N__63870\ : std_logic;
signal \N__63867\ : std_logic;
signal \N__63864\ : std_logic;
signal \N__63859\ : std_logic;
signal \N__63854\ : std_logic;
signal \N__63851\ : std_logic;
signal \N__63844\ : std_logic;
signal \N__63837\ : std_logic;
signal \N__63834\ : std_logic;
signal \N__63831\ : std_logic;
signal \N__63828\ : std_logic;
signal \N__63827\ : std_logic;
signal \N__63826\ : std_logic;
signal \N__63823\ : std_logic;
signal \N__63822\ : std_logic;
signal \N__63819\ : std_logic;
signal \N__63816\ : std_logic;
signal \N__63813\ : std_logic;
signal \N__63810\ : std_logic;
signal \N__63809\ : std_logic;
signal \N__63806\ : std_logic;
signal \N__63803\ : std_logic;
signal \N__63800\ : std_logic;
signal \N__63799\ : std_logic;
signal \N__63796\ : std_logic;
signal \N__63793\ : std_logic;
signal \N__63790\ : std_logic;
signal \N__63789\ : std_logic;
signal \N__63786\ : std_logic;
signal \N__63785\ : std_logic;
signal \N__63782\ : std_logic;
signal \N__63779\ : std_logic;
signal \N__63776\ : std_logic;
signal \N__63775\ : std_logic;
signal \N__63770\ : std_logic;
signal \N__63767\ : std_logic;
signal \N__63764\ : std_logic;
signal \N__63761\ : std_logic;
signal \N__63756\ : std_logic;
signal \N__63753\ : std_logic;
signal \N__63750\ : std_logic;
signal \N__63747\ : std_logic;
signal \N__63742\ : std_logic;
signal \N__63739\ : std_logic;
signal \N__63736\ : std_logic;
signal \N__63733\ : std_logic;
signal \N__63730\ : std_logic;
signal \N__63727\ : std_logic;
signal \N__63724\ : std_logic;
signal \N__63719\ : std_logic;
signal \N__63708\ : std_logic;
signal \N__63705\ : std_logic;
signal \N__63702\ : std_logic;
signal \N__63701\ : std_logic;
signal \N__63698\ : std_logic;
signal \N__63697\ : std_logic;
signal \N__63694\ : std_logic;
signal \N__63691\ : std_logic;
signal \N__63688\ : std_logic;
signal \N__63687\ : std_logic;
signal \N__63684\ : std_logic;
signal \N__63681\ : std_logic;
signal \N__63678\ : std_logic;
signal \N__63677\ : std_logic;
signal \N__63674\ : std_logic;
signal \N__63671\ : std_logic;
signal \N__63670\ : std_logic;
signal \N__63665\ : std_logic;
signal \N__63662\ : std_logic;
signal \N__63661\ : std_logic;
signal \N__63658\ : std_logic;
signal \N__63657\ : std_logic;
signal \N__63654\ : std_logic;
signal \N__63651\ : std_logic;
signal \N__63646\ : std_logic;
signal \N__63645\ : std_logic;
signal \N__63642\ : std_logic;
signal \N__63639\ : std_logic;
signal \N__63636\ : std_logic;
signal \N__63633\ : std_logic;
signal \N__63630\ : std_logic;
signal \N__63627\ : std_logic;
signal \N__63624\ : std_logic;
signal \N__63621\ : std_logic;
signal \N__63612\ : std_logic;
signal \N__63609\ : std_logic;
signal \N__63606\ : std_logic;
signal \N__63603\ : std_logic;
signal \N__63600\ : std_logic;
signal \N__63591\ : std_logic;
signal \N__63588\ : std_logic;
signal \N__63585\ : std_logic;
signal \N__63584\ : std_logic;
signal \N__63583\ : std_logic;
signal \N__63582\ : std_logic;
signal \N__63581\ : std_logic;
signal \N__63580\ : std_logic;
signal \N__63577\ : std_logic;
signal \N__63574\ : std_logic;
signal \N__63569\ : std_logic;
signal \N__63568\ : std_logic;
signal \N__63565\ : std_logic;
signal \N__63562\ : std_logic;
signal \N__63559\ : std_logic;
signal \N__63556\ : std_logic;
signal \N__63553\ : std_logic;
signal \N__63550\ : std_logic;
signal \N__63547\ : std_logic;
signal \N__63544\ : std_logic;
signal \N__63543\ : std_logic;
signal \N__63540\ : std_logic;
signal \N__63537\ : std_logic;
signal \N__63532\ : std_logic;
signal \N__63527\ : std_logic;
signal \N__63526\ : std_logic;
signal \N__63523\ : std_logic;
signal \N__63520\ : std_logic;
signal \N__63517\ : std_logic;
signal \N__63514\ : std_logic;
signal \N__63511\ : std_logic;
signal \N__63508\ : std_logic;
signal \N__63503\ : std_logic;
signal \N__63498\ : std_logic;
signal \N__63489\ : std_logic;
signal \N__63486\ : std_logic;
signal \N__63483\ : std_logic;
signal \N__63482\ : std_logic;
signal \N__63481\ : std_logic;
signal \N__63478\ : std_logic;
signal \N__63477\ : std_logic;
signal \N__63476\ : std_logic;
signal \N__63473\ : std_logic;
signal \N__63472\ : std_logic;
signal \N__63471\ : std_logic;
signal \N__63468\ : std_logic;
signal \N__63467\ : std_logic;
signal \N__63464\ : std_logic;
signal \N__63461\ : std_logic;
signal \N__63458\ : std_logic;
signal \N__63455\ : std_logic;
signal \N__63452\ : std_logic;
signal \N__63449\ : std_logic;
signal \N__63448\ : std_logic;
signal \N__63445\ : std_logic;
signal \N__63442\ : std_logic;
signal \N__63439\ : std_logic;
signal \N__63436\ : std_logic;
signal \N__63433\ : std_logic;
signal \N__63430\ : std_logic;
signal \N__63427\ : std_logic;
signal \N__63424\ : std_logic;
signal \N__63421\ : std_logic;
signal \N__63418\ : std_logic;
signal \N__63407\ : std_logic;
signal \N__63400\ : std_logic;
signal \N__63397\ : std_logic;
signal \N__63394\ : std_logic;
signal \N__63391\ : std_logic;
signal \N__63384\ : std_logic;
signal \N__63383\ : std_logic;
signal \N__63382\ : std_logic;
signal \N__63381\ : std_logic;
signal \N__63380\ : std_logic;
signal \N__63379\ : std_logic;
signal \N__63378\ : std_logic;
signal \N__63377\ : std_logic;
signal \N__63376\ : std_logic;
signal \N__63359\ : std_logic;
signal \N__63356\ : std_logic;
signal \N__63355\ : std_logic;
signal \N__63354\ : std_logic;
signal \N__63353\ : std_logic;
signal \N__63352\ : std_logic;
signal \N__63351\ : std_logic;
signal \N__63350\ : std_logic;
signal \N__63349\ : std_logic;
signal \N__63348\ : std_logic;
signal \N__63347\ : std_logic;
signal \N__63346\ : std_logic;
signal \N__63345\ : std_logic;
signal \N__63344\ : std_logic;
signal \N__63343\ : std_logic;
signal \N__63342\ : std_logic;
signal \N__63341\ : std_logic;
signal \N__63338\ : std_logic;
signal \N__63327\ : std_logic;
signal \N__63310\ : std_logic;
signal \N__63303\ : std_logic;
signal \N__63302\ : std_logic;
signal \N__63301\ : std_logic;
signal \N__63300\ : std_logic;
signal \N__63299\ : std_logic;
signal \N__63298\ : std_logic;
signal \N__63297\ : std_logic;
signal \N__63296\ : std_logic;
signal \N__63295\ : std_logic;
signal \N__63294\ : std_logic;
signal \N__63293\ : std_logic;
signal \N__63292\ : std_logic;
signal \N__63285\ : std_logic;
signal \N__63282\ : std_logic;
signal \N__63281\ : std_logic;
signal \N__63278\ : std_logic;
signal \N__63275\ : std_logic;
signal \N__63274\ : std_logic;
signal \N__63273\ : std_logic;
signal \N__63270\ : std_logic;
signal \N__63255\ : std_logic;
signal \N__63252\ : std_logic;
signal \N__63247\ : std_logic;
signal \N__63246\ : std_logic;
signal \N__63243\ : std_logic;
signal \N__63238\ : std_logic;
signal \N__63235\ : std_logic;
signal \N__63232\ : std_logic;
signal \N__63231\ : std_logic;
signal \N__63230\ : std_logic;
signal \N__63225\ : std_logic;
signal \N__63222\ : std_logic;
signal \N__63219\ : std_logic;
signal \N__63216\ : std_logic;
signal \N__63211\ : std_logic;
signal \N__63202\ : std_logic;
signal \N__63199\ : std_logic;
signal \N__63198\ : std_logic;
signal \N__63197\ : std_logic;
signal \N__63194\ : std_logic;
signal \N__63191\ : std_logic;
signal \N__63188\ : std_logic;
signal \N__63183\ : std_logic;
signal \N__63180\ : std_logic;
signal \N__63175\ : std_logic;
signal \N__63170\ : std_logic;
signal \N__63163\ : std_logic;
signal \N__63156\ : std_logic;
signal \N__63153\ : std_logic;
signal \N__63150\ : std_logic;
signal \N__63149\ : std_logic;
signal \N__63146\ : std_logic;
signal \N__63145\ : std_logic;
signal \N__63144\ : std_logic;
signal \N__63141\ : std_logic;
signal \N__63138\ : std_logic;
signal \N__63135\ : std_logic;
signal \N__63134\ : std_logic;
signal \N__63131\ : std_logic;
signal \N__63128\ : std_logic;
signal \N__63123\ : std_logic;
signal \N__63120\ : std_logic;
signal \N__63119\ : std_logic;
signal \N__63118\ : std_logic;
signal \N__63115\ : std_logic;
signal \N__63110\ : std_logic;
signal \N__63107\ : std_logic;
signal \N__63104\ : std_logic;
signal \N__63103\ : std_logic;
signal \N__63102\ : std_logic;
signal \N__63099\ : std_logic;
signal \N__63094\ : std_logic;
signal \N__63091\ : std_logic;
signal \N__63088\ : std_logic;
signal \N__63083\ : std_logic;
signal \N__63080\ : std_logic;
signal \N__63077\ : std_logic;
signal \N__63074\ : std_logic;
signal \N__63071\ : std_logic;
signal \N__63068\ : std_logic;
signal \N__63065\ : std_logic;
signal \N__63062\ : std_logic;
signal \N__63059\ : std_logic;
signal \N__63054\ : std_logic;
signal \N__63045\ : std_logic;
signal \N__63042\ : std_logic;
signal \N__63039\ : std_logic;
signal \N__63036\ : std_logic;
signal \N__63033\ : std_logic;
signal \N__63030\ : std_logic;
signal \N__63029\ : std_logic;
signal \N__63026\ : std_logic;
signal \N__63025\ : std_logic;
signal \N__63022\ : std_logic;
signal \N__63019\ : std_logic;
signal \N__63016\ : std_logic;
signal \N__63015\ : std_logic;
signal \N__63012\ : std_logic;
signal \N__63007\ : std_logic;
signal \N__63004\ : std_logic;
signal \N__63003\ : std_logic;
signal \N__63002\ : std_logic;
signal \N__62999\ : std_logic;
signal \N__62994\ : std_logic;
signal \N__62991\ : std_logic;
signal \N__62988\ : std_logic;
signal \N__62985\ : std_logic;
signal \N__62980\ : std_logic;
signal \N__62977\ : std_logic;
signal \N__62974\ : std_logic;
signal \N__62971\ : std_logic;
signal \N__62968\ : std_logic;
signal \N__62961\ : std_logic;
signal \N__62960\ : std_logic;
signal \N__62959\ : std_logic;
signal \N__62958\ : std_logic;
signal \N__62957\ : std_logic;
signal \N__62956\ : std_logic;
signal \N__62955\ : std_logic;
signal \N__62954\ : std_logic;
signal \N__62953\ : std_logic;
signal \N__62952\ : std_logic;
signal \N__62951\ : std_logic;
signal \N__62950\ : std_logic;
signal \N__62949\ : std_logic;
signal \N__62948\ : std_logic;
signal \N__62947\ : std_logic;
signal \N__62946\ : std_logic;
signal \N__62945\ : std_logic;
signal \N__62944\ : std_logic;
signal \N__62943\ : std_logic;
signal \N__62942\ : std_logic;
signal \N__62941\ : std_logic;
signal \N__62940\ : std_logic;
signal \N__62939\ : std_logic;
signal \N__62938\ : std_logic;
signal \N__62937\ : std_logic;
signal \N__62936\ : std_logic;
signal \N__62935\ : std_logic;
signal \N__62934\ : std_logic;
signal \N__62933\ : std_logic;
signal \N__62932\ : std_logic;
signal \N__62931\ : std_logic;
signal \N__62930\ : std_logic;
signal \N__62929\ : std_logic;
signal \N__62928\ : std_logic;
signal \N__62927\ : std_logic;
signal \N__62926\ : std_logic;
signal \N__62925\ : std_logic;
signal \N__62924\ : std_logic;
signal \N__62923\ : std_logic;
signal \N__62922\ : std_logic;
signal \N__62921\ : std_logic;
signal \N__62920\ : std_logic;
signal \N__62919\ : std_logic;
signal \N__62918\ : std_logic;
signal \N__62917\ : std_logic;
signal \N__62916\ : std_logic;
signal \N__62915\ : std_logic;
signal \N__62914\ : std_logic;
signal \N__62913\ : std_logic;
signal \N__62912\ : std_logic;
signal \N__62911\ : std_logic;
signal \N__62910\ : std_logic;
signal \N__62909\ : std_logic;
signal \N__62908\ : std_logic;
signal \N__62907\ : std_logic;
signal \N__62906\ : std_logic;
signal \N__62905\ : std_logic;
signal \N__62904\ : std_logic;
signal \N__62903\ : std_logic;
signal \N__62902\ : std_logic;
signal \N__62901\ : std_logic;
signal \N__62900\ : std_logic;
signal \N__62899\ : std_logic;
signal \N__62898\ : std_logic;
signal \N__62897\ : std_logic;
signal \N__62896\ : std_logic;
signal \N__62895\ : std_logic;
signal \N__62894\ : std_logic;
signal \N__62893\ : std_logic;
signal \N__62892\ : std_logic;
signal \N__62891\ : std_logic;
signal \N__62890\ : std_logic;
signal \N__62889\ : std_logic;
signal \N__62888\ : std_logic;
signal \N__62887\ : std_logic;
signal \N__62886\ : std_logic;
signal \N__62885\ : std_logic;
signal \N__62884\ : std_logic;
signal \N__62883\ : std_logic;
signal \N__62882\ : std_logic;
signal \N__62881\ : std_logic;
signal \N__62880\ : std_logic;
signal \N__62879\ : std_logic;
signal \N__62878\ : std_logic;
signal \N__62877\ : std_logic;
signal \N__62876\ : std_logic;
signal \N__62875\ : std_logic;
signal \N__62874\ : std_logic;
signal \N__62873\ : std_logic;
signal \N__62872\ : std_logic;
signal \N__62871\ : std_logic;
signal \N__62870\ : std_logic;
signal \N__62869\ : std_logic;
signal \N__62868\ : std_logic;
signal \N__62867\ : std_logic;
signal \N__62866\ : std_logic;
signal \N__62865\ : std_logic;
signal \N__62864\ : std_logic;
signal \N__62863\ : std_logic;
signal \N__62862\ : std_logic;
signal \N__62861\ : std_logic;
signal \N__62860\ : std_logic;
signal \N__62859\ : std_logic;
signal \N__62858\ : std_logic;
signal \N__62857\ : std_logic;
signal \N__62856\ : std_logic;
signal \N__62855\ : std_logic;
signal \N__62854\ : std_logic;
signal \N__62853\ : std_logic;
signal \N__62852\ : std_logic;
signal \N__62851\ : std_logic;
signal \N__62850\ : std_logic;
signal \N__62849\ : std_logic;
signal \N__62848\ : std_logic;
signal \N__62847\ : std_logic;
signal \N__62846\ : std_logic;
signal \N__62845\ : std_logic;
signal \N__62844\ : std_logic;
signal \N__62843\ : std_logic;
signal \N__62842\ : std_logic;
signal \N__62841\ : std_logic;
signal \N__62840\ : std_logic;
signal \N__62839\ : std_logic;
signal \N__62838\ : std_logic;
signal \N__62837\ : std_logic;
signal \N__62836\ : std_logic;
signal \N__62835\ : std_logic;
signal \N__62834\ : std_logic;
signal \N__62833\ : std_logic;
signal \N__62832\ : std_logic;
signal \N__62831\ : std_logic;
signal \N__62830\ : std_logic;
signal \N__62829\ : std_logic;
signal \N__62828\ : std_logic;
signal \N__62827\ : std_logic;
signal \N__62826\ : std_logic;
signal \N__62825\ : std_logic;
signal \N__62824\ : std_logic;
signal \N__62823\ : std_logic;
signal \N__62822\ : std_logic;
signal \N__62821\ : std_logic;
signal \N__62820\ : std_logic;
signal \N__62819\ : std_logic;
signal \N__62818\ : std_logic;
signal \N__62817\ : std_logic;
signal \N__62816\ : std_logic;
signal \N__62815\ : std_logic;
signal \N__62814\ : std_logic;
signal \N__62813\ : std_logic;
signal \N__62812\ : std_logic;
signal \N__62811\ : std_logic;
signal \N__62810\ : std_logic;
signal \N__62809\ : std_logic;
signal \N__62808\ : std_logic;
signal \N__62807\ : std_logic;
signal \N__62806\ : std_logic;
signal \N__62805\ : std_logic;
signal \N__62804\ : std_logic;
signal \N__62487\ : std_logic;
signal \N__62484\ : std_logic;
signal \N__62481\ : std_logic;
signal \N__62480\ : std_logic;
signal \N__62479\ : std_logic;
signal \N__62476\ : std_logic;
signal \N__62473\ : std_logic;
signal \N__62472\ : std_logic;
signal \N__62469\ : std_logic;
signal \N__62466\ : std_logic;
signal \N__62463\ : std_logic;
signal \N__62460\ : std_logic;
signal \N__62457\ : std_logic;
signal \N__62456\ : std_logic;
signal \N__62455\ : std_logic;
signal \N__62452\ : std_logic;
signal \N__62447\ : std_logic;
signal \N__62444\ : std_logic;
signal \N__62441\ : std_logic;
signal \N__62438\ : std_logic;
signal \N__62433\ : std_logic;
signal \N__62428\ : std_logic;
signal \N__62421\ : std_logic;
signal \N__62420\ : std_logic;
signal \N__62417\ : std_logic;
signal \N__62414\ : std_logic;
signal \N__62411\ : std_logic;
signal \N__62406\ : std_logic;
signal \N__62403\ : std_logic;
signal \N__62402\ : std_logic;
signal \N__62399\ : std_logic;
signal \N__62396\ : std_logic;
signal \N__62393\ : std_logic;
signal \N__62390\ : std_logic;
signal \N__62387\ : std_logic;
signal \N__62382\ : std_logic;
signal \N__62379\ : std_logic;
signal \N__62376\ : std_logic;
signal \N__62373\ : std_logic;
signal \N__62370\ : std_logic;
signal \N__62369\ : std_logic;
signal \N__62368\ : std_logic;
signal \N__62367\ : std_logic;
signal \N__62364\ : std_logic;
signal \N__62361\ : std_logic;
signal \N__62358\ : std_logic;
signal \N__62357\ : std_logic;
signal \N__62356\ : std_logic;
signal \N__62353\ : std_logic;
signal \N__62350\ : std_logic;
signal \N__62347\ : std_logic;
signal \N__62344\ : std_logic;
signal \N__62341\ : std_logic;
signal \N__62338\ : std_logic;
signal \N__62337\ : std_logic;
signal \N__62336\ : std_logic;
signal \N__62333\ : std_logic;
signal \N__62330\ : std_logic;
signal \N__62327\ : std_logic;
signal \N__62320\ : std_logic;
signal \N__62317\ : std_logic;
signal \N__62314\ : std_logic;
signal \N__62311\ : std_logic;
signal \N__62306\ : std_logic;
signal \N__62303\ : std_logic;
signal \N__62300\ : std_logic;
signal \N__62295\ : std_logic;
signal \N__62292\ : std_logic;
signal \N__62289\ : std_logic;
signal \N__62286\ : std_logic;
signal \N__62281\ : std_logic;
signal \N__62276\ : std_logic;
signal \N__62271\ : std_logic;
signal \N__62268\ : std_logic;
signal \N__62265\ : std_logic;
signal \N__62264\ : std_logic;
signal \N__62263\ : std_logic;
signal \N__62262\ : std_logic;
signal \N__62261\ : std_logic;
signal \N__62260\ : std_logic;
signal \N__62259\ : std_logic;
signal \N__62256\ : std_logic;
signal \N__62253\ : std_logic;
signal \N__62250\ : std_logic;
signal \N__62247\ : std_logic;
signal \N__62246\ : std_logic;
signal \N__62243\ : std_logic;
signal \N__62240\ : std_logic;
signal \N__62237\ : std_logic;
signal \N__62234\ : std_logic;
signal \N__62231\ : std_logic;
signal \N__62226\ : std_logic;
signal \N__62223\ : std_logic;
signal \N__62218\ : std_logic;
signal \N__62215\ : std_logic;
signal \N__62212\ : std_logic;
signal \N__62209\ : std_logic;
signal \N__62206\ : std_logic;
signal \N__62197\ : std_logic;
signal \N__62190\ : std_logic;
signal \N__62187\ : std_logic;
signal \N__62184\ : std_logic;
signal \N__62183\ : std_logic;
signal \N__62180\ : std_logic;
signal \N__62179\ : std_logic;
signal \N__62176\ : std_logic;
signal \N__62173\ : std_logic;
signal \N__62170\ : std_logic;
signal \N__62169\ : std_logic;
signal \N__62166\ : std_logic;
signal \N__62165\ : std_logic;
signal \N__62160\ : std_logic;
signal \N__62157\ : std_logic;
signal \N__62154\ : std_logic;
signal \N__62151\ : std_logic;
signal \N__62148\ : std_logic;
signal \N__62147\ : std_logic;
signal \N__62144\ : std_logic;
signal \N__62139\ : std_logic;
signal \N__62136\ : std_logic;
signal \N__62133\ : std_logic;
signal \N__62132\ : std_logic;
signal \N__62129\ : std_logic;
signal \N__62126\ : std_logic;
signal \N__62125\ : std_logic;
signal \N__62120\ : std_logic;
signal \N__62117\ : std_logic;
signal \N__62114\ : std_logic;
signal \N__62111\ : std_logic;
signal \N__62108\ : std_logic;
signal \N__62105\ : std_logic;
signal \N__62102\ : std_logic;
signal \N__62097\ : std_logic;
signal \N__62090\ : std_logic;
signal \N__62087\ : std_logic;
signal \N__62084\ : std_logic;
signal \N__62079\ : std_logic;
signal \N__62076\ : std_logic;
signal \N__62073\ : std_logic;
signal \N__62072\ : std_logic;
signal \N__62071\ : std_logic;
signal \N__62070\ : std_logic;
signal \N__62067\ : std_logic;
signal \N__62064\ : std_logic;
signal \N__62061\ : std_logic;
signal \N__62060\ : std_logic;
signal \N__62059\ : std_logic;
signal \N__62056\ : std_logic;
signal \N__62051\ : std_logic;
signal \N__62048\ : std_logic;
signal \N__62045\ : std_logic;
signal \N__62044\ : std_logic;
signal \N__62041\ : std_logic;
signal \N__62038\ : std_logic;
signal \N__62033\ : std_logic;
signal \N__62028\ : std_logic;
signal \N__62025\ : std_logic;
signal \N__62024\ : std_logic;
signal \N__62019\ : std_logic;
signal \N__62016\ : std_logic;
signal \N__62013\ : std_logic;
signal \N__62010\ : std_logic;
signal \N__62007\ : std_logic;
signal \N__62004\ : std_logic;
signal \N__62001\ : std_logic;
signal \N__61994\ : std_logic;
signal \N__61989\ : std_logic;
signal \N__61986\ : std_logic;
signal \N__61983\ : std_logic;
signal \N__61980\ : std_logic;
signal \N__61977\ : std_logic;
signal \N__61974\ : std_logic;
signal \N__61971\ : std_logic;
signal \N__61970\ : std_logic;
signal \N__61969\ : std_logic;
signal \N__61968\ : std_logic;
signal \N__61965\ : std_logic;
signal \N__61964\ : std_logic;
signal \N__61963\ : std_logic;
signal \N__61960\ : std_logic;
signal \N__61959\ : std_logic;
signal \N__61956\ : std_logic;
signal \N__61953\ : std_logic;
signal \N__61950\ : std_logic;
signal \N__61947\ : std_logic;
signal \N__61944\ : std_logic;
signal \N__61943\ : std_logic;
signal \N__61940\ : std_logic;
signal \N__61937\ : std_logic;
signal \N__61934\ : std_logic;
signal \N__61931\ : std_logic;
signal \N__61930\ : std_logic;
signal \N__61927\ : std_logic;
signal \N__61922\ : std_logic;
signal \N__61919\ : std_logic;
signal \N__61910\ : std_logic;
signal \N__61907\ : std_logic;
signal \N__61904\ : std_logic;
signal \N__61901\ : std_logic;
signal \N__61898\ : std_logic;
signal \N__61895\ : std_logic;
signal \N__61890\ : std_logic;
signal \N__61887\ : std_logic;
signal \N__61878\ : std_logic;
signal \N__61875\ : std_logic;
signal \N__61872\ : std_logic;
signal \N__61871\ : std_logic;
signal \N__61868\ : std_logic;
signal \N__61867\ : std_logic;
signal \N__61864\ : std_logic;
signal \N__61863\ : std_logic;
signal \N__61862\ : std_logic;
signal \N__61861\ : std_logic;
signal \N__61860\ : std_logic;
signal \N__61859\ : std_logic;
signal \N__61856\ : std_logic;
signal \N__61853\ : std_logic;
signal \N__61850\ : std_logic;
signal \N__61847\ : std_logic;
signal \N__61844\ : std_logic;
signal \N__61841\ : std_logic;
signal \N__61838\ : std_logic;
signal \N__61835\ : std_logic;
signal \N__61832\ : std_logic;
signal \N__61827\ : std_logic;
signal \N__61824\ : std_logic;
signal \N__61821\ : std_logic;
signal \N__61820\ : std_logic;
signal \N__61817\ : std_logic;
signal \N__61814\ : std_logic;
signal \N__61811\ : std_logic;
signal \N__61808\ : std_logic;
signal \N__61803\ : std_logic;
signal \N__61800\ : std_logic;
signal \N__61797\ : std_logic;
signal \N__61794\ : std_logic;
signal \N__61791\ : std_logic;
signal \N__61788\ : std_logic;
signal \N__61785\ : std_logic;
signal \N__61782\ : std_logic;
signal \N__61779\ : std_logic;
signal \N__61776\ : std_logic;
signal \N__61773\ : std_logic;
signal \N__61766\ : std_logic;
signal \N__61759\ : std_logic;
signal \N__61752\ : std_logic;
signal \N__61749\ : std_logic;
signal \N__61746\ : std_logic;
signal \N__61745\ : std_logic;
signal \N__61742\ : std_logic;
signal \N__61739\ : std_logic;
signal \N__61738\ : std_logic;
signal \N__61737\ : std_logic;
signal \N__61734\ : std_logic;
signal \N__61731\ : std_logic;
signal \N__61730\ : std_logic;
signal \N__61729\ : std_logic;
signal \N__61726\ : std_logic;
signal \N__61723\ : std_logic;
signal \N__61720\ : std_logic;
signal \N__61719\ : std_logic;
signal \N__61716\ : std_logic;
signal \N__61713\ : std_logic;
signal \N__61712\ : std_logic;
signal \N__61711\ : std_logic;
signal \N__61708\ : std_logic;
signal \N__61705\ : std_logic;
signal \N__61700\ : std_logic;
signal \N__61697\ : std_logic;
signal \N__61694\ : std_logic;
signal \N__61691\ : std_logic;
signal \N__61688\ : std_logic;
signal \N__61685\ : std_logic;
signal \N__61682\ : std_logic;
signal \N__61675\ : std_logic;
signal \N__61670\ : std_logic;
signal \N__61667\ : std_logic;
signal \N__61662\ : std_logic;
signal \N__61659\ : std_logic;
signal \N__61656\ : std_logic;
signal \N__61647\ : std_logic;
signal \N__61646\ : std_logic;
signal \N__61645\ : std_logic;
signal \N__61644\ : std_logic;
signal \N__61641\ : std_logic;
signal \N__61640\ : std_logic;
signal \N__61639\ : std_logic;
signal \N__61636\ : std_logic;
signal \N__61633\ : std_logic;
signal \N__61632\ : std_logic;
signal \N__61631\ : std_logic;
signal \N__61628\ : std_logic;
signal \N__61625\ : std_logic;
signal \N__61622\ : std_logic;
signal \N__61619\ : std_logic;
signal \N__61614\ : std_logic;
signal \N__61613\ : std_logic;
signal \N__61610\ : std_logic;
signal \N__61607\ : std_logic;
signal \N__61604\ : std_logic;
signal \N__61599\ : std_logic;
signal \N__61596\ : std_logic;
signal \N__61593\ : std_logic;
signal \N__61590\ : std_logic;
signal \N__61587\ : std_logic;
signal \N__61580\ : std_logic;
signal \N__61575\ : std_logic;
signal \N__61572\ : std_logic;
signal \N__61569\ : std_logic;
signal \N__61566\ : std_logic;
signal \N__61559\ : std_logic;
signal \N__61554\ : std_logic;
signal \N__61551\ : std_logic;
signal \N__61548\ : std_logic;
signal \N__61547\ : std_logic;
signal \N__61546\ : std_logic;
signal \N__61545\ : std_logic;
signal \N__61544\ : std_logic;
signal \N__61541\ : std_logic;
signal \N__61538\ : std_logic;
signal \N__61535\ : std_logic;
signal \N__61532\ : std_logic;
signal \N__61531\ : std_logic;
signal \N__61530\ : std_logic;
signal \N__61527\ : std_logic;
signal \N__61526\ : std_logic;
signal \N__61525\ : std_logic;
signal \N__61522\ : std_logic;
signal \N__61517\ : std_logic;
signal \N__61514\ : std_logic;
signal \N__61511\ : std_logic;
signal \N__61508\ : std_logic;
signal \N__61505\ : std_logic;
signal \N__61502\ : std_logic;
signal \N__61499\ : std_logic;
signal \N__61494\ : std_logic;
signal \N__61491\ : std_logic;
signal \N__61486\ : std_logic;
signal \N__61483\ : std_logic;
signal \N__61478\ : std_logic;
signal \N__61473\ : std_logic;
signal \N__61468\ : std_logic;
signal \N__61461\ : std_logic;
signal \N__61458\ : std_logic;
signal \N__61455\ : std_logic;
signal \N__61452\ : std_logic;
signal \N__61449\ : std_logic;
signal \N__61448\ : std_logic;
signal \N__61447\ : std_logic;
signal \N__61444\ : std_logic;
signal \N__61441\ : std_logic;
signal \N__61438\ : std_logic;
signal \N__61437\ : std_logic;
signal \N__61436\ : std_logic;
signal \N__61435\ : std_logic;
signal \N__61434\ : std_logic;
signal \N__61431\ : std_logic;
signal \N__61428\ : std_logic;
signal \N__61425\ : std_logic;
signal \N__61422\ : std_logic;
signal \N__61421\ : std_logic;
signal \N__61418\ : std_logic;
signal \N__61415\ : std_logic;
signal \N__61412\ : std_logic;
signal \N__61407\ : std_logic;
signal \N__61406\ : std_logic;
signal \N__61401\ : std_logic;
signal \N__61398\ : std_logic;
signal \N__61395\ : std_logic;
signal \N__61390\ : std_logic;
signal \N__61387\ : std_logic;
signal \N__61384\ : std_logic;
signal \N__61381\ : std_logic;
signal \N__61376\ : std_logic;
signal \N__61371\ : std_logic;
signal \N__61362\ : std_logic;
signal \N__61359\ : std_logic;
signal \N__61356\ : std_logic;
signal \N__61355\ : std_logic;
signal \N__61354\ : std_logic;
signal \N__61353\ : std_logic;
signal \N__61352\ : std_logic;
signal \N__61349\ : std_logic;
signal \N__61348\ : std_logic;
signal \N__61345\ : std_logic;
signal \N__61342\ : std_logic;
signal \N__61339\ : std_logic;
signal \N__61336\ : std_logic;
signal \N__61333\ : std_logic;
signal \N__61330\ : std_logic;
signal \N__61327\ : std_logic;
signal \N__61320\ : std_logic;
signal \N__61319\ : std_logic;
signal \N__61318\ : std_logic;
signal \N__61311\ : std_logic;
signal \N__61310\ : std_logic;
signal \N__61307\ : std_logic;
signal \N__61304\ : std_logic;
signal \N__61301\ : std_logic;
signal \N__61298\ : std_logic;
signal \N__61295\ : std_logic;
signal \N__61290\ : std_logic;
signal \N__61287\ : std_logic;
signal \N__61284\ : std_logic;
signal \N__61281\ : std_logic;
signal \N__61276\ : std_logic;
signal \N__61273\ : std_logic;
signal \N__61270\ : std_logic;
signal \N__61267\ : std_logic;
signal \N__61260\ : std_logic;
signal \N__61257\ : std_logic;
signal \N__61254\ : std_logic;
signal \N__61253\ : std_logic;
signal \N__61252\ : std_logic;
signal \N__61249\ : std_logic;
signal \N__61248\ : std_logic;
signal \N__61247\ : std_logic;
signal \N__61246\ : std_logic;
signal \N__61243\ : std_logic;
signal \N__61242\ : std_logic;
signal \N__61239\ : std_logic;
signal \N__61236\ : std_logic;
signal \N__61233\ : std_logic;
signal \N__61230\ : std_logic;
signal \N__61229\ : std_logic;
signal \N__61226\ : std_logic;
signal \N__61223\ : std_logic;
signal \N__61220\ : std_logic;
signal \N__61217\ : std_logic;
signal \N__61212\ : std_logic;
signal \N__61209\ : std_logic;
signal \N__61206\ : std_logic;
signal \N__61203\ : std_logic;
signal \N__61200\ : std_logic;
signal \N__61197\ : std_logic;
signal \N__61194\ : std_logic;
signal \N__61193\ : std_logic;
signal \N__61188\ : std_logic;
signal \N__61185\ : std_logic;
signal \N__61182\ : std_logic;
signal \N__61177\ : std_logic;
signal \N__61174\ : std_logic;
signal \N__61171\ : std_logic;
signal \N__61166\ : std_logic;
signal \N__61163\ : std_logic;
signal \N__61158\ : std_logic;
signal \N__61155\ : std_logic;
signal \N__61152\ : std_logic;
signal \N__61149\ : std_logic;
signal \N__61146\ : std_logic;
signal \N__61137\ : std_logic;
signal \N__61134\ : std_logic;
signal \N__61131\ : std_logic;
signal \N__61130\ : std_logic;
signal \N__61127\ : std_logic;
signal \N__61126\ : std_logic;
signal \N__61125\ : std_logic;
signal \N__61124\ : std_logic;
signal \N__61121\ : std_logic;
signal \N__61118\ : std_logic;
signal \N__61117\ : std_logic;
signal \N__61114\ : std_logic;
signal \N__61113\ : std_logic;
signal \N__61110\ : std_logic;
signal \N__61107\ : std_logic;
signal \N__61104\ : std_logic;
signal \N__61103\ : std_logic;
signal \N__61100\ : std_logic;
signal \N__61097\ : std_logic;
signal \N__61094\ : std_logic;
signal \N__61091\ : std_logic;
signal \N__61088\ : std_logic;
signal \N__61085\ : std_logic;
signal \N__61082\ : std_logic;
signal \N__61079\ : std_logic;
signal \N__61076\ : std_logic;
signal \N__61073\ : std_logic;
signal \N__61070\ : std_logic;
signal \N__61063\ : std_logic;
signal \N__61060\ : std_logic;
signal \N__61057\ : std_logic;
signal \N__61054\ : std_logic;
signal \N__61051\ : std_logic;
signal \N__61048\ : std_logic;
signal \N__61045\ : std_logic;
signal \N__61038\ : std_logic;
signal \N__61033\ : std_logic;
signal \N__61026\ : std_logic;
signal \N__61023\ : std_logic;
signal \N__61020\ : std_logic;
signal \N__61019\ : std_logic;
signal \N__61018\ : std_logic;
signal \N__61015\ : std_logic;
signal \N__61014\ : std_logic;
signal \N__61013\ : std_logic;
signal \N__61010\ : std_logic;
signal \N__61007\ : std_logic;
signal \N__61004\ : std_logic;
signal \N__61001\ : std_logic;
signal \N__61000\ : std_logic;
signal \N__60997\ : std_logic;
signal \N__60994\ : std_logic;
signal \N__60991\ : std_logic;
signal \N__60988\ : std_logic;
signal \N__60985\ : std_logic;
signal \N__60982\ : std_logic;
signal \N__60981\ : std_logic;
signal \N__60980\ : std_logic;
signal \N__60977\ : std_logic;
signal \N__60972\ : std_logic;
signal \N__60967\ : std_logic;
signal \N__60964\ : std_logic;
signal \N__60961\ : std_logic;
signal \N__60958\ : std_logic;
signal \N__60955\ : std_logic;
signal \N__60952\ : std_logic;
signal \N__60949\ : std_logic;
signal \N__60946\ : std_logic;
signal \N__60939\ : std_logic;
signal \N__60934\ : std_logic;
signal \N__60927\ : std_logic;
signal \N__60924\ : std_logic;
signal \N__60921\ : std_logic;
signal \N__60918\ : std_logic;
signal \N__60915\ : std_logic;
signal \N__60914\ : std_logic;
signal \N__60913\ : std_logic;
signal \N__60912\ : std_logic;
signal \N__60909\ : std_logic;
signal \N__60906\ : std_logic;
signal \N__60905\ : std_logic;
signal \N__60902\ : std_logic;
signal \N__60901\ : std_logic;
signal \N__60898\ : std_logic;
signal \N__60897\ : std_logic;
signal \N__60892\ : std_logic;
signal \N__60889\ : std_logic;
signal \N__60886\ : std_logic;
signal \N__60883\ : std_logic;
signal \N__60880\ : std_logic;
signal \N__60877\ : std_logic;
signal \N__60872\ : std_logic;
signal \N__60869\ : std_logic;
signal \N__60866\ : std_logic;
signal \N__60863\ : std_logic;
signal \N__60860\ : std_logic;
signal \N__60857\ : std_logic;
signal \N__60850\ : std_logic;
signal \N__60849\ : std_logic;
signal \N__60846\ : std_logic;
signal \N__60843\ : std_logic;
signal \N__60840\ : std_logic;
signal \N__60837\ : std_logic;
signal \N__60834\ : std_logic;
signal \N__60829\ : std_logic;
signal \N__60822\ : std_logic;
signal \N__60819\ : std_logic;
signal \N__60816\ : std_logic;
signal \N__60813\ : std_logic;
signal \N__60810\ : std_logic;
signal \N__60807\ : std_logic;
signal \N__60806\ : std_logic;
signal \N__60805\ : std_logic;
signal \N__60802\ : std_logic;
signal \N__60799\ : std_logic;
signal \N__60798\ : std_logic;
signal \N__60797\ : std_logic;
signal \N__60794\ : std_logic;
signal \N__60791\ : std_logic;
signal \N__60788\ : std_logic;
signal \N__60787\ : std_logic;
signal \N__60786\ : std_logic;
signal \N__60783\ : std_logic;
signal \N__60780\ : std_logic;
signal \N__60777\ : std_logic;
signal \N__60776\ : std_logic;
signal \N__60771\ : std_logic;
signal \N__60768\ : std_logic;
signal \N__60765\ : std_logic;
signal \N__60762\ : std_logic;
signal \N__60759\ : std_logic;
signal \N__60756\ : std_logic;
signal \N__60753\ : std_logic;
signal \N__60746\ : std_logic;
signal \N__60743\ : std_logic;
signal \N__60740\ : std_logic;
signal \N__60737\ : std_logic;
signal \N__60734\ : std_logic;
signal \N__60731\ : std_logic;
signal \N__60728\ : std_logic;
signal \N__60723\ : std_logic;
signal \N__60714\ : std_logic;
signal \N__60711\ : std_logic;
signal \N__60710\ : std_logic;
signal \N__60709\ : std_logic;
signal \N__60706\ : std_logic;
signal \N__60703\ : std_logic;
signal \N__60700\ : std_logic;
signal \N__60697\ : std_logic;
signal \N__60694\ : std_logic;
signal \N__60691\ : std_logic;
signal \N__60688\ : std_logic;
signal \N__60683\ : std_logic;
signal \N__60678\ : std_logic;
signal \N__60675\ : std_logic;
signal \N__60672\ : std_logic;
signal \N__60669\ : std_logic;
signal \N__60666\ : std_logic;
signal \N__60663\ : std_logic;
signal \N__60660\ : std_logic;
signal \N__60657\ : std_logic;
signal \N__60654\ : std_logic;
signal \N__60651\ : std_logic;
signal \N__60648\ : std_logic;
signal \N__60645\ : std_logic;
signal \N__60642\ : std_logic;
signal \N__60641\ : std_logic;
signal \N__60640\ : std_logic;
signal \N__60637\ : std_logic;
signal \N__60634\ : std_logic;
signal \N__60631\ : std_logic;
signal \N__60626\ : std_logic;
signal \N__60623\ : std_logic;
signal \N__60618\ : std_logic;
signal \N__60617\ : std_logic;
signal \N__60616\ : std_logic;
signal \N__60615\ : std_logic;
signal \N__60614\ : std_logic;
signal \N__60613\ : std_logic;
signal \N__60612\ : std_logic;
signal \N__60609\ : std_logic;
signal \N__60606\ : std_logic;
signal \N__60605\ : std_logic;
signal \N__60604\ : std_logic;
signal \N__60599\ : std_logic;
signal \N__60598\ : std_logic;
signal \N__60597\ : std_logic;
signal \N__60592\ : std_logic;
signal \N__60591\ : std_logic;
signal \N__60590\ : std_logic;
signal \N__60589\ : std_logic;
signal \N__60586\ : std_logic;
signal \N__60581\ : std_logic;
signal \N__60578\ : std_logic;
signal \N__60575\ : std_logic;
signal \N__60572\ : std_logic;
signal \N__60569\ : std_logic;
signal \N__60566\ : std_logic;
signal \N__60565\ : std_logic;
signal \N__60562\ : std_logic;
signal \N__60559\ : std_logic;
signal \N__60558\ : std_logic;
signal \N__60557\ : std_logic;
signal \N__60552\ : std_logic;
signal \N__60549\ : std_logic;
signal \N__60544\ : std_logic;
signal \N__60541\ : std_logic;
signal \N__60540\ : std_logic;
signal \N__60535\ : std_logic;
signal \N__60532\ : std_logic;
signal \N__60529\ : std_logic;
signal \N__60524\ : std_logic;
signal \N__60521\ : std_logic;
signal \N__60518\ : std_logic;
signal \N__60517\ : std_logic;
signal \N__60516\ : std_logic;
signal \N__60515\ : std_logic;
signal \N__60512\ : std_logic;
signal \N__60507\ : std_logic;
signal \N__60504\ : std_logic;
signal \N__60501\ : std_logic;
signal \N__60496\ : std_logic;
signal \N__60489\ : std_logic;
signal \N__60486\ : std_logic;
signal \N__60483\ : std_logic;
signal \N__60478\ : std_logic;
signal \N__60475\ : std_logic;
signal \N__60474\ : std_logic;
signal \N__60473\ : std_logic;
signal \N__60472\ : std_logic;
signal \N__60469\ : std_logic;
signal \N__60464\ : std_logic;
signal \N__60461\ : std_logic;
signal \N__60456\ : std_logic;
signal \N__60451\ : std_logic;
signal \N__60448\ : std_logic;
signal \N__60445\ : std_logic;
signal \N__60440\ : std_logic;
signal \N__60435\ : std_logic;
signal \N__60430\ : std_logic;
signal \N__60427\ : std_logic;
signal \N__60420\ : std_logic;
signal \N__60411\ : std_logic;
signal \N__60408\ : std_logic;
signal \N__60405\ : std_logic;
signal \N__60402\ : std_logic;
signal \N__60399\ : std_logic;
signal \N__60396\ : std_logic;
signal \N__60393\ : std_logic;
signal \N__60390\ : std_logic;
signal \N__60387\ : std_logic;
signal \N__60386\ : std_logic;
signal \N__60385\ : std_logic;
signal \N__60384\ : std_logic;
signal \N__60383\ : std_logic;
signal \N__60382\ : std_logic;
signal \N__60381\ : std_logic;
signal \N__60380\ : std_logic;
signal \N__60379\ : std_logic;
signal \N__60378\ : std_logic;
signal \N__60377\ : std_logic;
signal \N__60376\ : std_logic;
signal \N__60375\ : std_logic;
signal \N__60374\ : std_logic;
signal \N__60369\ : std_logic;
signal \N__60364\ : std_logic;
signal \N__60359\ : std_logic;
signal \N__60358\ : std_logic;
signal \N__60357\ : std_logic;
signal \N__60356\ : std_logic;
signal \N__60355\ : std_logic;
signal \N__60354\ : std_logic;
signal \N__60353\ : std_logic;
signal \N__60350\ : std_logic;
signal \N__60347\ : std_logic;
signal \N__60346\ : std_logic;
signal \N__60345\ : std_logic;
signal \N__60340\ : std_logic;
signal \N__60335\ : std_logic;
signal \N__60330\ : std_logic;
signal \N__60329\ : std_logic;
signal \N__60328\ : std_logic;
signal \N__60325\ : std_logic;
signal \N__60320\ : std_logic;
signal \N__60317\ : std_logic;
signal \N__60312\ : std_logic;
signal \N__60307\ : std_logic;
signal \N__60304\ : std_logic;
signal \N__60299\ : std_logic;
signal \N__60294\ : std_logic;
signal \N__60287\ : std_logic;
signal \N__60282\ : std_logic;
signal \N__60277\ : std_logic;
signal \N__60272\ : std_logic;
signal \N__60269\ : std_logic;
signal \N__60266\ : std_logic;
signal \N__60263\ : std_logic;
signal \N__60260\ : std_logic;
signal \N__60257\ : std_logic;
signal \N__60254\ : std_logic;
signal \N__60249\ : std_logic;
signal \N__60246\ : std_logic;
signal \N__60243\ : std_logic;
signal \N__60240\ : std_logic;
signal \N__60235\ : std_logic;
signal \N__60230\ : std_logic;
signal \N__60219\ : std_logic;
signal \N__60216\ : std_logic;
signal \N__60213\ : std_logic;
signal \N__60210\ : std_logic;
signal \N__60207\ : std_logic;
signal \N__60206\ : std_logic;
signal \N__60205\ : std_logic;
signal \N__60204\ : std_logic;
signal \N__60203\ : std_logic;
signal \N__60202\ : std_logic;
signal \N__60197\ : std_logic;
signal \N__60196\ : std_logic;
signal \N__60195\ : std_logic;
signal \N__60194\ : std_logic;
signal \N__60193\ : std_logic;
signal \N__60188\ : std_logic;
signal \N__60187\ : std_logic;
signal \N__60186\ : std_logic;
signal \N__60181\ : std_logic;
signal \N__60178\ : std_logic;
signal \N__60173\ : std_logic;
signal \N__60168\ : std_logic;
signal \N__60167\ : std_logic;
signal \N__60166\ : std_logic;
signal \N__60165\ : std_logic;
signal \N__60164\ : std_logic;
signal \N__60163\ : std_logic;
signal \N__60162\ : std_logic;
signal \N__60159\ : std_logic;
signal \N__60158\ : std_logic;
signal \N__60157\ : std_logic;
signal \N__60152\ : std_logic;
signal \N__60151\ : std_logic;
signal \N__60150\ : std_logic;
signal \N__60149\ : std_logic;
signal \N__60148\ : std_logic;
signal \N__60145\ : std_logic;
signal \N__60138\ : std_logic;
signal \N__60133\ : std_logic;
signal \N__60128\ : std_logic;
signal \N__60127\ : std_logic;
signal \N__60122\ : std_logic;
signal \N__60119\ : std_logic;
signal \N__60114\ : std_logic;
signal \N__60111\ : std_logic;
signal \N__60106\ : std_logic;
signal \N__60101\ : std_logic;
signal \N__60098\ : std_logic;
signal \N__60093\ : std_logic;
signal \N__60090\ : std_logic;
signal \N__60087\ : std_logic;
signal \N__60084\ : std_logic;
signal \N__60081\ : std_logic;
signal \N__60078\ : std_logic;
signal \N__60073\ : std_logic;
signal \N__60070\ : std_logic;
signal \N__60063\ : std_logic;
signal \N__60060\ : std_logic;
signal \N__60057\ : std_logic;
signal \N__60054\ : std_logic;
signal \N__60051\ : std_logic;
signal \N__60046\ : std_logic;
signal \N__60041\ : std_logic;
signal \N__60030\ : std_logic;
signal \N__60027\ : std_logic;
signal \N__60024\ : std_logic;
signal \N__60023\ : std_logic;
signal \N__60022\ : std_logic;
signal \N__60019\ : std_logic;
signal \N__60018\ : std_logic;
signal \N__60017\ : std_logic;
signal \N__60016\ : std_logic;
signal \N__60013\ : std_logic;
signal \N__60010\ : std_logic;
signal \N__60009\ : std_logic;
signal \N__60006\ : std_logic;
signal \N__60005\ : std_logic;
signal \N__60004\ : std_logic;
signal \N__60001\ : std_logic;
signal \N__59998\ : std_logic;
signal \N__59995\ : std_logic;
signal \N__59994\ : std_logic;
signal \N__59991\ : std_logic;
signal \N__59988\ : std_logic;
signal \N__59985\ : std_logic;
signal \N__59984\ : std_logic;
signal \N__59981\ : std_logic;
signal \N__59978\ : std_logic;
signal \N__59975\ : std_logic;
signal \N__59972\ : std_logic;
signal \N__59969\ : std_logic;
signal \N__59966\ : std_logic;
signal \N__59963\ : std_logic;
signal \N__59958\ : std_logic;
signal \N__59955\ : std_logic;
signal \N__59952\ : std_logic;
signal \N__59947\ : std_logic;
signal \N__59944\ : std_logic;
signal \N__59941\ : std_logic;
signal \N__59940\ : std_logic;
signal \N__59935\ : std_logic;
signal \N__59932\ : std_logic;
signal \N__59929\ : std_logic;
signal \N__59926\ : std_logic;
signal \N__59923\ : std_logic;
signal \N__59920\ : std_logic;
signal \N__59917\ : std_logic;
signal \N__59914\ : std_logic;
signal \N__59911\ : std_logic;
signal \N__59906\ : std_logic;
signal \N__59901\ : std_logic;
signal \N__59896\ : std_logic;
signal \N__59893\ : std_logic;
signal \N__59888\ : std_logic;
signal \N__59885\ : std_logic;
signal \N__59882\ : std_logic;
signal \N__59879\ : std_logic;
signal \N__59874\ : std_logic;
signal \N__59865\ : std_logic;
signal \N__59864\ : std_logic;
signal \N__59863\ : std_logic;
signal \N__59860\ : std_logic;
signal \N__59857\ : std_logic;
signal \N__59854\ : std_logic;
signal \N__59853\ : std_logic;
signal \N__59852\ : std_logic;
signal \N__59851\ : std_logic;
signal \N__59850\ : std_logic;
signal \N__59845\ : std_logic;
signal \N__59844\ : std_logic;
signal \N__59841\ : std_logic;
signal \N__59838\ : std_logic;
signal \N__59835\ : std_logic;
signal \N__59834\ : std_logic;
signal \N__59831\ : std_logic;
signal \N__59828\ : std_logic;
signal \N__59825\ : std_logic;
signal \N__59822\ : std_logic;
signal \N__59817\ : std_logic;
signal \N__59814\ : std_logic;
signal \N__59811\ : std_logic;
signal \N__59808\ : std_logic;
signal \N__59805\ : std_logic;
signal \N__59802\ : std_logic;
signal \N__59797\ : std_logic;
signal \N__59794\ : std_logic;
signal \N__59791\ : std_logic;
signal \N__59788\ : std_logic;
signal \N__59783\ : std_logic;
signal \N__59780\ : std_logic;
signal \N__59775\ : std_logic;
signal \N__59772\ : std_logic;
signal \N__59763\ : std_logic;
signal \N__59760\ : std_logic;
signal \N__59757\ : std_logic;
signal \N__59754\ : std_logic;
signal \N__59751\ : std_logic;
signal \N__59748\ : std_logic;
signal \N__59745\ : std_logic;
signal \N__59742\ : std_logic;
signal \N__59739\ : std_logic;
signal \N__59736\ : std_logic;
signal \N__59733\ : std_logic;
signal \N__59730\ : std_logic;
signal \N__59729\ : std_logic;
signal \N__59728\ : std_logic;
signal \N__59727\ : std_logic;
signal \N__59726\ : std_logic;
signal \N__59723\ : std_logic;
signal \N__59720\ : std_logic;
signal \N__59719\ : std_logic;
signal \N__59718\ : std_logic;
signal \N__59717\ : std_logic;
signal \N__59716\ : std_logic;
signal \N__59715\ : std_logic;
signal \N__59714\ : std_logic;
signal \N__59713\ : std_logic;
signal \N__59712\ : std_logic;
signal \N__59711\ : std_logic;
signal \N__59710\ : std_logic;
signal \N__59709\ : std_logic;
signal \N__59708\ : std_logic;
signal \N__59707\ : std_logic;
signal \N__59706\ : std_logic;
signal \N__59705\ : std_logic;
signal \N__59704\ : std_logic;
signal \N__59703\ : std_logic;
signal \N__59702\ : std_logic;
signal \N__59699\ : std_logic;
signal \N__59698\ : std_logic;
signal \N__59697\ : std_logic;
signal \N__59696\ : std_logic;
signal \N__59695\ : std_logic;
signal \N__59690\ : std_logic;
signal \N__59677\ : std_logic;
signal \N__59676\ : std_logic;
signal \N__59675\ : std_logic;
signal \N__59674\ : std_logic;
signal \N__59673\ : std_logic;
signal \N__59672\ : std_logic;
signal \N__59671\ : std_logic;
signal \N__59654\ : std_logic;
signal \N__59653\ : std_logic;
signal \N__59652\ : std_logic;
signal \N__59651\ : std_logic;
signal \N__59650\ : std_logic;
signal \N__59649\ : std_logic;
signal \N__59648\ : std_logic;
signal \N__59647\ : std_logic;
signal \N__59646\ : std_logic;
signal \N__59645\ : std_logic;
signal \N__59644\ : std_logic;
signal \N__59643\ : std_logic;
signal \N__59642\ : std_logic;
signal \N__59641\ : std_logic;
signal \N__59640\ : std_logic;
signal \N__59639\ : std_logic;
signal \N__59638\ : std_logic;
signal \N__59637\ : std_logic;
signal \N__59636\ : std_logic;
signal \N__59635\ : std_logic;
signal \N__59634\ : std_logic;
signal \N__59633\ : std_logic;
signal \N__59632\ : std_logic;
signal \N__59625\ : std_logic;
signal \N__59608\ : std_logic;
signal \N__59607\ : std_logic;
signal \N__59606\ : std_logic;
signal \N__59605\ : std_logic;
signal \N__59604\ : std_logic;
signal \N__59603\ : std_logic;
signal \N__59602\ : std_logic;
signal \N__59601\ : std_logic;
signal \N__59600\ : std_logic;
signal \N__59599\ : std_logic;
signal \N__59598\ : std_logic;
signal \N__59597\ : std_logic;
signal \N__59596\ : std_logic;
signal \N__59595\ : std_logic;
signal \N__59594\ : std_logic;
signal \N__59593\ : std_logic;
signal \N__59592\ : std_logic;
signal \N__59591\ : std_logic;
signal \N__59590\ : std_logic;
signal \N__59589\ : std_logic;
signal \N__59588\ : std_logic;
signal \N__59587\ : std_logic;
signal \N__59582\ : std_logic;
signal \N__59569\ : std_logic;
signal \N__59566\ : std_logic;
signal \N__59559\ : std_logic;
signal \N__59558\ : std_logic;
signal \N__59557\ : std_logic;
signal \N__59556\ : std_logic;
signal \N__59555\ : std_logic;
signal \N__59554\ : std_logic;
signal \N__59553\ : std_logic;
signal \N__59552\ : std_logic;
signal \N__59551\ : std_logic;
signal \N__59550\ : std_logic;
signal \N__59549\ : std_logic;
signal \N__59548\ : std_logic;
signal \N__59547\ : std_logic;
signal \N__59546\ : std_logic;
signal \N__59545\ : std_logic;
signal \N__59544\ : std_logic;
signal \N__59543\ : std_logic;
signal \N__59542\ : std_logic;
signal \N__59541\ : std_logic;
signal \N__59524\ : std_logic;
signal \N__59517\ : std_logic;
signal \N__59516\ : std_logic;
signal \N__59515\ : std_logic;
signal \N__59514\ : std_logic;
signal \N__59513\ : std_logic;
signal \N__59512\ : std_logic;
signal \N__59511\ : std_logic;
signal \N__59510\ : std_logic;
signal \N__59509\ : std_logic;
signal \N__59508\ : std_logic;
signal \N__59507\ : std_logic;
signal \N__59506\ : std_logic;
signal \N__59505\ : std_logic;
signal \N__59504\ : std_logic;
signal \N__59487\ : std_logic;
signal \N__59482\ : std_logic;
signal \N__59465\ : std_logic;
signal \N__59460\ : std_logic;
signal \N__59449\ : std_logic;
signal \N__59448\ : std_logic;
signal \N__59447\ : std_logic;
signal \N__59446\ : std_logic;
signal \N__59445\ : std_logic;
signal \N__59444\ : std_logic;
signal \N__59443\ : std_logic;
signal \N__59442\ : std_logic;
signal \N__59441\ : std_logic;
signal \N__59440\ : std_logic;
signal \N__59439\ : std_logic;
signal \N__59438\ : std_logic;
signal \N__59437\ : std_logic;
signal \N__59436\ : std_logic;
signal \N__59435\ : std_logic;
signal \N__59434\ : std_logic;
signal \N__59433\ : std_logic;
signal \N__59432\ : std_logic;
signal \N__59431\ : std_logic;
signal \N__59430\ : std_logic;
signal \N__59429\ : std_logic;
signal \N__59428\ : std_logic;
signal \N__59427\ : std_logic;
signal \N__59426\ : std_logic;
signal \N__59425\ : std_logic;
signal \N__59424\ : std_logic;
signal \N__59423\ : std_logic;
signal \N__59422\ : std_logic;
signal \N__59421\ : std_logic;
signal \N__59420\ : std_logic;
signal \N__59419\ : std_logic;
signal \N__59418\ : std_logic;
signal \N__59417\ : std_logic;
signal \N__59416\ : std_logic;
signal \N__59415\ : std_logic;
signal \N__59414\ : std_logic;
signal \N__59413\ : std_logic;
signal \N__59412\ : std_logic;
signal \N__59399\ : std_logic;
signal \N__59394\ : std_logic;
signal \N__59389\ : std_logic;
signal \N__59388\ : std_logic;
signal \N__59387\ : std_logic;
signal \N__59386\ : std_logic;
signal \N__59385\ : std_logic;
signal \N__59384\ : std_logic;
signal \N__59383\ : std_logic;
signal \N__59382\ : std_logic;
signal \N__59381\ : std_logic;
signal \N__59374\ : std_logic;
signal \N__59371\ : std_logic;
signal \N__59368\ : std_logic;
signal \N__59365\ : std_logic;
signal \N__59348\ : std_logic;
signal \N__59345\ : std_logic;
signal \N__59342\ : std_logic;
signal \N__59339\ : std_logic;
signal \N__59336\ : std_logic;
signal \N__59335\ : std_logic;
signal \N__59334\ : std_logic;
signal \N__59333\ : std_logic;
signal \N__59328\ : std_logic;
signal \N__59311\ : std_logic;
signal \N__59308\ : std_logic;
signal \N__59299\ : std_logic;
signal \N__59294\ : std_logic;
signal \N__59287\ : std_logic;
signal \N__59284\ : std_logic;
signal \N__59281\ : std_logic;
signal \N__59278\ : std_logic;
signal \N__59277\ : std_logic;
signal \N__59276\ : std_logic;
signal \N__59275\ : std_logic;
signal \N__59272\ : std_logic;
signal \N__59269\ : std_logic;
signal \N__59262\ : std_logic;
signal \N__59245\ : std_logic;
signal \N__59240\ : std_logic;
signal \N__59223\ : std_logic;
signal \N__59216\ : std_logic;
signal \N__59199\ : std_logic;
signal \N__59194\ : std_logic;
signal \N__59191\ : std_logic;
signal \N__59190\ : std_logic;
signal \N__59189\ : std_logic;
signal \N__59188\ : std_logic;
signal \N__59187\ : std_logic;
signal \N__59186\ : std_logic;
signal \N__59185\ : std_logic;
signal \N__59184\ : std_logic;
signal \N__59183\ : std_logic;
signal \N__59180\ : std_logic;
signal \N__59171\ : std_logic;
signal \N__59166\ : std_logic;
signal \N__59165\ : std_logic;
signal \N__59164\ : std_logic;
signal \N__59163\ : std_logic;
signal \N__59162\ : std_logic;
signal \N__59161\ : std_logic;
signal \N__59160\ : std_logic;
signal \N__59157\ : std_logic;
signal \N__59150\ : std_logic;
signal \N__59149\ : std_logic;
signal \N__59148\ : std_logic;
signal \N__59147\ : std_logic;
signal \N__59146\ : std_logic;
signal \N__59145\ : std_logic;
signal \N__59144\ : std_logic;
signal \N__59143\ : std_logic;
signal \N__59142\ : std_logic;
signal \N__59141\ : std_logic;
signal \N__59140\ : std_logic;
signal \N__59139\ : std_logic;
signal \N__59134\ : std_logic;
signal \N__59119\ : std_logic;
signal \N__59106\ : std_logic;
signal \N__59093\ : std_logic;
signal \N__59090\ : std_logic;
signal \N__59085\ : std_logic;
signal \N__59082\ : std_logic;
signal \N__59071\ : std_logic;
signal \N__59068\ : std_logic;
signal \N__59051\ : std_logic;
signal \N__59046\ : std_logic;
signal \N__59043\ : std_logic;
signal \N__59038\ : std_logic;
signal \N__59035\ : std_logic;
signal \N__59032\ : std_logic;
signal \N__59029\ : std_logic;
signal \N__59026\ : std_logic;
signal \N__59025\ : std_logic;
signal \N__59024\ : std_logic;
signal \N__59023\ : std_logic;
signal \N__59020\ : std_logic;
signal \N__59017\ : std_logic;
signal \N__59016\ : std_logic;
signal \N__59015\ : std_logic;
signal \N__59014\ : std_logic;
signal \N__59013\ : std_logic;
signal \N__59012\ : std_logic;
signal \N__59011\ : std_logic;
signal \N__59010\ : std_logic;
signal \N__58993\ : std_logic;
signal \N__58988\ : std_logic;
signal \N__58985\ : std_logic;
signal \N__58978\ : std_logic;
signal \N__58971\ : std_logic;
signal \N__58964\ : std_logic;
signal \N__58955\ : std_logic;
signal \N__58940\ : std_logic;
signal \N__58935\ : std_logic;
signal \N__58926\ : std_logic;
signal \N__58919\ : std_logic;
signal \N__58916\ : std_logic;
signal \N__58909\ : std_logic;
signal \N__58902\ : std_logic;
signal \N__58897\ : std_logic;
signal \N__58884\ : std_logic;
signal \N__58881\ : std_logic;
signal \N__58880\ : std_logic;
signal \N__58879\ : std_logic;
signal \N__58876\ : std_logic;
signal \N__58873\ : std_logic;
signal \N__58870\ : std_logic;
signal \N__58869\ : std_logic;
signal \N__58868\ : std_logic;
signal \N__58867\ : std_logic;
signal \N__58862\ : std_logic;
signal \N__58859\ : std_logic;
signal \N__58856\ : std_logic;
signal \N__58853\ : std_logic;
signal \N__58850\ : std_logic;
signal \N__58843\ : std_logic;
signal \N__58840\ : std_logic;
signal \N__58837\ : std_logic;
signal \N__58834\ : std_logic;
signal \N__58831\ : std_logic;
signal \N__58828\ : std_logic;
signal \N__58825\ : std_logic;
signal \N__58818\ : std_logic;
signal \N__58815\ : std_logic;
signal \N__58812\ : std_logic;
signal \N__58809\ : std_logic;
signal \N__58806\ : std_logic;
signal \N__58803\ : std_logic;
signal \N__58800\ : std_logic;
signal \N__58797\ : std_logic;
signal \N__58796\ : std_logic;
signal \N__58795\ : std_logic;
signal \N__58792\ : std_logic;
signal \N__58789\ : std_logic;
signal \N__58788\ : std_logic;
signal \N__58787\ : std_logic;
signal \N__58784\ : std_logic;
signal \N__58783\ : std_logic;
signal \N__58780\ : std_logic;
signal \N__58779\ : std_logic;
signal \N__58776\ : std_logic;
signal \N__58773\ : std_logic;
signal \N__58770\ : std_logic;
signal \N__58767\ : std_logic;
signal \N__58766\ : std_logic;
signal \N__58763\ : std_logic;
signal \N__58760\ : std_logic;
signal \N__58757\ : std_logic;
signal \N__58750\ : std_logic;
signal \N__58749\ : std_logic;
signal \N__58746\ : std_logic;
signal \N__58743\ : std_logic;
signal \N__58738\ : std_logic;
signal \N__58733\ : std_logic;
signal \N__58730\ : std_logic;
signal \N__58727\ : std_logic;
signal \N__58724\ : std_logic;
signal \N__58721\ : std_logic;
signal \N__58716\ : std_logic;
signal \N__58707\ : std_logic;
signal \N__58704\ : std_logic;
signal \N__58701\ : std_logic;
signal \N__58700\ : std_logic;
signal \N__58697\ : std_logic;
signal \N__58696\ : std_logic;
signal \N__58693\ : std_logic;
signal \N__58692\ : std_logic;
signal \N__58691\ : std_logic;
signal \N__58688\ : std_logic;
signal \N__58685\ : std_logic;
signal \N__58684\ : std_logic;
signal \N__58681\ : std_logic;
signal \N__58678\ : std_logic;
signal \N__58675\ : std_logic;
signal \N__58670\ : std_logic;
signal \N__58667\ : std_logic;
signal \N__58666\ : std_logic;
signal \N__58661\ : std_logic;
signal \N__58660\ : std_logic;
signal \N__58657\ : std_logic;
signal \N__58652\ : std_logic;
signal \N__58649\ : std_logic;
signal \N__58646\ : std_logic;
signal \N__58643\ : std_logic;
signal \N__58638\ : std_logic;
signal \N__58635\ : std_logic;
signal \N__58634\ : std_logic;
signal \N__58629\ : std_logic;
signal \N__58626\ : std_logic;
signal \N__58623\ : std_logic;
signal \N__58620\ : std_logic;
signal \N__58617\ : std_logic;
signal \N__58612\ : std_logic;
signal \N__58609\ : std_logic;
signal \N__58602\ : std_logic;
signal \N__58599\ : std_logic;
signal \N__58596\ : std_logic;
signal \N__58595\ : std_logic;
signal \N__58594\ : std_logic;
signal \N__58593\ : std_logic;
signal \N__58592\ : std_logic;
signal \N__58591\ : std_logic;
signal \N__58590\ : std_logic;
signal \N__58589\ : std_logic;
signal \N__58586\ : std_logic;
signal \N__58583\ : std_logic;
signal \N__58580\ : std_logic;
signal \N__58577\ : std_logic;
signal \N__58574\ : std_logic;
signal \N__58571\ : std_logic;
signal \N__58568\ : std_logic;
signal \N__58565\ : std_logic;
signal \N__58562\ : std_logic;
signal \N__58561\ : std_logic;
signal \N__58556\ : std_logic;
signal \N__58553\ : std_logic;
signal \N__58550\ : std_logic;
signal \N__58545\ : std_logic;
signal \N__58540\ : std_logic;
signal \N__58537\ : std_logic;
signal \N__58534\ : std_logic;
signal \N__58531\ : std_logic;
signal \N__58524\ : std_logic;
signal \N__58521\ : std_logic;
signal \N__58518\ : std_logic;
signal \N__58515\ : std_logic;
signal \N__58512\ : std_logic;
signal \N__58509\ : std_logic;
signal \N__58500\ : std_logic;
signal \N__58499\ : std_logic;
signal \N__58498\ : std_logic;
signal \N__58497\ : std_logic;
signal \N__58496\ : std_logic;
signal \N__58493\ : std_logic;
signal \N__58490\ : std_logic;
signal \N__58489\ : std_logic;
signal \N__58486\ : std_logic;
signal \N__58483\ : std_logic;
signal \N__58480\ : std_logic;
signal \N__58477\ : std_logic;
signal \N__58474\ : std_logic;
signal \N__58473\ : std_logic;
signal \N__58470\ : std_logic;
signal \N__58465\ : std_logic;
signal \N__58462\ : std_logic;
signal \N__58459\ : std_logic;
signal \N__58456\ : std_logic;
signal \N__58455\ : std_logic;
signal \N__58452\ : std_logic;
signal \N__58449\ : std_logic;
signal \N__58444\ : std_logic;
signal \N__58441\ : std_logic;
signal \N__58440\ : std_logic;
signal \N__58437\ : std_logic;
signal \N__58434\ : std_logic;
signal \N__58431\ : std_logic;
signal \N__58428\ : std_logic;
signal \N__58425\ : std_logic;
signal \N__58422\ : std_logic;
signal \N__58419\ : std_logic;
signal \N__58416\ : std_logic;
signal \N__58413\ : std_logic;
signal \N__58406\ : std_logic;
signal \N__58403\ : std_logic;
signal \N__58400\ : std_logic;
signal \N__58395\ : std_logic;
signal \N__58386\ : std_logic;
signal \N__58383\ : std_logic;
signal \N__58380\ : std_logic;
signal \N__58377\ : std_logic;
signal \N__58376\ : std_logic;
signal \N__58373\ : std_logic;
signal \N__58370\ : std_logic;
signal \N__58365\ : std_logic;
signal \N__58364\ : std_logic;
signal \N__58361\ : std_logic;
signal \N__58358\ : std_logic;
signal \N__58357\ : std_logic;
signal \N__58352\ : std_logic;
signal \N__58351\ : std_logic;
signal \N__58350\ : std_logic;
signal \N__58349\ : std_logic;
signal \N__58348\ : std_logic;
signal \N__58345\ : std_logic;
signal \N__58342\ : std_logic;
signal \N__58339\ : std_logic;
signal \N__58336\ : std_logic;
signal \N__58333\ : std_logic;
signal \N__58332\ : std_logic;
signal \N__58329\ : std_logic;
signal \N__58326\ : std_logic;
signal \N__58323\ : std_logic;
signal \N__58316\ : std_logic;
signal \N__58313\ : std_logic;
signal \N__58310\ : std_logic;
signal \N__58307\ : std_logic;
signal \N__58302\ : std_logic;
signal \N__58299\ : std_logic;
signal \N__58296\ : std_logic;
signal \N__58293\ : std_logic;
signal \N__58290\ : std_logic;
signal \N__58287\ : std_logic;
signal \N__58284\ : std_logic;
signal \N__58281\ : std_logic;
signal \N__58276\ : std_logic;
signal \N__58269\ : std_logic;
signal \N__58266\ : std_logic;
signal \N__58263\ : std_logic;
signal \N__58260\ : std_logic;
signal \N__58257\ : std_logic;
signal \N__58256\ : std_logic;
signal \N__58253\ : std_logic;
signal \N__58250\ : std_logic;
signal \N__58247\ : std_logic;
signal \N__58246\ : std_logic;
signal \N__58243\ : std_logic;
signal \N__58240\ : std_logic;
signal \N__58237\ : std_logic;
signal \N__58232\ : std_logic;
signal \N__58227\ : std_logic;
signal \N__58224\ : std_logic;
signal \N__58223\ : std_logic;
signal \N__58220\ : std_logic;
signal \N__58217\ : std_logic;
signal \N__58212\ : std_logic;
signal \N__58211\ : std_logic;
signal \N__58208\ : std_logic;
signal \N__58205\ : std_logic;
signal \N__58200\ : std_logic;
signal \N__58199\ : std_logic;
signal \N__58198\ : std_logic;
signal \N__58197\ : std_logic;
signal \N__58196\ : std_logic;
signal \N__58191\ : std_logic;
signal \N__58190\ : std_logic;
signal \N__58187\ : std_logic;
signal \N__58186\ : std_logic;
signal \N__58185\ : std_logic;
signal \N__58184\ : std_logic;
signal \N__58183\ : std_logic;
signal \N__58182\ : std_logic;
signal \N__58181\ : std_logic;
signal \N__58180\ : std_logic;
signal \N__58179\ : std_logic;
signal \N__58174\ : std_logic;
signal \N__58171\ : std_logic;
signal \N__58166\ : std_logic;
signal \N__58165\ : std_logic;
signal \N__58160\ : std_logic;
signal \N__58159\ : std_logic;
signal \N__58158\ : std_logic;
signal \N__58157\ : std_logic;
signal \N__58156\ : std_logic;
signal \N__58153\ : std_logic;
signal \N__58148\ : std_logic;
signal \N__58143\ : std_logic;
signal \N__58140\ : std_logic;
signal \N__58135\ : std_logic;
signal \N__58132\ : std_logic;
signal \N__58129\ : std_logic;
signal \N__58126\ : std_logic;
signal \N__58121\ : std_logic;
signal \N__58120\ : std_logic;
signal \N__58117\ : std_logic;
signal \N__58114\ : std_logic;
signal \N__58113\ : std_logic;
signal \N__58112\ : std_logic;
signal \N__58111\ : std_logic;
signal \N__58110\ : std_logic;
signal \N__58105\ : std_logic;
signal \N__58102\ : std_logic;
signal \N__58099\ : std_logic;
signal \N__58094\ : std_logic;
signal \N__58089\ : std_logic;
signal \N__58086\ : std_logic;
signal \N__58083\ : std_logic;
signal \N__58078\ : std_logic;
signal \N__58073\ : std_logic;
signal \N__58068\ : std_logic;
signal \N__58065\ : std_logic;
signal \N__58060\ : std_logic;
signal \N__58057\ : std_logic;
signal \N__58050\ : std_logic;
signal \N__58045\ : std_logic;
signal \N__58038\ : std_logic;
signal \N__58035\ : std_logic;
signal \N__58032\ : std_logic;
signal \N__58027\ : std_logic;
signal \N__58024\ : std_logic;
signal \N__58017\ : std_logic;
signal \N__58016\ : std_logic;
signal \N__58015\ : std_logic;
signal \N__58014\ : std_logic;
signal \N__58013\ : std_logic;
signal \N__58008\ : std_logic;
signal \N__58007\ : std_logic;
signal \N__58006\ : std_logic;
signal \N__58005\ : std_logic;
signal \N__58004\ : std_logic;
signal \N__58001\ : std_logic;
signal \N__57996\ : std_logic;
signal \N__57993\ : std_logic;
signal \N__57992\ : std_logic;
signal \N__57991\ : std_logic;
signal \N__57990\ : std_logic;
signal \N__57989\ : std_logic;
signal \N__57988\ : std_logic;
signal \N__57987\ : std_logic;
signal \N__57982\ : std_logic;
signal \N__57981\ : std_logic;
signal \N__57980\ : std_logic;
signal \N__57979\ : std_logic;
signal \N__57978\ : std_logic;
signal \N__57973\ : std_logic;
signal \N__57970\ : std_logic;
signal \N__57967\ : std_logic;
signal \N__57964\ : std_logic;
signal \N__57959\ : std_logic;
signal \N__57954\ : std_logic;
signal \N__57949\ : std_logic;
signal \N__57946\ : std_logic;
signal \N__57943\ : std_logic;
signal \N__57942\ : std_logic;
signal \N__57941\ : std_logic;
signal \N__57936\ : std_logic;
signal \N__57935\ : std_logic;
signal \N__57932\ : std_logic;
signal \N__57927\ : std_logic;
signal \N__57926\ : std_logic;
signal \N__57923\ : std_logic;
signal \N__57918\ : std_logic;
signal \N__57915\ : std_logic;
signal \N__57914\ : std_logic;
signal \N__57911\ : std_logic;
signal \N__57906\ : std_logic;
signal \N__57901\ : std_logic;
signal \N__57898\ : std_logic;
signal \N__57895\ : std_logic;
signal \N__57890\ : std_logic;
signal \N__57887\ : std_logic;
signal \N__57880\ : std_logic;
signal \N__57877\ : std_logic;
signal \N__57872\ : std_logic;
signal \N__57869\ : std_logic;
signal \N__57866\ : std_logic;
signal \N__57861\ : std_logic;
signal \N__57852\ : std_logic;
signal \N__57849\ : std_logic;
signal \N__57846\ : std_logic;
signal \N__57841\ : std_logic;
signal \N__57834\ : std_logic;
signal \N__57833\ : std_logic;
signal \N__57830\ : std_logic;
signal \N__57827\ : std_logic;
signal \N__57826\ : std_logic;
signal \N__57823\ : std_logic;
signal \N__57820\ : std_logic;
signal \N__57817\ : std_logic;
signal \N__57814\ : std_logic;
signal \N__57811\ : std_logic;
signal \N__57808\ : std_logic;
signal \N__57801\ : std_logic;
signal \N__57800\ : std_logic;
signal \N__57799\ : std_logic;
signal \N__57796\ : std_logic;
signal \N__57793\ : std_logic;
signal \N__57790\ : std_logic;
signal \N__57787\ : std_logic;
signal \N__57784\ : std_logic;
signal \N__57781\ : std_logic;
signal \N__57778\ : std_logic;
signal \N__57775\ : std_logic;
signal \N__57772\ : std_logic;
signal \N__57769\ : std_logic;
signal \N__57764\ : std_logic;
signal \N__57761\ : std_logic;
signal \N__57758\ : std_logic;
signal \N__57753\ : std_logic;
signal \N__57750\ : std_logic;
signal \N__57747\ : std_logic;
signal \N__57744\ : std_logic;
signal \N__57743\ : std_logic;
signal \N__57740\ : std_logic;
signal \N__57737\ : std_logic;
signal \N__57736\ : std_logic;
signal \N__57731\ : std_logic;
signal \N__57728\ : std_logic;
signal \N__57723\ : std_logic;
signal \N__57720\ : std_logic;
signal \N__57719\ : std_logic;
signal \N__57718\ : std_logic;
signal \N__57715\ : std_logic;
signal \N__57710\ : std_logic;
signal \N__57705\ : std_logic;
signal \N__57702\ : std_logic;
signal \N__57699\ : std_logic;
signal \N__57696\ : std_logic;
signal \N__57693\ : std_logic;
signal \N__57690\ : std_logic;
signal \N__57687\ : std_logic;
signal \N__57686\ : std_logic;
signal \N__57685\ : std_logic;
signal \N__57682\ : std_logic;
signal \N__57679\ : std_logic;
signal \N__57676\ : std_logic;
signal \N__57671\ : std_logic;
signal \N__57668\ : std_logic;
signal \N__57665\ : std_logic;
signal \N__57662\ : std_logic;
signal \N__57659\ : std_logic;
signal \N__57656\ : std_logic;
signal \N__57653\ : std_logic;
signal \N__57650\ : std_logic;
signal \N__57645\ : std_logic;
signal \N__57642\ : std_logic;
signal \N__57639\ : std_logic;
signal \N__57636\ : std_logic;
signal \N__57633\ : std_logic;
signal \N__57632\ : std_logic;
signal \N__57629\ : std_logic;
signal \N__57628\ : std_logic;
signal \N__57627\ : std_logic;
signal \N__57624\ : std_logic;
signal \N__57621\ : std_logic;
signal \N__57620\ : std_logic;
signal \N__57619\ : std_logic;
signal \N__57618\ : std_logic;
signal \N__57615\ : std_logic;
signal \N__57612\ : std_logic;
signal \N__57609\ : std_logic;
signal \N__57608\ : std_logic;
signal \N__57605\ : std_logic;
signal \N__57602\ : std_logic;
signal \N__57601\ : std_logic;
signal \N__57598\ : std_logic;
signal \N__57595\ : std_logic;
signal \N__57592\ : std_logic;
signal \N__57589\ : std_logic;
signal \N__57586\ : std_logic;
signal \N__57583\ : std_logic;
signal \N__57580\ : std_logic;
signal \N__57577\ : std_logic;
signal \N__57574\ : std_logic;
signal \N__57571\ : std_logic;
signal \N__57568\ : std_logic;
signal \N__57561\ : std_logic;
signal \N__57558\ : std_logic;
signal \N__57555\ : std_logic;
signal \N__57540\ : std_logic;
signal \N__57537\ : std_logic;
signal \N__57536\ : std_logic;
signal \N__57535\ : std_logic;
signal \N__57534\ : std_logic;
signal \N__57531\ : std_logic;
signal \N__57528\ : std_logic;
signal \N__57525\ : std_logic;
signal \N__57524\ : std_logic;
signal \N__57521\ : std_logic;
signal \N__57520\ : std_logic;
signal \N__57513\ : std_logic;
signal \N__57510\ : std_logic;
signal \N__57509\ : std_logic;
signal \N__57506\ : std_logic;
signal \N__57503\ : std_logic;
signal \N__57500\ : std_logic;
signal \N__57497\ : std_logic;
signal \N__57496\ : std_logic;
signal \N__57493\ : std_logic;
signal \N__57490\ : std_logic;
signal \N__57487\ : std_logic;
signal \N__57482\ : std_logic;
signal \N__57479\ : std_logic;
signal \N__57476\ : std_logic;
signal \N__57475\ : std_logic;
signal \N__57472\ : std_logic;
signal \N__57469\ : std_logic;
signal \N__57464\ : std_logic;
signal \N__57461\ : std_logic;
signal \N__57458\ : std_logic;
signal \N__57453\ : std_logic;
signal \N__57450\ : std_logic;
signal \N__57447\ : std_logic;
signal \N__57444\ : std_logic;
signal \N__57435\ : std_logic;
signal \N__57432\ : std_logic;
signal \N__57429\ : std_logic;
signal \N__57426\ : std_logic;
signal \N__57423\ : std_logic;
signal \N__57420\ : std_logic;
signal \N__57419\ : std_logic;
signal \N__57418\ : std_logic;
signal \N__57415\ : std_logic;
signal \N__57414\ : std_logic;
signal \N__57413\ : std_logic;
signal \N__57412\ : std_logic;
signal \N__57409\ : std_logic;
signal \N__57406\ : std_logic;
signal \N__57403\ : std_logic;
signal \N__57400\ : std_logic;
signal \N__57397\ : std_logic;
signal \N__57394\ : std_logic;
signal \N__57393\ : std_logic;
signal \N__57392\ : std_logic;
signal \N__57389\ : std_logic;
signal \N__57386\ : std_logic;
signal \N__57383\ : std_logic;
signal \N__57380\ : std_logic;
signal \N__57375\ : std_logic;
signal \N__57374\ : std_logic;
signal \N__57371\ : std_logic;
signal \N__57368\ : std_logic;
signal \N__57361\ : std_logic;
signal \N__57356\ : std_logic;
signal \N__57353\ : std_logic;
signal \N__57350\ : std_logic;
signal \N__57343\ : std_logic;
signal \N__57340\ : std_logic;
signal \N__57337\ : std_logic;
signal \N__57330\ : std_logic;
signal \N__57327\ : std_logic;
signal \N__57324\ : std_logic;
signal \N__57323\ : std_logic;
signal \N__57320\ : std_logic;
signal \N__57319\ : std_logic;
signal \N__57316\ : std_logic;
signal \N__57313\ : std_logic;
signal \N__57310\ : std_logic;
signal \N__57307\ : std_logic;
signal \N__57300\ : std_logic;
signal \N__57297\ : std_logic;
signal \N__57294\ : std_logic;
signal \N__57291\ : std_logic;
signal \N__57288\ : std_logic;
signal \N__57287\ : std_logic;
signal \N__57284\ : std_logic;
signal \N__57281\ : std_logic;
signal \N__57278\ : std_logic;
signal \N__57275\ : std_logic;
signal \N__57272\ : std_logic;
signal \N__57267\ : std_logic;
signal \N__57264\ : std_logic;
signal \N__57261\ : std_logic;
signal \N__57258\ : std_logic;
signal \N__57255\ : std_logic;
signal \N__57252\ : std_logic;
signal \N__57249\ : std_logic;
signal \N__57248\ : std_logic;
signal \N__57243\ : std_logic;
signal \N__57242\ : std_logic;
signal \N__57239\ : std_logic;
signal \N__57238\ : std_logic;
signal \N__57237\ : std_logic;
signal \N__57234\ : std_logic;
signal \N__57231\ : std_logic;
signal \N__57228\ : std_logic;
signal \N__57227\ : std_logic;
signal \N__57224\ : std_logic;
signal \N__57223\ : std_logic;
signal \N__57220\ : std_logic;
signal \N__57217\ : std_logic;
signal \N__57216\ : std_logic;
signal \N__57213\ : std_logic;
signal \N__57210\ : std_logic;
signal \N__57209\ : std_logic;
signal \N__57208\ : std_logic;
signal \N__57205\ : std_logic;
signal \N__57202\ : std_logic;
signal \N__57197\ : std_logic;
signal \N__57194\ : std_logic;
signal \N__57191\ : std_logic;
signal \N__57188\ : std_logic;
signal \N__57185\ : std_logic;
signal \N__57182\ : std_logic;
signal \N__57179\ : std_logic;
signal \N__57176\ : std_logic;
signal \N__57173\ : std_logic;
signal \N__57170\ : std_logic;
signal \N__57167\ : std_logic;
signal \N__57150\ : std_logic;
signal \N__57147\ : std_logic;
signal \N__57146\ : std_logic;
signal \N__57143\ : std_logic;
signal \N__57138\ : std_logic;
signal \N__57135\ : std_logic;
signal \N__57132\ : std_logic;
signal \N__57131\ : std_logic;
signal \N__57128\ : std_logic;
signal \N__57125\ : std_logic;
signal \N__57124\ : std_logic;
signal \N__57123\ : std_logic;
signal \N__57120\ : std_logic;
signal \N__57117\ : std_logic;
signal \N__57114\ : std_logic;
signal \N__57111\ : std_logic;
signal \N__57104\ : std_logic;
signal \N__57101\ : std_logic;
signal \N__57098\ : std_logic;
signal \N__57093\ : std_logic;
signal \N__57090\ : std_logic;
signal \N__57089\ : std_logic;
signal \N__57086\ : std_logic;
signal \N__57083\ : std_logic;
signal \N__57082\ : std_logic;
signal \N__57079\ : std_logic;
signal \N__57076\ : std_logic;
signal \N__57073\ : std_logic;
signal \N__57066\ : std_logic;
signal \N__57063\ : std_logic;
signal \N__57060\ : std_logic;
signal \N__57057\ : std_logic;
signal \N__57056\ : std_logic;
signal \N__57053\ : std_logic;
signal \N__57050\ : std_logic;
signal \N__57047\ : std_logic;
signal \N__57044\ : std_logic;
signal \N__57041\ : std_logic;
signal \N__57036\ : std_logic;
signal \N__57033\ : std_logic;
signal \N__57030\ : std_logic;
signal \N__57029\ : std_logic;
signal \N__57028\ : std_logic;
signal \N__57023\ : std_logic;
signal \N__57020\ : std_logic;
signal \N__57015\ : std_logic;
signal \N__57014\ : std_logic;
signal \N__57013\ : std_logic;
signal \N__57012\ : std_logic;
signal \N__57009\ : std_logic;
signal \N__57006\ : std_logic;
signal \N__57003\ : std_logic;
signal \N__57002\ : std_logic;
signal \N__56999\ : std_logic;
signal \N__56996\ : std_logic;
signal \N__56995\ : std_logic;
signal \N__56994\ : std_logic;
signal \N__56993\ : std_logic;
signal \N__56990\ : std_logic;
signal \N__56985\ : std_logic;
signal \N__56980\ : std_logic;
signal \N__56973\ : std_logic;
signal \N__56964\ : std_logic;
signal \N__56961\ : std_logic;
signal \N__56958\ : std_logic;
signal \N__56955\ : std_logic;
signal \N__56952\ : std_logic;
signal \N__56949\ : std_logic;
signal \N__56948\ : std_logic;
signal \N__56947\ : std_logic;
signal \N__56946\ : std_logic;
signal \N__56943\ : std_logic;
signal \N__56940\ : std_logic;
signal \N__56935\ : std_logic;
signal \N__56932\ : std_logic;
signal \N__56929\ : std_logic;
signal \N__56926\ : std_logic;
signal \N__56921\ : std_logic;
signal \N__56916\ : std_logic;
signal \N__56915\ : std_logic;
signal \N__56910\ : std_logic;
signal \N__56909\ : std_logic;
signal \N__56908\ : std_logic;
signal \N__56905\ : std_logic;
signal \N__56902\ : std_logic;
signal \N__56899\ : std_logic;
signal \N__56896\ : std_logic;
signal \N__56889\ : std_logic;
signal \N__56886\ : std_logic;
signal \N__56885\ : std_logic;
signal \N__56882\ : std_logic;
signal \N__56879\ : std_logic;
signal \N__56878\ : std_logic;
signal \N__56873\ : std_logic;
signal \N__56870\ : std_logic;
signal \N__56869\ : std_logic;
signal \N__56868\ : std_logic;
signal \N__56863\ : std_logic;
signal \N__56858\ : std_logic;
signal \N__56853\ : std_logic;
signal \N__56850\ : std_logic;
signal \N__56847\ : std_logic;
signal \N__56844\ : std_logic;
signal \N__56843\ : std_logic;
signal \N__56840\ : std_logic;
signal \N__56837\ : std_logic;
signal \N__56834\ : std_logic;
signal \N__56829\ : std_logic;
signal \N__56828\ : std_logic;
signal \N__56825\ : std_logic;
signal \N__56822\ : std_logic;
signal \N__56819\ : std_logic;
signal \N__56818\ : std_logic;
signal \N__56817\ : std_logic;
signal \N__56816\ : std_logic;
signal \N__56815\ : std_logic;
signal \N__56812\ : std_logic;
signal \N__56809\ : std_logic;
signal \N__56806\ : std_logic;
signal \N__56799\ : std_logic;
signal \N__56796\ : std_logic;
signal \N__56787\ : std_logic;
signal \N__56784\ : std_logic;
signal \N__56781\ : std_logic;
signal \N__56778\ : std_logic;
signal \N__56775\ : std_logic;
signal \N__56772\ : std_logic;
signal \N__56771\ : std_logic;
signal \N__56770\ : std_logic;
signal \N__56767\ : std_logic;
signal \N__56762\ : std_logic;
signal \N__56757\ : std_logic;
signal \N__56754\ : std_logic;
signal \N__56751\ : std_logic;
signal \N__56748\ : std_logic;
signal \N__56745\ : std_logic;
signal \N__56742\ : std_logic;
signal \N__56739\ : std_logic;
signal \N__56736\ : std_logic;
signal \N__56733\ : std_logic;
signal \N__56730\ : std_logic;
signal \N__56729\ : std_logic;
signal \N__56728\ : std_logic;
signal \N__56727\ : std_logic;
signal \N__56726\ : std_logic;
signal \N__56725\ : std_logic;
signal \N__56722\ : std_logic;
signal \N__56719\ : std_logic;
signal \N__56718\ : std_logic;
signal \N__56713\ : std_logic;
signal \N__56708\ : std_logic;
signal \N__56705\ : std_logic;
signal \N__56702\ : std_logic;
signal \N__56701\ : std_logic;
signal \N__56700\ : std_logic;
signal \N__56697\ : std_logic;
signal \N__56692\ : std_logic;
signal \N__56687\ : std_logic;
signal \N__56684\ : std_logic;
signal \N__56681\ : std_logic;
signal \N__56670\ : std_logic;
signal \N__56667\ : std_logic;
signal \N__56664\ : std_logic;
signal \N__56661\ : std_logic;
signal \N__56660\ : std_logic;
signal \N__56657\ : std_logic;
signal \N__56654\ : std_logic;
signal \N__56651\ : std_logic;
signal \N__56650\ : std_logic;
signal \N__56649\ : std_logic;
signal \N__56646\ : std_logic;
signal \N__56643\ : std_logic;
signal \N__56638\ : std_logic;
signal \N__56631\ : std_logic;
signal \N__56628\ : std_logic;
signal \N__56627\ : std_logic;
signal \N__56622\ : std_logic;
signal \N__56621\ : std_logic;
signal \N__56620\ : std_logic;
signal \N__56617\ : std_logic;
signal \N__56612\ : std_logic;
signal \N__56607\ : std_logic;
signal \N__56606\ : std_logic;
signal \N__56601\ : std_logic;
signal \N__56598\ : std_logic;
signal \N__56595\ : std_logic;
signal \N__56594\ : std_logic;
signal \N__56593\ : std_logic;
signal \N__56592\ : std_logic;
signal \N__56591\ : std_logic;
signal \N__56588\ : std_logic;
signal \N__56585\ : std_logic;
signal \N__56584\ : std_logic;
signal \N__56583\ : std_logic;
signal \N__56578\ : std_logic;
signal \N__56575\ : std_logic;
signal \N__56574\ : std_logic;
signal \N__56569\ : std_logic;
signal \N__56564\ : std_logic;
signal \N__56561\ : std_logic;
signal \N__56560\ : std_logic;
signal \N__56559\ : std_logic;
signal \N__56554\ : std_logic;
signal \N__56549\ : std_logic;
signal \N__56546\ : std_logic;
signal \N__56543\ : std_logic;
signal \N__56540\ : std_logic;
signal \N__56537\ : std_logic;
signal \N__56534\ : std_logic;
signal \N__56529\ : std_logic;
signal \N__56520\ : std_logic;
signal \N__56517\ : std_logic;
signal \N__56516\ : std_logic;
signal \N__56513\ : std_logic;
signal \N__56512\ : std_logic;
signal \N__56511\ : std_logic;
signal \N__56508\ : std_logic;
signal \N__56505\ : std_logic;
signal \N__56500\ : std_logic;
signal \N__56493\ : std_logic;
signal \N__56490\ : std_logic;
signal \N__56489\ : std_logic;
signal \N__56486\ : std_logic;
signal \N__56483\ : std_logic;
signal \N__56480\ : std_logic;
signal \N__56477\ : std_logic;
signal \N__56472\ : std_logic;
signal \N__56469\ : std_logic;
signal \N__56468\ : std_logic;
signal \N__56465\ : std_logic;
signal \N__56462\ : std_logic;
signal \N__56459\ : std_logic;
signal \N__56456\ : std_logic;
signal \N__56453\ : std_logic;
signal \N__56448\ : std_logic;
signal \N__56447\ : std_logic;
signal \N__56446\ : std_logic;
signal \N__56443\ : std_logic;
signal \N__56442\ : std_logic;
signal \N__56441\ : std_logic;
signal \N__56440\ : std_logic;
signal \N__56439\ : std_logic;
signal \N__56434\ : std_logic;
signal \N__56431\ : std_logic;
signal \N__56428\ : std_logic;
signal \N__56425\ : std_logic;
signal \N__56422\ : std_logic;
signal \N__56419\ : std_logic;
signal \N__56416\ : std_logic;
signal \N__56411\ : std_logic;
signal \N__56408\ : std_logic;
signal \N__56407\ : std_logic;
signal \N__56406\ : std_logic;
signal \N__56403\ : std_logic;
signal \N__56394\ : std_logic;
signal \N__56389\ : std_logic;
signal \N__56384\ : std_logic;
signal \N__56379\ : std_logic;
signal \N__56376\ : std_logic;
signal \N__56373\ : std_logic;
signal \N__56370\ : std_logic;
signal \N__56367\ : std_logic;
signal \N__56364\ : std_logic;
signal \N__56361\ : std_logic;
signal \N__56360\ : std_logic;
signal \N__56359\ : std_logic;
signal \N__56358\ : std_logic;
signal \N__56357\ : std_logic;
signal \N__56354\ : std_logic;
signal \N__56353\ : std_logic;
signal \N__56352\ : std_logic;
signal \N__56351\ : std_logic;
signal \N__56350\ : std_logic;
signal \N__56347\ : std_logic;
signal \N__56340\ : std_logic;
signal \N__56337\ : std_logic;
signal \N__56336\ : std_logic;
signal \N__56333\ : std_logic;
signal \N__56330\ : std_logic;
signal \N__56327\ : std_logic;
signal \N__56324\ : std_logic;
signal \N__56317\ : std_logic;
signal \N__56312\ : std_logic;
signal \N__56309\ : std_logic;
signal \N__56308\ : std_logic;
signal \N__56299\ : std_logic;
signal \N__56296\ : std_logic;
signal \N__56293\ : std_logic;
signal \N__56290\ : std_logic;
signal \N__56283\ : std_logic;
signal \N__56280\ : std_logic;
signal \N__56277\ : std_logic;
signal \N__56274\ : std_logic;
signal \N__56271\ : std_logic;
signal \N__56268\ : std_logic;
signal \N__56265\ : std_logic;
signal \N__56262\ : std_logic;
signal \N__56259\ : std_logic;
signal \N__56256\ : std_logic;
signal \N__56253\ : std_logic;
signal \N__56250\ : std_logic;
signal \N__56249\ : std_logic;
signal \N__56248\ : std_logic;
signal \N__56247\ : std_logic;
signal \N__56246\ : std_logic;
signal \N__56245\ : std_logic;
signal \N__56242\ : std_logic;
signal \N__56239\ : std_logic;
signal \N__56236\ : std_logic;
signal \N__56233\ : std_logic;
signal \N__56232\ : std_logic;
signal \N__56229\ : std_logic;
signal \N__56226\ : std_logic;
signal \N__56223\ : std_logic;
signal \N__56216\ : std_logic;
signal \N__56213\ : std_logic;
signal \N__56210\ : std_logic;
signal \N__56207\ : std_logic;
signal \N__56204\ : std_logic;
signal \N__56201\ : std_logic;
signal \N__56198\ : std_logic;
signal \N__56195\ : std_logic;
signal \N__56186\ : std_logic;
signal \N__56181\ : std_logic;
signal \N__56180\ : std_logic;
signal \N__56177\ : std_logic;
signal \N__56174\ : std_logic;
signal \N__56173\ : std_logic;
signal \N__56170\ : std_logic;
signal \N__56167\ : std_logic;
signal \N__56164\ : std_logic;
signal \N__56159\ : std_logic;
signal \N__56154\ : std_logic;
signal \N__56151\ : std_logic;
signal \N__56148\ : std_logic;
signal \N__56147\ : std_logic;
signal \N__56146\ : std_logic;
signal \N__56145\ : std_logic;
signal \N__56144\ : std_logic;
signal \N__56141\ : std_logic;
signal \N__56138\ : std_logic;
signal \N__56131\ : std_logic;
signal \N__56130\ : std_logic;
signal \N__56129\ : std_logic;
signal \N__56128\ : std_logic;
signal \N__56127\ : std_logic;
signal \N__56124\ : std_logic;
signal \N__56123\ : std_logic;
signal \N__56122\ : std_logic;
signal \N__56119\ : std_logic;
signal \N__56116\ : std_logic;
signal \N__56113\ : std_logic;
signal \N__56110\ : std_logic;
signal \N__56105\ : std_logic;
signal \N__56102\ : std_logic;
signal \N__56099\ : std_logic;
signal \N__56096\ : std_logic;
signal \N__56093\ : std_logic;
signal \N__56088\ : std_logic;
signal \N__56081\ : std_logic;
signal \N__56070\ : std_logic;
signal \N__56069\ : std_logic;
signal \N__56066\ : std_logic;
signal \N__56063\ : std_logic;
signal \N__56058\ : std_logic;
signal \N__56057\ : std_logic;
signal \N__56056\ : std_logic;
signal \N__56053\ : std_logic;
signal \N__56050\ : std_logic;
signal \N__56047\ : std_logic;
signal \N__56040\ : std_logic;
signal \N__56037\ : std_logic;
signal \N__56036\ : std_logic;
signal \N__56031\ : std_logic;
signal \N__56028\ : std_logic;
signal \N__56027\ : std_logic;
signal \N__56022\ : std_logic;
signal \N__56019\ : std_logic;
signal \N__56016\ : std_logic;
signal \N__56013\ : std_logic;
signal \N__56010\ : std_logic;
signal \N__56007\ : std_logic;
signal \N__56004\ : std_logic;
signal \N__56001\ : std_logic;
signal \N__55998\ : std_logic;
signal \N__55995\ : std_logic;
signal \N__55992\ : std_logic;
signal \N__55989\ : std_logic;
signal \N__55988\ : std_logic;
signal \N__55983\ : std_logic;
signal \N__55982\ : std_logic;
signal \N__55979\ : std_logic;
signal \N__55976\ : std_logic;
signal \N__55971\ : std_logic;
signal \N__55968\ : std_logic;
signal \N__55965\ : std_logic;
signal \N__55964\ : std_logic;
signal \N__55961\ : std_logic;
signal \N__55960\ : std_logic;
signal \N__55957\ : std_logic;
signal \N__55954\ : std_logic;
signal \N__55951\ : std_logic;
signal \N__55944\ : std_logic;
signal \N__55943\ : std_logic;
signal \N__55940\ : std_logic;
signal \N__55937\ : std_logic;
signal \N__55934\ : std_logic;
signal \N__55929\ : std_logic;
signal \N__55928\ : std_logic;
signal \N__55927\ : std_logic;
signal \N__55924\ : std_logic;
signal \N__55921\ : std_logic;
signal \N__55920\ : std_logic;
signal \N__55917\ : std_logic;
signal \N__55916\ : std_logic;
signal \N__55913\ : std_logic;
signal \N__55910\ : std_logic;
signal \N__55907\ : std_logic;
signal \N__55904\ : std_logic;
signal \N__55901\ : std_logic;
signal \N__55896\ : std_logic;
signal \N__55893\ : std_logic;
signal \N__55890\ : std_logic;
signal \N__55887\ : std_logic;
signal \N__55884\ : std_logic;
signal \N__55875\ : std_logic;
signal \N__55872\ : std_logic;
signal \N__55869\ : std_logic;
signal \N__55868\ : std_logic;
signal \N__55865\ : std_logic;
signal \N__55864\ : std_logic;
signal \N__55863\ : std_logic;
signal \N__55862\ : std_logic;
signal \N__55861\ : std_logic;
signal \N__55858\ : std_logic;
signal \N__55857\ : std_logic;
signal \N__55856\ : std_logic;
signal \N__55855\ : std_logic;
signal \N__55854\ : std_logic;
signal \N__55853\ : std_logic;
signal \N__55850\ : std_logic;
signal \N__55847\ : std_logic;
signal \N__55844\ : std_logic;
signal \N__55841\ : std_logic;
signal \N__55838\ : std_logic;
signal \N__55835\ : std_logic;
signal \N__55824\ : std_logic;
signal \N__55817\ : std_logic;
signal \N__55808\ : std_logic;
signal \N__55805\ : std_logic;
signal \N__55800\ : std_logic;
signal \N__55797\ : std_logic;
signal \N__55796\ : std_logic;
signal \N__55795\ : std_logic;
signal \N__55794\ : std_logic;
signal \N__55791\ : std_logic;
signal \N__55788\ : std_logic;
signal \N__55785\ : std_logic;
signal \N__55782\ : std_logic;
signal \N__55775\ : std_logic;
signal \N__55770\ : std_logic;
signal \N__55767\ : std_logic;
signal \N__55764\ : std_logic;
signal \N__55761\ : std_logic;
signal \N__55758\ : std_logic;
signal \N__55755\ : std_logic;
signal \N__55752\ : std_logic;
signal \N__55749\ : std_logic;
signal \N__55746\ : std_logic;
signal \N__55745\ : std_logic;
signal \N__55744\ : std_logic;
signal \N__55743\ : std_logic;
signal \N__55742\ : std_logic;
signal \N__55741\ : std_logic;
signal \N__55740\ : std_logic;
signal \N__55735\ : std_logic;
signal \N__55728\ : std_logic;
signal \N__55727\ : std_logic;
signal \N__55726\ : std_logic;
signal \N__55725\ : std_logic;
signal \N__55724\ : std_logic;
signal \N__55723\ : std_logic;
signal \N__55722\ : std_logic;
signal \N__55717\ : std_logic;
signal \N__55712\ : std_logic;
signal \N__55707\ : std_logic;
signal \N__55702\ : std_logic;
signal \N__55697\ : std_logic;
signal \N__55696\ : std_logic;
signal \N__55695\ : std_logic;
signal \N__55694\ : std_logic;
signal \N__55693\ : std_logic;
signal \N__55690\ : std_logic;
signal \N__55689\ : std_logic;
signal \N__55688\ : std_logic;
signal \N__55687\ : std_logic;
signal \N__55686\ : std_logic;
signal \N__55683\ : std_logic;
signal \N__55680\ : std_logic;
signal \N__55675\ : std_logic;
signal \N__55670\ : std_logic;
signal \N__55665\ : std_logic;
signal \N__55662\ : std_logic;
signal \N__55653\ : std_logic;
signal \N__55652\ : std_logic;
signal \N__55651\ : std_logic;
signal \N__55650\ : std_logic;
signal \N__55645\ : std_logic;
signal \N__55640\ : std_logic;
signal \N__55637\ : std_logic;
signal \N__55632\ : std_logic;
signal \N__55625\ : std_logic;
signal \N__55622\ : std_logic;
signal \N__55619\ : std_logic;
signal \N__55612\ : std_logic;
signal \N__55609\ : std_logic;
signal \N__55606\ : std_logic;
signal \N__55603\ : std_logic;
signal \N__55596\ : std_logic;
signal \N__55593\ : std_logic;
signal \N__55590\ : std_logic;
signal \N__55587\ : std_logic;
signal \N__55584\ : std_logic;
signal \N__55581\ : std_logic;
signal \N__55578\ : std_logic;
signal \N__55575\ : std_logic;
signal \N__55572\ : std_logic;
signal \N__55571\ : std_logic;
signal \N__55570\ : std_logic;
signal \N__55567\ : std_logic;
signal \N__55564\ : std_logic;
signal \N__55563\ : std_logic;
signal \N__55560\ : std_logic;
signal \N__55559\ : std_logic;
signal \N__55558\ : std_logic;
signal \N__55555\ : std_logic;
signal \N__55552\ : std_logic;
signal \N__55549\ : std_logic;
signal \N__55546\ : std_logic;
signal \N__55543\ : std_logic;
signal \N__55540\ : std_logic;
signal \N__55539\ : std_logic;
signal \N__55538\ : std_logic;
signal \N__55531\ : std_logic;
signal \N__55526\ : std_logic;
signal \N__55523\ : std_logic;
signal \N__55522\ : std_logic;
signal \N__55521\ : std_logic;
signal \N__55518\ : std_logic;
signal \N__55515\ : std_logic;
signal \N__55512\ : std_logic;
signal \N__55507\ : std_logic;
signal \N__55504\ : std_logic;
signal \N__55501\ : std_logic;
signal \N__55498\ : std_logic;
signal \N__55495\ : std_logic;
signal \N__55492\ : std_logic;
signal \N__55489\ : std_logic;
signal \N__55484\ : std_logic;
signal \N__55481\ : std_logic;
signal \N__55478\ : std_logic;
signal \N__55475\ : std_logic;
signal \N__55472\ : std_logic;
signal \N__55467\ : std_logic;
signal \N__55460\ : std_logic;
signal \N__55455\ : std_logic;
signal \N__55454\ : std_logic;
signal \N__55453\ : std_logic;
signal \N__55452\ : std_logic;
signal \N__55451\ : std_logic;
signal \N__55450\ : std_logic;
signal \N__55449\ : std_logic;
signal \N__55448\ : std_logic;
signal \N__55447\ : std_logic;
signal \N__55446\ : std_logic;
signal \N__55445\ : std_logic;
signal \N__55444\ : std_logic;
signal \N__55439\ : std_logic;
signal \N__55438\ : std_logic;
signal \N__55435\ : std_logic;
signal \N__55432\ : std_logic;
signal \N__55431\ : std_logic;
signal \N__55430\ : std_logic;
signal \N__55429\ : std_logic;
signal \N__55428\ : std_logic;
signal \N__55427\ : std_logic;
signal \N__55424\ : std_logic;
signal \N__55423\ : std_logic;
signal \N__55420\ : std_logic;
signal \N__55417\ : std_logic;
signal \N__55410\ : std_logic;
signal \N__55409\ : std_logic;
signal \N__55406\ : std_logic;
signal \N__55403\ : std_logic;
signal \N__55400\ : std_logic;
signal \N__55399\ : std_logic;
signal \N__55396\ : std_logic;
signal \N__55391\ : std_logic;
signal \N__55388\ : std_logic;
signal \N__55387\ : std_logic;
signal \N__55386\ : std_logic;
signal \N__55383\ : std_logic;
signal \N__55376\ : std_logic;
signal \N__55373\ : std_logic;
signal \N__55370\ : std_logic;
signal \N__55367\ : std_logic;
signal \N__55362\ : std_logic;
signal \N__55359\ : std_logic;
signal \N__55352\ : std_logic;
signal \N__55351\ : std_logic;
signal \N__55348\ : std_logic;
signal \N__55345\ : std_logic;
signal \N__55342\ : std_logic;
signal \N__55339\ : std_logic;
signal \N__55336\ : std_logic;
signal \N__55333\ : std_logic;
signal \N__55328\ : std_logic;
signal \N__55319\ : std_logic;
signal \N__55314\ : std_logic;
signal \N__55311\ : std_logic;
signal \N__55306\ : std_logic;
signal \N__55303\ : std_logic;
signal \N__55296\ : std_logic;
signal \N__55291\ : std_logic;
signal \N__55288\ : std_logic;
signal \N__55283\ : std_logic;
signal \N__55278\ : std_logic;
signal \N__55275\ : std_logic;
signal \N__55272\ : std_logic;
signal \N__55263\ : std_logic;
signal \N__55262\ : std_logic;
signal \N__55259\ : std_logic;
signal \N__55258\ : std_logic;
signal \N__55257\ : std_logic;
signal \N__55256\ : std_logic;
signal \N__55255\ : std_logic;
signal \N__55254\ : std_logic;
signal \N__55251\ : std_logic;
signal \N__55250\ : std_logic;
signal \N__55249\ : std_logic;
signal \N__55246\ : std_logic;
signal \N__55239\ : std_logic;
signal \N__55236\ : std_logic;
signal \N__55233\ : std_logic;
signal \N__55232\ : std_logic;
signal \N__55231\ : std_logic;
signal \N__55230\ : std_logic;
signal \N__55229\ : std_logic;
signal \N__55228\ : std_logic;
signal \N__55225\ : std_logic;
signal \N__55222\ : std_logic;
signal \N__55221\ : std_logic;
signal \N__55218\ : std_logic;
signal \N__55217\ : std_logic;
signal \N__55212\ : std_logic;
signal \N__55209\ : std_logic;
signal \N__55206\ : std_logic;
signal \N__55199\ : std_logic;
signal \N__55198\ : std_logic;
signal \N__55193\ : std_logic;
signal \N__55192\ : std_logic;
signal \N__55187\ : std_logic;
signal \N__55184\ : std_logic;
signal \N__55183\ : std_logic;
signal \N__55180\ : std_logic;
signal \N__55177\ : std_logic;
signal \N__55174\ : std_logic;
signal \N__55167\ : std_logic;
signal \N__55164\ : std_logic;
signal \N__55163\ : std_logic;
signal \N__55160\ : std_logic;
signal \N__55157\ : std_logic;
signal \N__55156\ : std_logic;
signal \N__55155\ : std_logic;
signal \N__55154\ : std_logic;
signal \N__55151\ : std_logic;
signal \N__55148\ : std_logic;
signal \N__55145\ : std_logic;
signal \N__55140\ : std_logic;
signal \N__55135\ : std_logic;
signal \N__55132\ : std_logic;
signal \N__55129\ : std_logic;
signal \N__55126\ : std_logic;
signal \N__55123\ : std_logic;
signal \N__55120\ : std_logic;
signal \N__55117\ : std_logic;
signal \N__55114\ : std_logic;
signal \N__55113\ : std_logic;
signal \N__55110\ : std_logic;
signal \N__55105\ : std_logic;
signal \N__55098\ : std_logic;
signal \N__55085\ : std_logic;
signal \N__55082\ : std_logic;
signal \N__55079\ : std_logic;
signal \N__55076\ : std_logic;
signal \N__55069\ : std_logic;
signal \N__55062\ : std_logic;
signal \N__55059\ : std_logic;
signal \N__55058\ : std_logic;
signal \N__55057\ : std_logic;
signal \N__55056\ : std_logic;
signal \N__55055\ : std_logic;
signal \N__55054\ : std_logic;
signal \N__55053\ : std_logic;
signal \N__55052\ : std_logic;
signal \N__55049\ : std_logic;
signal \N__55046\ : std_logic;
signal \N__55043\ : std_logic;
signal \N__55040\ : std_logic;
signal \N__55037\ : std_logic;
signal \N__55036\ : std_logic;
signal \N__55035\ : std_logic;
signal \N__55032\ : std_logic;
signal \N__55031\ : std_logic;
signal \N__55030\ : std_logic;
signal \N__55029\ : std_logic;
signal \N__55026\ : std_logic;
signal \N__55023\ : std_logic;
signal \N__55022\ : std_logic;
signal \N__55021\ : std_logic;
signal \N__55020\ : std_logic;
signal \N__55019\ : std_logic;
signal \N__55014\ : std_logic;
signal \N__55011\ : std_logic;
signal \N__55010\ : std_logic;
signal \N__55005\ : std_logic;
signal \N__55002\ : std_logic;
signal \N__55001\ : std_logic;
signal \N__54998\ : std_logic;
signal \N__54995\ : std_logic;
signal \N__54992\ : std_logic;
signal \N__54989\ : std_logic;
signal \N__54986\ : std_logic;
signal \N__54979\ : std_logic;
signal \N__54976\ : std_logic;
signal \N__54973\ : std_logic;
signal \N__54970\ : std_logic;
signal \N__54967\ : std_logic;
signal \N__54964\ : std_logic;
signal \N__54963\ : std_logic;
signal \N__54960\ : std_logic;
signal \N__54955\ : std_logic;
signal \N__54954\ : std_logic;
signal \N__54953\ : std_logic;
signal \N__54950\ : std_logic;
signal \N__54947\ : std_logic;
signal \N__54944\ : std_logic;
signal \N__54939\ : std_logic;
signal \N__54930\ : std_logic;
signal \N__54929\ : std_logic;
signal \N__54928\ : std_logic;
signal \N__54925\ : std_logic;
signal \N__54920\ : std_logic;
signal \N__54917\ : std_logic;
signal \N__54914\ : std_logic;
signal \N__54911\ : std_logic;
signal \N__54908\ : std_logic;
signal \N__54905\ : std_logic;
signal \N__54902\ : std_logic;
signal \N__54893\ : std_logic;
signal \N__54888\ : std_logic;
signal \N__54885\ : std_logic;
signal \N__54882\ : std_logic;
signal \N__54879\ : std_logic;
signal \N__54874\ : std_logic;
signal \N__54871\ : std_logic;
signal \N__54862\ : std_logic;
signal \N__54859\ : std_logic;
signal \N__54854\ : std_logic;
signal \N__54851\ : std_logic;
signal \N__54846\ : std_logic;
signal \N__54837\ : std_logic;
signal \N__54836\ : std_logic;
signal \N__54835\ : std_logic;
signal \N__54834\ : std_logic;
signal \N__54833\ : std_logic;
signal \N__54832\ : std_logic;
signal \N__54829\ : std_logic;
signal \N__54826\ : std_logic;
signal \N__54825\ : std_logic;
signal \N__54822\ : std_logic;
signal \N__54821\ : std_logic;
signal \N__54820\ : std_logic;
signal \N__54819\ : std_logic;
signal \N__54818\ : std_logic;
signal \N__54817\ : std_logic;
signal \N__54816\ : std_logic;
signal \N__54813\ : std_logic;
signal \N__54810\ : std_logic;
signal \N__54807\ : std_logic;
signal \N__54806\ : std_logic;
signal \N__54803\ : std_logic;
signal \N__54802\ : std_logic;
signal \N__54799\ : std_logic;
signal \N__54798\ : std_logic;
signal \N__54795\ : std_logic;
signal \N__54792\ : std_logic;
signal \N__54789\ : std_logic;
signal \N__54784\ : std_logic;
signal \N__54783\ : std_logic;
signal \N__54782\ : std_logic;
signal \N__54781\ : std_logic;
signal \N__54780\ : std_logic;
signal \N__54775\ : std_logic;
signal \N__54772\ : std_logic;
signal \N__54769\ : std_logic;
signal \N__54764\ : std_logic;
signal \N__54761\ : std_logic;
signal \N__54758\ : std_logic;
signal \N__54757\ : std_logic;
signal \N__54756\ : std_logic;
signal \N__54753\ : std_logic;
signal \N__54750\ : std_logic;
signal \N__54747\ : std_logic;
signal \N__54744\ : std_logic;
signal \N__54737\ : std_logic;
signal \N__54736\ : std_logic;
signal \N__54735\ : std_logic;
signal \N__54732\ : std_logic;
signal \N__54729\ : std_logic;
signal \N__54724\ : std_logic;
signal \N__54721\ : std_logic;
signal \N__54712\ : std_logic;
signal \N__54709\ : std_logic;
signal \N__54706\ : std_logic;
signal \N__54703\ : std_logic;
signal \N__54698\ : std_logic;
signal \N__54691\ : std_logic;
signal \N__54686\ : std_logic;
signal \N__54675\ : std_logic;
signal \N__54672\ : std_logic;
signal \N__54669\ : std_logic;
signal \N__54660\ : std_logic;
signal \N__54657\ : std_logic;
signal \N__54654\ : std_logic;
signal \N__54649\ : std_logic;
signal \N__54646\ : std_logic;
signal \N__54639\ : std_logic;
signal \N__54638\ : std_logic;
signal \N__54635\ : std_logic;
signal \N__54634\ : std_logic;
signal \N__54631\ : std_logic;
signal \N__54628\ : std_logic;
signal \N__54623\ : std_logic;
signal \N__54620\ : std_logic;
signal \N__54617\ : std_logic;
signal \N__54614\ : std_logic;
signal \N__54611\ : std_logic;
signal \N__54606\ : std_logic;
signal \N__54603\ : std_logic;
signal \N__54600\ : std_logic;
signal \N__54599\ : std_logic;
signal \N__54598\ : std_logic;
signal \N__54595\ : std_logic;
signal \N__54592\ : std_logic;
signal \N__54589\ : std_logic;
signal \N__54586\ : std_logic;
signal \N__54581\ : std_logic;
signal \N__54576\ : std_logic;
signal \N__54573\ : std_logic;
signal \N__54570\ : std_logic;
signal \N__54567\ : std_logic;
signal \N__54564\ : std_logic;
signal \N__54561\ : std_logic;
signal \N__54558\ : std_logic;
signal \N__54555\ : std_logic;
signal \N__54552\ : std_logic;
signal \N__54549\ : std_logic;
signal \N__54546\ : std_logic;
signal \N__54543\ : std_logic;
signal \N__54540\ : std_logic;
signal \N__54537\ : std_logic;
signal \N__54534\ : std_logic;
signal \N__54531\ : std_logic;
signal \N__54528\ : std_logic;
signal \N__54525\ : std_logic;
signal \N__54524\ : std_logic;
signal \N__54523\ : std_logic;
signal \N__54522\ : std_logic;
signal \N__54521\ : std_logic;
signal \N__54520\ : std_logic;
signal \N__54519\ : std_logic;
signal \N__54518\ : std_logic;
signal \N__54517\ : std_logic;
signal \N__54516\ : std_logic;
signal \N__54515\ : std_logic;
signal \N__54514\ : std_logic;
signal \N__54513\ : std_logic;
signal \N__54512\ : std_logic;
signal \N__54511\ : std_logic;
signal \N__54510\ : std_logic;
signal \N__54509\ : std_logic;
signal \N__54508\ : std_logic;
signal \N__54507\ : std_logic;
signal \N__54506\ : std_logic;
signal \N__54505\ : std_logic;
signal \N__54504\ : std_logic;
signal \N__54503\ : std_logic;
signal \N__54502\ : std_logic;
signal \N__54501\ : std_logic;
signal \N__54500\ : std_logic;
signal \N__54499\ : std_logic;
signal \N__54498\ : std_logic;
signal \N__54497\ : std_logic;
signal \N__54496\ : std_logic;
signal \N__54495\ : std_logic;
signal \N__54494\ : std_logic;
signal \N__54429\ : std_logic;
signal \N__54426\ : std_logic;
signal \N__54423\ : std_logic;
signal \N__54420\ : std_logic;
signal \N__54419\ : std_logic;
signal \N__54416\ : std_logic;
signal \N__54413\ : std_logic;
signal \N__54410\ : std_logic;
signal \N__54405\ : std_logic;
signal \N__54404\ : std_logic;
signal \N__54403\ : std_logic;
signal \N__54402\ : std_logic;
signal \N__54399\ : std_logic;
signal \N__54398\ : std_logic;
signal \N__54395\ : std_logic;
signal \N__54392\ : std_logic;
signal \N__54389\ : std_logic;
signal \N__54384\ : std_logic;
signal \N__54381\ : std_logic;
signal \N__54380\ : std_logic;
signal \N__54373\ : std_logic;
signal \N__54370\ : std_logic;
signal \N__54367\ : std_logic;
signal \N__54364\ : std_logic;
signal \N__54359\ : std_logic;
signal \N__54356\ : std_logic;
signal \N__54351\ : std_logic;
signal \N__54348\ : std_logic;
signal \N__54345\ : std_logic;
signal \N__54344\ : std_logic;
signal \N__54343\ : std_logic;
signal \N__54342\ : std_logic;
signal \N__54339\ : std_logic;
signal \N__54338\ : std_logic;
signal \N__54337\ : std_logic;
signal \N__54336\ : std_logic;
signal \N__54335\ : std_logic;
signal \N__54334\ : std_logic;
signal \N__54331\ : std_logic;
signal \N__54326\ : std_logic;
signal \N__54323\ : std_logic;
signal \N__54320\ : std_logic;
signal \N__54315\ : std_logic;
signal \N__54312\ : std_logic;
signal \N__54309\ : std_logic;
signal \N__54306\ : std_logic;
signal \N__54303\ : std_logic;
signal \N__54300\ : std_logic;
signal \N__54293\ : std_logic;
signal \N__54290\ : std_logic;
signal \N__54289\ : std_logic;
signal \N__54288\ : std_logic;
signal \N__54285\ : std_logic;
signal \N__54282\ : std_logic;
signal \N__54277\ : std_logic;
signal \N__54274\ : std_logic;
signal \N__54269\ : std_logic;
signal \N__54258\ : std_logic;
signal \N__54255\ : std_logic;
signal \N__54252\ : std_logic;
signal \N__54251\ : std_logic;
signal \N__54248\ : std_logic;
signal \N__54245\ : std_logic;
signal \N__54240\ : std_logic;
signal \N__54237\ : std_logic;
signal \N__54234\ : std_logic;
signal \N__54231\ : std_logic;
signal \N__54228\ : std_logic;
signal \N__54225\ : std_logic;
signal \N__54222\ : std_logic;
signal \N__54219\ : std_logic;
signal \N__54216\ : std_logic;
signal \N__54213\ : std_logic;
signal \N__54210\ : std_logic;
signal \N__54207\ : std_logic;
signal \N__54206\ : std_logic;
signal \N__54203\ : std_logic;
signal \N__54200\ : std_logic;
signal \N__54197\ : std_logic;
signal \N__54194\ : std_logic;
signal \N__54193\ : std_logic;
signal \N__54190\ : std_logic;
signal \N__54187\ : std_logic;
signal \N__54184\ : std_logic;
signal \N__54177\ : std_logic;
signal \N__54174\ : std_logic;
signal \N__54171\ : std_logic;
signal \N__54168\ : std_logic;
signal \N__54165\ : std_logic;
signal \N__54162\ : std_logic;
signal \N__54159\ : std_logic;
signal \N__54156\ : std_logic;
signal \N__54153\ : std_logic;
signal \N__54152\ : std_logic;
signal \N__54149\ : std_logic;
signal \N__54146\ : std_logic;
signal \N__54143\ : std_logic;
signal \N__54142\ : std_logic;
signal \N__54139\ : std_logic;
signal \N__54136\ : std_logic;
signal \N__54133\ : std_logic;
signal \N__54130\ : std_logic;
signal \N__54123\ : std_logic;
signal \N__54120\ : std_logic;
signal \N__54119\ : std_logic;
signal \N__54118\ : std_logic;
signal \N__54115\ : std_logic;
signal \N__54114\ : std_logic;
signal \N__54113\ : std_logic;
signal \N__54112\ : std_logic;
signal \N__54109\ : std_logic;
signal \N__54106\ : std_logic;
signal \N__54103\ : std_logic;
signal \N__54100\ : std_logic;
signal \N__54097\ : std_logic;
signal \N__54094\ : std_logic;
signal \N__54091\ : std_logic;
signal \N__54086\ : std_logic;
signal \N__54083\ : std_logic;
signal \N__54080\ : std_logic;
signal \N__54077\ : std_logic;
signal \N__54074\ : std_logic;
signal \N__54071\ : std_logic;
signal \N__54068\ : std_logic;
signal \N__54065\ : std_logic;
signal \N__54060\ : std_logic;
signal \N__54057\ : std_logic;
signal \N__54048\ : std_logic;
signal \N__54045\ : std_logic;
signal \N__54042\ : std_logic;
signal \N__54039\ : std_logic;
signal \N__54036\ : std_logic;
signal \N__54033\ : std_logic;
signal \N__54030\ : std_logic;
signal \N__54027\ : std_logic;
signal \N__54024\ : std_logic;
signal \N__54021\ : std_logic;
signal \N__54018\ : std_logic;
signal \N__54015\ : std_logic;
signal \N__54012\ : std_logic;
signal \N__54009\ : std_logic;
signal \N__54006\ : std_logic;
signal \N__54005\ : std_logic;
signal \N__54004\ : std_logic;
signal \N__54003\ : std_logic;
signal \N__54002\ : std_logic;
signal \N__54001\ : std_logic;
signal \N__53998\ : std_logic;
signal \N__53995\ : std_logic;
signal \N__53994\ : std_logic;
signal \N__53993\ : std_logic;
signal \N__53992\ : std_logic;
signal \N__53991\ : std_logic;
signal \N__53988\ : std_logic;
signal \N__53985\ : std_logic;
signal \N__53980\ : std_logic;
signal \N__53979\ : std_logic;
signal \N__53978\ : std_logic;
signal \N__53977\ : std_logic;
signal \N__53976\ : std_logic;
signal \N__53973\ : std_logic;
signal \N__53970\ : std_logic;
signal \N__53969\ : std_logic;
signal \N__53968\ : std_logic;
signal \N__53967\ : std_logic;
signal \N__53966\ : std_logic;
signal \N__53963\ : std_logic;
signal \N__53962\ : std_logic;
signal \N__53961\ : std_logic;
signal \N__53960\ : std_logic;
signal \N__53959\ : std_logic;
signal \N__53956\ : std_logic;
signal \N__53953\ : std_logic;
signal \N__53950\ : std_logic;
signal \N__53949\ : std_logic;
signal \N__53948\ : std_logic;
signal \N__53945\ : std_logic;
signal \N__53942\ : std_logic;
signal \N__53939\ : std_logic;
signal \N__53934\ : std_logic;
signal \N__53931\ : std_logic;
signal \N__53928\ : std_logic;
signal \N__53925\ : std_logic;
signal \N__53922\ : std_logic;
signal \N__53919\ : std_logic;
signal \N__53914\ : std_logic;
signal \N__53911\ : std_logic;
signal \N__53908\ : std_logic;
signal \N__53905\ : std_logic;
signal \N__53902\ : std_logic;
signal \N__53899\ : std_logic;
signal \N__53896\ : std_logic;
signal \N__53893\ : std_logic;
signal \N__53888\ : std_logic;
signal \N__53885\ : std_logic;
signal \N__53882\ : std_logic;
signal \N__53879\ : std_logic;
signal \N__53874\ : std_logic;
signal \N__53871\ : std_logic;
signal \N__53868\ : std_logic;
signal \N__53865\ : std_logic;
signal \N__53858\ : std_logic;
signal \N__53853\ : std_logic;
signal \N__53832\ : std_logic;
signal \N__53827\ : std_logic;
signal \N__53824\ : std_logic;
signal \N__53819\ : std_logic;
signal \N__53816\ : std_logic;
signal \N__53813\ : std_logic;
signal \N__53810\ : std_logic;
signal \N__53805\ : std_logic;
signal \N__53802\ : std_logic;
signal \N__53793\ : std_logic;
signal \N__53792\ : std_logic;
signal \N__53789\ : std_logic;
signal \N__53788\ : std_logic;
signal \N__53785\ : std_logic;
signal \N__53782\ : std_logic;
signal \N__53779\ : std_logic;
signal \N__53776\ : std_logic;
signal \N__53773\ : std_logic;
signal \N__53770\ : std_logic;
signal \N__53767\ : std_logic;
signal \N__53764\ : std_logic;
signal \N__53761\ : std_logic;
signal \N__53756\ : std_logic;
signal \N__53753\ : std_logic;
signal \N__53750\ : std_logic;
signal \N__53745\ : std_logic;
signal \N__53742\ : std_logic;
signal \N__53739\ : std_logic;
signal \N__53736\ : std_logic;
signal \N__53733\ : std_logic;
signal \N__53730\ : std_logic;
signal \N__53727\ : std_logic;
signal \N__53724\ : std_logic;
signal \N__53721\ : std_logic;
signal \N__53720\ : std_logic;
signal \N__53719\ : std_logic;
signal \N__53718\ : std_logic;
signal \N__53717\ : std_logic;
signal \N__53716\ : std_logic;
signal \N__53715\ : std_logic;
signal \N__53714\ : std_logic;
signal \N__53713\ : std_logic;
signal \N__53712\ : std_logic;
signal \N__53709\ : std_logic;
signal \N__53704\ : std_logic;
signal \N__53701\ : std_logic;
signal \N__53696\ : std_logic;
signal \N__53695\ : std_logic;
signal \N__53694\ : std_logic;
signal \N__53693\ : std_logic;
signal \N__53692\ : std_logic;
signal \N__53691\ : std_logic;
signal \N__53690\ : std_logic;
signal \N__53689\ : std_logic;
signal \N__53684\ : std_logic;
signal \N__53679\ : std_logic;
signal \N__53676\ : std_logic;
signal \N__53675\ : std_logic;
signal \N__53674\ : std_logic;
signal \N__53673\ : std_logic;
signal \N__53672\ : std_logic;
signal \N__53671\ : std_logic;
signal \N__53670\ : std_logic;
signal \N__53669\ : std_logic;
signal \N__53666\ : std_logic;
signal \N__53661\ : std_logic;
signal \N__53656\ : std_logic;
signal \N__53651\ : std_logic;
signal \N__53648\ : std_logic;
signal \N__53643\ : std_logic;
signal \N__53640\ : std_logic;
signal \N__53637\ : std_logic;
signal \N__53634\ : std_logic;
signal \N__53629\ : std_logic;
signal \N__53626\ : std_logic;
signal \N__53623\ : std_logic;
signal \N__53620\ : std_logic;
signal \N__53615\ : std_logic;
signal \N__53610\ : std_logic;
signal \N__53607\ : std_logic;
signal \N__53596\ : std_logic;
signal \N__53593\ : std_logic;
signal \N__53588\ : std_logic;
signal \N__53585\ : std_logic;
signal \N__53578\ : std_logic;
signal \N__53573\ : std_logic;
signal \N__53568\ : std_logic;
signal \N__53565\ : std_logic;
signal \N__53562\ : std_logic;
signal \N__53559\ : std_logic;
signal \N__53556\ : std_logic;
signal \N__53547\ : std_logic;
signal \N__53544\ : std_logic;
signal \N__53541\ : std_logic;
signal \N__53538\ : std_logic;
signal \N__53535\ : std_logic;
signal \N__53532\ : std_logic;
signal \N__53529\ : std_logic;
signal \N__53526\ : std_logic;
signal \N__53525\ : std_logic;
signal \N__53524\ : std_logic;
signal \N__53521\ : std_logic;
signal \N__53518\ : std_logic;
signal \N__53515\ : std_logic;
signal \N__53512\ : std_logic;
signal \N__53509\ : std_logic;
signal \N__53504\ : std_logic;
signal \N__53501\ : std_logic;
signal \N__53496\ : std_logic;
signal \N__53493\ : std_logic;
signal \N__53490\ : std_logic;
signal \N__53487\ : std_logic;
signal \N__53484\ : std_logic;
signal \N__53481\ : std_logic;
signal \N__53478\ : std_logic;
signal \N__53475\ : std_logic;
signal \N__53472\ : std_logic;
signal \N__53469\ : std_logic;
signal \N__53466\ : std_logic;
signal \N__53463\ : std_logic;
signal \N__53460\ : std_logic;
signal \N__53457\ : std_logic;
signal \N__53454\ : std_logic;
signal \N__53451\ : std_logic;
signal \N__53448\ : std_logic;
signal \N__53445\ : std_logic;
signal \N__53442\ : std_logic;
signal \N__53439\ : std_logic;
signal \N__53436\ : std_logic;
signal \N__53433\ : std_logic;
signal \N__53430\ : std_logic;
signal \N__53427\ : std_logic;
signal \N__53424\ : std_logic;
signal \N__53421\ : std_logic;
signal \N__53420\ : std_logic;
signal \N__53419\ : std_logic;
signal \N__53416\ : std_logic;
signal \N__53413\ : std_logic;
signal \N__53410\ : std_logic;
signal \N__53407\ : std_logic;
signal \N__53404\ : std_logic;
signal \N__53401\ : std_logic;
signal \N__53398\ : std_logic;
signal \N__53393\ : std_logic;
signal \N__53390\ : std_logic;
signal \N__53387\ : std_logic;
signal \N__53382\ : std_logic;
signal \N__53379\ : std_logic;
signal \N__53376\ : std_logic;
signal \N__53375\ : std_logic;
signal \N__53372\ : std_logic;
signal \N__53371\ : std_logic;
signal \N__53368\ : std_logic;
signal \N__53365\ : std_logic;
signal \N__53362\ : std_logic;
signal \N__53359\ : std_logic;
signal \N__53356\ : std_logic;
signal \N__53351\ : std_logic;
signal \N__53348\ : std_logic;
signal \N__53345\ : std_logic;
signal \N__53340\ : std_logic;
signal \N__53337\ : std_logic;
signal \N__53334\ : std_logic;
signal \N__53331\ : std_logic;
signal \N__53330\ : std_logic;
signal \N__53329\ : std_logic;
signal \N__53328\ : std_logic;
signal \N__53325\ : std_logic;
signal \N__53324\ : std_logic;
signal \N__53323\ : std_logic;
signal \N__53320\ : std_logic;
signal \N__53319\ : std_logic;
signal \N__53318\ : std_logic;
signal \N__53317\ : std_logic;
signal \N__53316\ : std_logic;
signal \N__53315\ : std_logic;
signal \N__53314\ : std_logic;
signal \N__53311\ : std_logic;
signal \N__53310\ : std_logic;
signal \N__53307\ : std_logic;
signal \N__53306\ : std_logic;
signal \N__53303\ : std_logic;
signal \N__53300\ : std_logic;
signal \N__53297\ : std_logic;
signal \N__53296\ : std_logic;
signal \N__53293\ : std_logic;
signal \N__53290\ : std_logic;
signal \N__53287\ : std_logic;
signal \N__53286\ : std_logic;
signal \N__53283\ : std_logic;
signal \N__53282\ : std_logic;
signal \N__53281\ : std_logic;
signal \N__53278\ : std_logic;
signal \N__53275\ : std_logic;
signal \N__53272\ : std_logic;
signal \N__53271\ : std_logic;
signal \N__53270\ : std_logic;
signal \N__53267\ : std_logic;
signal \N__53266\ : std_logic;
signal \N__53263\ : std_logic;
signal \N__53262\ : std_logic;
signal \N__53259\ : std_logic;
signal \N__53258\ : std_logic;
signal \N__53257\ : std_logic;
signal \N__53256\ : std_logic;
signal \N__53253\ : std_logic;
signal \N__53250\ : std_logic;
signal \N__53247\ : std_logic;
signal \N__53244\ : std_logic;
signal \N__53241\ : std_logic;
signal \N__53238\ : std_logic;
signal \N__53235\ : std_logic;
signal \N__53232\ : std_logic;
signal \N__53229\ : std_logic;
signal \N__53226\ : std_logic;
signal \N__53223\ : std_logic;
signal \N__53220\ : std_logic;
signal \N__53217\ : std_logic;
signal \N__53214\ : std_logic;
signal \N__53211\ : std_logic;
signal \N__53208\ : std_logic;
signal \N__53205\ : std_logic;
signal \N__53202\ : std_logic;
signal \N__53199\ : std_logic;
signal \N__53196\ : std_logic;
signal \N__53195\ : std_logic;
signal \N__53194\ : std_logic;
signal \N__53191\ : std_logic;
signal \N__53188\ : std_logic;
signal \N__53185\ : std_logic;
signal \N__53182\ : std_logic;
signal \N__53181\ : std_logic;
signal \N__53180\ : std_logic;
signal \N__53179\ : std_logic;
signal \N__53176\ : std_logic;
signal \N__53175\ : std_logic;
signal \N__53172\ : std_logic;
signal \N__53167\ : std_logic;
signal \N__53162\ : std_logic;
signal \N__53157\ : std_logic;
signal \N__53154\ : std_logic;
signal \N__53147\ : std_logic;
signal \N__53142\ : std_logic;
signal \N__53137\ : std_logic;
signal \N__53130\ : std_logic;
signal \N__53127\ : std_logic;
signal \N__53124\ : std_logic;
signal \N__53119\ : std_logic;
signal \N__53116\ : std_logic;
signal \N__53111\ : std_logic;
signal \N__53108\ : std_logic;
signal \N__53097\ : std_logic;
signal \N__53090\ : std_logic;
signal \N__53087\ : std_logic;
signal \N__53082\ : std_logic;
signal \N__53075\ : std_logic;
signal \N__53068\ : std_logic;
signal \N__53059\ : std_logic;
signal \N__53056\ : std_logic;
signal \N__53053\ : std_logic;
signal \N__53048\ : std_logic;
signal \N__53043\ : std_logic;
signal \N__53034\ : std_logic;
signal \N__53031\ : std_logic;
signal \N__53028\ : std_logic;
signal \N__53025\ : std_logic;
signal \N__53022\ : std_logic;
signal \N__53019\ : std_logic;
signal \N__53016\ : std_logic;
signal \N__53015\ : std_logic;
signal \N__53014\ : std_logic;
signal \N__53013\ : std_logic;
signal \N__53012\ : std_logic;
signal \N__53011\ : std_logic;
signal \N__53010\ : std_logic;
signal \N__53009\ : std_logic;
signal \N__53008\ : std_logic;
signal \N__53005\ : std_logic;
signal \N__53004\ : std_logic;
signal \N__53001\ : std_logic;
signal \N__53000\ : std_logic;
signal \N__52999\ : std_logic;
signal \N__52998\ : std_logic;
signal \N__52995\ : std_logic;
signal \N__52994\ : std_logic;
signal \N__52991\ : std_logic;
signal \N__52990\ : std_logic;
signal \N__52989\ : std_logic;
signal \N__52988\ : std_logic;
signal \N__52987\ : std_logic;
signal \N__52984\ : std_logic;
signal \N__52983\ : std_logic;
signal \N__52982\ : std_logic;
signal \N__52979\ : std_logic;
signal \N__52976\ : std_logic;
signal \N__52973\ : std_logic;
signal \N__52970\ : std_logic;
signal \N__52967\ : std_logic;
signal \N__52964\ : std_logic;
signal \N__52961\ : std_logic;
signal \N__52958\ : std_logic;
signal \N__52955\ : std_logic;
signal \N__52952\ : std_logic;
signal \N__52949\ : std_logic;
signal \N__52946\ : std_logic;
signal \N__52943\ : std_logic;
signal \N__52940\ : std_logic;
signal \N__52937\ : std_logic;
signal \N__52934\ : std_logic;
signal \N__52931\ : std_logic;
signal \N__52928\ : std_logic;
signal \N__52927\ : std_logic;
signal \N__52926\ : std_logic;
signal \N__52925\ : std_logic;
signal \N__52924\ : std_logic;
signal \N__52923\ : std_logic;
signal \N__52922\ : std_logic;
signal \N__52919\ : std_logic;
signal \N__52916\ : std_logic;
signal \N__52911\ : std_logic;
signal \N__52908\ : std_logic;
signal \N__52905\ : std_logic;
signal \N__52904\ : std_logic;
signal \N__52903\ : std_logic;
signal \N__52902\ : std_logic;
signal \N__52901\ : std_logic;
signal \N__52894\ : std_logic;
signal \N__52885\ : std_logic;
signal \N__52882\ : std_logic;
signal \N__52877\ : std_logic;
signal \N__52872\ : std_logic;
signal \N__52867\ : std_logic;
signal \N__52854\ : std_logic;
signal \N__52847\ : std_logic;
signal \N__52842\ : std_logic;
signal \N__52833\ : std_logic;
signal \N__52830\ : std_logic;
signal \N__52827\ : std_logic;
signal \N__52816\ : std_logic;
signal \N__52803\ : std_logic;
signal \N__52800\ : std_logic;
signal \N__52797\ : std_logic;
signal \N__52794\ : std_logic;
signal \N__52791\ : std_logic;
signal \N__52788\ : std_logic;
signal \N__52785\ : std_logic;
signal \N__52782\ : std_logic;
signal \N__52781\ : std_logic;
signal \N__52780\ : std_logic;
signal \N__52779\ : std_logic;
signal \N__52776\ : std_logic;
signal \N__52773\ : std_logic;
signal \N__52772\ : std_logic;
signal \N__52771\ : std_logic;
signal \N__52770\ : std_logic;
signal \N__52769\ : std_logic;
signal \N__52768\ : std_logic;
signal \N__52765\ : std_logic;
signal \N__52762\ : std_logic;
signal \N__52761\ : std_logic;
signal \N__52760\ : std_logic;
signal \N__52757\ : std_logic;
signal \N__52756\ : std_logic;
signal \N__52755\ : std_logic;
signal \N__52752\ : std_logic;
signal \N__52749\ : std_logic;
signal \N__52746\ : std_logic;
signal \N__52745\ : std_logic;
signal \N__52744\ : std_logic;
signal \N__52743\ : std_logic;
signal \N__52742\ : std_logic;
signal \N__52741\ : std_logic;
signal \N__52740\ : std_logic;
signal \N__52739\ : std_logic;
signal \N__52738\ : std_logic;
signal \N__52737\ : std_logic;
signal \N__52736\ : std_logic;
signal \N__52733\ : std_logic;
signal \N__52730\ : std_logic;
signal \N__52727\ : std_logic;
signal \N__52722\ : std_logic;
signal \N__52719\ : std_logic;
signal \N__52716\ : std_logic;
signal \N__52713\ : std_logic;
signal \N__52710\ : std_logic;
signal \N__52707\ : std_logic;
signal \N__52702\ : std_logic;
signal \N__52701\ : std_logic;
signal \N__52700\ : std_logic;
signal \N__52697\ : std_logic;
signal \N__52694\ : std_logic;
signal \N__52691\ : std_logic;
signal \N__52688\ : std_logic;
signal \N__52685\ : std_logic;
signal \N__52682\ : std_logic;
signal \N__52677\ : std_logic;
signal \N__52676\ : std_logic;
signal \N__52675\ : std_logic;
signal \N__52674\ : std_logic;
signal \N__52673\ : std_logic;
signal \N__52672\ : std_logic;
signal \N__52669\ : std_logic;
signal \N__52666\ : std_logic;
signal \N__52663\ : std_logic;
signal \N__52660\ : std_logic;
signal \N__52657\ : std_logic;
signal \N__52648\ : std_logic;
signal \N__52643\ : std_logic;
signal \N__52640\ : std_logic;
signal \N__52637\ : std_logic;
signal \N__52634\ : std_logic;
signal \N__52631\ : std_logic;
signal \N__52626\ : std_logic;
signal \N__52621\ : std_logic;
signal \N__52614\ : std_logic;
signal \N__52611\ : std_logic;
signal \N__52608\ : std_logic;
signal \N__52605\ : std_logic;
signal \N__52602\ : std_logic;
signal \N__52599\ : std_logic;
signal \N__52592\ : std_logic;
signal \N__52585\ : std_logic;
signal \N__52578\ : std_logic;
signal \N__52567\ : std_logic;
signal \N__52548\ : std_logic;
signal \N__52545\ : std_logic;
signal \N__52542\ : std_logic;
signal \N__52539\ : std_logic;
signal \N__52536\ : std_logic;
signal \N__52533\ : std_logic;
signal \N__52530\ : std_logic;
signal \N__52527\ : std_logic;
signal \N__52526\ : std_logic;
signal \N__52525\ : std_logic;
signal \N__52524\ : std_logic;
signal \N__52523\ : std_logic;
signal \N__52522\ : std_logic;
signal \N__52521\ : std_logic;
signal \N__52520\ : std_logic;
signal \N__52517\ : std_logic;
signal \N__52514\ : std_logic;
signal \N__52513\ : std_logic;
signal \N__52512\ : std_logic;
signal \N__52509\ : std_logic;
signal \N__52506\ : std_logic;
signal \N__52503\ : std_logic;
signal \N__52500\ : std_logic;
signal \N__52497\ : std_logic;
signal \N__52496\ : std_logic;
signal \N__52495\ : std_logic;
signal \N__52494\ : std_logic;
signal \N__52493\ : std_logic;
signal \N__52492\ : std_logic;
signal \N__52489\ : std_logic;
signal \N__52488\ : std_logic;
signal \N__52487\ : std_logic;
signal \N__52486\ : std_logic;
signal \N__52485\ : std_logic;
signal \N__52484\ : std_logic;
signal \N__52481\ : std_logic;
signal \N__52478\ : std_logic;
signal \N__52475\ : std_logic;
signal \N__52472\ : std_logic;
signal \N__52471\ : std_logic;
signal \N__52468\ : std_logic;
signal \N__52463\ : std_logic;
signal \N__52458\ : std_logic;
signal \N__52455\ : std_logic;
signal \N__52450\ : std_logic;
signal \N__52447\ : std_logic;
signal \N__52446\ : std_logic;
signal \N__52445\ : std_logic;
signal \N__52442\ : std_logic;
signal \N__52441\ : std_logic;
signal \N__52440\ : std_logic;
signal \N__52439\ : std_logic;
signal \N__52438\ : std_logic;
signal \N__52437\ : std_logic;
signal \N__52434\ : std_logic;
signal \N__52431\ : std_logic;
signal \N__52428\ : std_logic;
signal \N__52425\ : std_logic;
signal \N__52422\ : std_logic;
signal \N__52419\ : std_logic;
signal \N__52410\ : std_logic;
signal \N__52407\ : std_logic;
signal \N__52404\ : std_logic;
signal \N__52399\ : std_logic;
signal \N__52396\ : std_logic;
signal \N__52391\ : std_logic;
signal \N__52388\ : std_logic;
signal \N__52385\ : std_logic;
signal \N__52382\ : std_logic;
signal \N__52381\ : std_logic;
signal \N__52378\ : std_logic;
signal \N__52375\ : std_logic;
signal \N__52372\ : std_logic;
signal \N__52371\ : std_logic;
signal \N__52370\ : std_logic;
signal \N__52367\ : std_logic;
signal \N__52364\ : std_logic;
signal \N__52357\ : std_logic;
signal \N__52354\ : std_logic;
signal \N__52349\ : std_logic;
signal \N__52344\ : std_logic;
signal \N__52333\ : std_logic;
signal \N__52330\ : std_logic;
signal \N__52327\ : std_logic;
signal \N__52324\ : std_logic;
signal \N__52319\ : std_logic;
signal \N__52316\ : std_logic;
signal \N__52311\ : std_logic;
signal \N__52308\ : std_logic;
signal \N__52303\ : std_logic;
signal \N__52298\ : std_logic;
signal \N__52293\ : std_logic;
signal \N__52284\ : std_logic;
signal \N__52279\ : std_logic;
signal \N__52276\ : std_logic;
signal \N__52271\ : std_logic;
signal \N__52268\ : std_logic;
signal \N__52263\ : std_logic;
signal \N__52254\ : std_logic;
signal \N__52251\ : std_logic;
signal \N__52248\ : std_logic;
signal \N__52245\ : std_logic;
signal \N__52242\ : std_logic;
signal \N__52239\ : std_logic;
signal \N__52236\ : std_logic;
signal \N__52235\ : std_logic;
signal \N__52234\ : std_logic;
signal \N__52233\ : std_logic;
signal \N__52232\ : std_logic;
signal \N__52231\ : std_logic;
signal \N__52228\ : std_logic;
signal \N__52227\ : std_logic;
signal \N__52224\ : std_logic;
signal \N__52223\ : std_logic;
signal \N__52222\ : std_logic;
signal \N__52221\ : std_logic;
signal \N__52220\ : std_logic;
signal \N__52217\ : std_logic;
signal \N__52216\ : std_logic;
signal \N__52215\ : std_logic;
signal \N__52214\ : std_logic;
signal \N__52213\ : std_logic;
signal \N__52210\ : std_logic;
signal \N__52207\ : std_logic;
signal \N__52206\ : std_logic;
signal \N__52205\ : std_logic;
signal \N__52204\ : std_logic;
signal \N__52203\ : std_logic;
signal \N__52200\ : std_logic;
signal \N__52199\ : std_logic;
signal \N__52198\ : std_logic;
signal \N__52195\ : std_logic;
signal \N__52192\ : std_logic;
signal \N__52191\ : std_logic;
signal \N__52188\ : std_logic;
signal \N__52187\ : std_logic;
signal \N__52186\ : std_logic;
signal \N__52183\ : std_logic;
signal \N__52182\ : std_logic;
signal \N__52179\ : std_logic;
signal \N__52176\ : std_logic;
signal \N__52173\ : std_logic;
signal \N__52170\ : std_logic;
signal \N__52167\ : std_logic;
signal \N__52164\ : std_logic;
signal \N__52161\ : std_logic;
signal \N__52158\ : std_logic;
signal \N__52153\ : std_logic;
signal \N__52150\ : std_logic;
signal \N__52147\ : std_logic;
signal \N__52146\ : std_logic;
signal \N__52145\ : std_logic;
signal \N__52142\ : std_logic;
signal \N__52139\ : std_logic;
signal \N__52136\ : std_logic;
signal \N__52133\ : std_logic;
signal \N__52130\ : std_logic;
signal \N__52125\ : std_logic;
signal \N__52124\ : std_logic;
signal \N__52123\ : std_logic;
signal \N__52122\ : std_logic;
signal \N__52119\ : std_logic;
signal \N__52116\ : std_logic;
signal \N__52113\ : std_logic;
signal \N__52110\ : std_logic;
signal \N__52107\ : std_logic;
signal \N__52104\ : std_logic;
signal \N__52099\ : std_logic;
signal \N__52090\ : std_logic;
signal \N__52087\ : std_logic;
signal \N__52080\ : std_logic;
signal \N__52077\ : std_logic;
signal \N__52074\ : std_logic;
signal \N__52071\ : std_logic;
signal \N__52066\ : std_logic;
signal \N__52061\ : std_logic;
signal \N__52058\ : std_logic;
signal \N__52055\ : std_logic;
signal \N__52054\ : std_logic;
signal \N__52051\ : std_logic;
signal \N__52048\ : std_logic;
signal \N__52045\ : std_logic;
signal \N__52038\ : std_logic;
signal \N__52027\ : std_logic;
signal \N__52020\ : std_logic;
signal \N__52017\ : std_logic;
signal \N__52006\ : std_logic;
signal \N__52003\ : std_logic;
signal \N__51984\ : std_logic;
signal \N__51981\ : std_logic;
signal \N__51978\ : std_logic;
signal \N__51975\ : std_logic;
signal \N__51972\ : std_logic;
signal \N__51969\ : std_logic;
signal \N__51966\ : std_logic;
signal \N__51963\ : std_logic;
signal \N__51960\ : std_logic;
signal \N__51957\ : std_logic;
signal \N__51954\ : std_logic;
signal \N__51951\ : std_logic;
signal \N__51950\ : std_logic;
signal \N__51947\ : std_logic;
signal \N__51946\ : std_logic;
signal \N__51943\ : std_logic;
signal \N__51940\ : std_logic;
signal \N__51937\ : std_logic;
signal \N__51936\ : std_logic;
signal \N__51931\ : std_logic;
signal \N__51928\ : std_logic;
signal \N__51927\ : std_logic;
signal \N__51926\ : std_logic;
signal \N__51925\ : std_logic;
signal \N__51924\ : std_logic;
signal \N__51923\ : std_logic;
signal \N__51922\ : std_logic;
signal \N__51921\ : std_logic;
signal \N__51920\ : std_logic;
signal \N__51919\ : std_logic;
signal \N__51916\ : std_logic;
signal \N__51915\ : std_logic;
signal \N__51910\ : std_logic;
signal \N__51907\ : std_logic;
signal \N__51906\ : std_logic;
signal \N__51905\ : std_logic;
signal \N__51904\ : std_logic;
signal \N__51903\ : std_logic;
signal \N__51902\ : std_logic;
signal \N__51899\ : std_logic;
signal \N__51896\ : std_logic;
signal \N__51893\ : std_logic;
signal \N__51892\ : std_logic;
signal \N__51891\ : std_logic;
signal \N__51890\ : std_logic;
signal \N__51887\ : std_logic;
signal \N__51884\ : std_logic;
signal \N__51881\ : std_logic;
signal \N__51878\ : std_logic;
signal \N__51875\ : std_logic;
signal \N__51872\ : std_logic;
signal \N__51871\ : std_logic;
signal \N__51868\ : std_logic;
signal \N__51867\ : std_logic;
signal \N__51866\ : std_logic;
signal \N__51861\ : std_logic;
signal \N__51860\ : std_logic;
signal \N__51859\ : std_logic;
signal \N__51856\ : std_logic;
signal \N__51853\ : std_logic;
signal \N__51850\ : std_logic;
signal \N__51847\ : std_logic;
signal \N__51846\ : std_logic;
signal \N__51843\ : std_logic;
signal \N__51840\ : std_logic;
signal \N__51837\ : std_logic;
signal \N__51834\ : std_logic;
signal \N__51831\ : std_logic;
signal \N__51828\ : std_logic;
signal \N__51825\ : std_logic;
signal \N__51824\ : std_logic;
signal \N__51821\ : std_logic;
signal \N__51814\ : std_logic;
signal \N__51809\ : std_logic;
signal \N__51804\ : std_logic;
signal \N__51801\ : std_logic;
signal \N__51798\ : std_logic;
signal \N__51795\ : std_logic;
signal \N__51792\ : std_logic;
signal \N__51791\ : std_logic;
signal \N__51790\ : std_logic;
signal \N__51787\ : std_logic;
signal \N__51784\ : std_logic;
signal \N__51781\ : std_logic;
signal \N__51776\ : std_logic;
signal \N__51773\ : std_logic;
signal \N__51770\ : std_logic;
signal \N__51765\ : std_logic;
signal \N__51760\ : std_logic;
signal \N__51755\ : std_logic;
signal \N__51752\ : std_logic;
signal \N__51743\ : std_logic;
signal \N__51740\ : std_logic;
signal \N__51733\ : std_logic;
signal \N__51730\ : std_logic;
signal \N__51727\ : std_logic;
signal \N__51718\ : std_logic;
signal \N__51707\ : std_logic;
signal \N__51702\ : std_logic;
signal \N__51697\ : std_logic;
signal \N__51684\ : std_logic;
signal \N__51681\ : std_logic;
signal \N__51678\ : std_logic;
signal \N__51675\ : std_logic;
signal \N__51672\ : std_logic;
signal \N__51669\ : std_logic;
signal \N__51666\ : std_logic;
signal \N__51663\ : std_logic;
signal \N__51660\ : std_logic;
signal \N__51657\ : std_logic;
signal \N__51656\ : std_logic;
signal \N__51653\ : std_logic;
signal \N__51652\ : std_logic;
signal \N__51649\ : std_logic;
signal \N__51646\ : std_logic;
signal \N__51643\ : std_logic;
signal \N__51640\ : std_logic;
signal \N__51637\ : std_logic;
signal \N__51634\ : std_logic;
signal \N__51631\ : std_logic;
signal \N__51624\ : std_logic;
signal \N__51621\ : std_logic;
signal \N__51620\ : std_logic;
signal \N__51617\ : std_logic;
signal \N__51614\ : std_logic;
signal \N__51611\ : std_logic;
signal \N__51610\ : std_logic;
signal \N__51607\ : std_logic;
signal \N__51604\ : std_logic;
signal \N__51601\ : std_logic;
signal \N__51598\ : std_logic;
signal \N__51591\ : std_logic;
signal \N__51588\ : std_logic;
signal \N__51587\ : std_logic;
signal \N__51586\ : std_logic;
signal \N__51583\ : std_logic;
signal \N__51580\ : std_logic;
signal \N__51577\ : std_logic;
signal \N__51574\ : std_logic;
signal \N__51571\ : std_logic;
signal \N__51568\ : std_logic;
signal \N__51565\ : std_logic;
signal \N__51562\ : std_logic;
signal \N__51555\ : std_logic;
signal \N__51552\ : std_logic;
signal \N__51549\ : std_logic;
signal \N__51546\ : std_logic;
signal \N__51543\ : std_logic;
signal \N__51540\ : std_logic;
signal \N__51537\ : std_logic;
signal \N__51534\ : std_logic;
signal \N__51531\ : std_logic;
signal \N__51528\ : std_logic;
signal \N__51525\ : std_logic;
signal \N__51522\ : std_logic;
signal \N__51519\ : std_logic;
signal \N__51516\ : std_logic;
signal \N__51513\ : std_logic;
signal \N__51510\ : std_logic;
signal \N__51507\ : std_logic;
signal \N__51506\ : std_logic;
signal \N__51505\ : std_logic;
signal \N__51502\ : std_logic;
signal \N__51499\ : std_logic;
signal \N__51496\ : std_logic;
signal \N__51493\ : std_logic;
signal \N__51490\ : std_logic;
signal \N__51487\ : std_logic;
signal \N__51482\ : std_logic;
signal \N__51477\ : std_logic;
signal \N__51476\ : std_logic;
signal \N__51473\ : std_logic;
signal \N__51470\ : std_logic;
signal \N__51467\ : std_logic;
signal \N__51464\ : std_logic;
signal \N__51463\ : std_logic;
signal \N__51460\ : std_logic;
signal \N__51457\ : std_logic;
signal \N__51454\ : std_logic;
signal \N__51447\ : std_logic;
signal \N__51444\ : std_logic;
signal \N__51441\ : std_logic;
signal \N__51438\ : std_logic;
signal \N__51435\ : std_logic;
signal \N__51434\ : std_logic;
signal \N__51431\ : std_logic;
signal \N__51430\ : std_logic;
signal \N__51427\ : std_logic;
signal \N__51424\ : std_logic;
signal \N__51421\ : std_logic;
signal \N__51418\ : std_logic;
signal \N__51415\ : std_logic;
signal \N__51412\ : std_logic;
signal \N__51409\ : std_logic;
signal \N__51402\ : std_logic;
signal \N__51399\ : std_logic;
signal \N__51396\ : std_logic;
signal \N__51395\ : std_logic;
signal \N__51392\ : std_logic;
signal \N__51389\ : std_logic;
signal \N__51386\ : std_logic;
signal \N__51383\ : std_logic;
signal \N__51382\ : std_logic;
signal \N__51377\ : std_logic;
signal \N__51374\ : std_logic;
signal \N__51369\ : std_logic;
signal \N__51368\ : std_logic;
signal \N__51365\ : std_logic;
signal \N__51364\ : std_logic;
signal \N__51361\ : std_logic;
signal \N__51358\ : std_logic;
signal \N__51355\ : std_logic;
signal \N__51352\ : std_logic;
signal \N__51347\ : std_logic;
signal \N__51342\ : std_logic;
signal \N__51339\ : std_logic;
signal \N__51336\ : std_logic;
signal \N__51333\ : std_logic;
signal \N__51330\ : std_logic;
signal \N__51327\ : std_logic;
signal \N__51324\ : std_logic;
signal \N__51321\ : std_logic;
signal \N__51318\ : std_logic;
signal \N__51315\ : std_logic;
signal \N__51312\ : std_logic;
signal \N__51309\ : std_logic;
signal \N__51306\ : std_logic;
signal \N__51303\ : std_logic;
signal \N__51300\ : std_logic;
signal \N__51299\ : std_logic;
signal \N__51296\ : std_logic;
signal \N__51293\ : std_logic;
signal \N__51290\ : std_logic;
signal \N__51285\ : std_logic;
signal \N__51282\ : std_logic;
signal \N__51279\ : std_logic;
signal \N__51276\ : std_logic;
signal \N__51273\ : std_logic;
signal \N__51270\ : std_logic;
signal \N__51267\ : std_logic;
signal \N__51264\ : std_logic;
signal \N__51261\ : std_logic;
signal \N__51258\ : std_logic;
signal \N__51255\ : std_logic;
signal \N__51252\ : std_logic;
signal \N__51251\ : std_logic;
signal \N__51248\ : std_logic;
signal \N__51245\ : std_logic;
signal \N__51242\ : std_logic;
signal \N__51241\ : std_logic;
signal \N__51238\ : std_logic;
signal \N__51235\ : std_logic;
signal \N__51232\ : std_logic;
signal \N__51229\ : std_logic;
signal \N__51224\ : std_logic;
signal \N__51221\ : std_logic;
signal \N__51218\ : std_logic;
signal \N__51213\ : std_logic;
signal \N__51210\ : std_logic;
signal \N__51207\ : std_logic;
signal \N__51206\ : std_logic;
signal \N__51203\ : std_logic;
signal \N__51200\ : std_logic;
signal \N__51197\ : std_logic;
signal \N__51194\ : std_logic;
signal \N__51191\ : std_logic;
signal \N__51190\ : std_logic;
signal \N__51187\ : std_logic;
signal \N__51186\ : std_logic;
signal \N__51183\ : std_logic;
signal \N__51180\ : std_logic;
signal \N__51177\ : std_logic;
signal \N__51174\ : std_logic;
signal \N__51171\ : std_logic;
signal \N__51168\ : std_logic;
signal \N__51163\ : std_logic;
signal \N__51160\ : std_logic;
signal \N__51157\ : std_logic;
signal \N__51154\ : std_logic;
signal \N__51151\ : std_logic;
signal \N__51148\ : std_logic;
signal \N__51145\ : std_logic;
signal \N__51142\ : std_logic;
signal \N__51139\ : std_logic;
signal \N__51136\ : std_logic;
signal \N__51129\ : std_logic;
signal \N__51126\ : std_logic;
signal \N__51123\ : std_logic;
signal \N__51122\ : std_logic;
signal \N__51121\ : std_logic;
signal \N__51120\ : std_logic;
signal \N__51119\ : std_logic;
signal \N__51118\ : std_logic;
signal \N__51113\ : std_logic;
signal \N__51104\ : std_logic;
signal \N__51101\ : std_logic;
signal \N__51098\ : std_logic;
signal \N__51095\ : std_logic;
signal \N__51092\ : std_logic;
signal \N__51089\ : std_logic;
signal \N__51086\ : std_logic;
signal \N__51081\ : std_logic;
signal \N__51080\ : std_logic;
signal \N__51079\ : std_logic;
signal \N__51078\ : std_logic;
signal \N__51077\ : std_logic;
signal \N__51076\ : std_logic;
signal \N__51075\ : std_logic;
signal \N__51070\ : std_logic;
signal \N__51059\ : std_logic;
signal \N__51054\ : std_logic;
signal \N__51053\ : std_logic;
signal \N__51052\ : std_logic;
signal \N__51049\ : std_logic;
signal \N__51048\ : std_logic;
signal \N__51045\ : std_logic;
signal \N__51044\ : std_logic;
signal \N__51037\ : std_logic;
signal \N__51032\ : std_logic;
signal \N__51029\ : std_logic;
signal \N__51024\ : std_logic;
signal \N__51023\ : std_logic;
signal \N__51022\ : std_logic;
signal \N__51019\ : std_logic;
signal \N__51016\ : std_logic;
signal \N__51015\ : std_logic;
signal \N__51014\ : std_logic;
signal \N__51013\ : std_logic;
signal \N__51008\ : std_logic;
signal \N__50999\ : std_logic;
signal \N__50994\ : std_logic;
signal \N__50993\ : std_logic;
signal \N__50990\ : std_logic;
signal \N__50987\ : std_logic;
signal \N__50984\ : std_logic;
signal \N__50983\ : std_logic;
signal \N__50980\ : std_logic;
signal \N__50979\ : std_logic;
signal \N__50976\ : std_logic;
signal \N__50973\ : std_logic;
signal \N__50970\ : std_logic;
signal \N__50967\ : std_logic;
signal \N__50960\ : std_logic;
signal \N__50955\ : std_logic;
signal \N__50952\ : std_logic;
signal \N__50949\ : std_logic;
signal \N__50946\ : std_logic;
signal \N__50943\ : std_logic;
signal \N__50940\ : std_logic;
signal \N__50937\ : std_logic;
signal \N__50934\ : std_logic;
signal \N__50933\ : std_logic;
signal \N__50932\ : std_logic;
signal \N__50931\ : std_logic;
signal \N__50930\ : std_logic;
signal \N__50927\ : std_logic;
signal \N__50924\ : std_logic;
signal \N__50923\ : std_logic;
signal \N__50922\ : std_logic;
signal \N__50921\ : std_logic;
signal \N__50914\ : std_logic;
signal \N__50909\ : std_logic;
signal \N__50902\ : std_logic;
signal \N__50899\ : std_logic;
signal \N__50896\ : std_logic;
signal \N__50893\ : std_logic;
signal \N__50886\ : std_logic;
signal \N__50885\ : std_logic;
signal \N__50884\ : std_logic;
signal \N__50883\ : std_logic;
signal \N__50882\ : std_logic;
signal \N__50881\ : std_logic;
signal \N__50878\ : std_logic;
signal \N__50875\ : std_logic;
signal \N__50874\ : std_logic;
signal \N__50873\ : std_logic;
signal \N__50872\ : std_logic;
signal \N__50871\ : std_logic;
signal \N__50866\ : std_logic;
signal \N__50865\ : std_logic;
signal \N__50864\ : std_logic;
signal \N__50861\ : std_logic;
signal \N__50858\ : std_logic;
signal \N__50855\ : std_logic;
signal \N__50844\ : std_logic;
signal \N__50841\ : std_logic;
signal \N__50836\ : std_logic;
signal \N__50833\ : std_logic;
signal \N__50830\ : std_logic;
signal \N__50821\ : std_logic;
signal \N__50820\ : std_logic;
signal \N__50817\ : std_logic;
signal \N__50814\ : std_logic;
signal \N__50811\ : std_logic;
signal \N__50808\ : std_logic;
signal \N__50805\ : std_logic;
signal \N__50802\ : std_logic;
signal \N__50797\ : std_logic;
signal \N__50790\ : std_logic;
signal \N__50787\ : std_logic;
signal \N__50784\ : std_logic;
signal \N__50781\ : std_logic;
signal \N__50778\ : std_logic;
signal \N__50775\ : std_logic;
signal \N__50772\ : std_logic;
signal \N__50769\ : std_logic;
signal \N__50766\ : std_logic;
signal \N__50763\ : std_logic;
signal \N__50760\ : std_logic;
signal \N__50757\ : std_logic;
signal \N__50754\ : std_logic;
signal \N__50751\ : std_logic;
signal \N__50748\ : std_logic;
signal \N__50747\ : std_logic;
signal \N__50746\ : std_logic;
signal \N__50743\ : std_logic;
signal \N__50738\ : std_logic;
signal \N__50735\ : std_logic;
signal \N__50732\ : std_logic;
signal \N__50727\ : std_logic;
signal \N__50724\ : std_logic;
signal \N__50721\ : std_logic;
signal \N__50718\ : std_logic;
signal \N__50717\ : std_logic;
signal \N__50716\ : std_logic;
signal \N__50715\ : std_logic;
signal \N__50714\ : std_logic;
signal \N__50711\ : std_logic;
signal \N__50706\ : std_logic;
signal \N__50701\ : std_logic;
signal \N__50698\ : std_logic;
signal \N__50693\ : std_logic;
signal \N__50690\ : std_logic;
signal \N__50687\ : std_logic;
signal \N__50682\ : std_logic;
signal \N__50681\ : std_logic;
signal \N__50678\ : std_logic;
signal \N__50675\ : std_logic;
signal \N__50670\ : std_logic;
signal \N__50667\ : std_logic;
signal \N__50666\ : std_logic;
signal \N__50663\ : std_logic;
signal \N__50660\ : std_logic;
signal \N__50655\ : std_logic;
signal \N__50652\ : std_logic;
signal \N__50649\ : std_logic;
signal \N__50646\ : std_logic;
signal \N__50643\ : std_logic;
signal \N__50642\ : std_logic;
signal \N__50637\ : std_logic;
signal \N__50634\ : std_logic;
signal \N__50631\ : std_logic;
signal \N__50628\ : std_logic;
signal \N__50625\ : std_logic;
signal \N__50622\ : std_logic;
signal \N__50621\ : std_logic;
signal \N__50618\ : std_logic;
signal \N__50615\ : std_logic;
signal \N__50612\ : std_logic;
signal \N__50611\ : std_logic;
signal \N__50608\ : std_logic;
signal \N__50605\ : std_logic;
signal \N__50602\ : std_logic;
signal \N__50597\ : std_logic;
signal \N__50592\ : std_logic;
signal \N__50589\ : std_logic;
signal \N__50586\ : std_logic;
signal \N__50585\ : std_logic;
signal \N__50582\ : std_logic;
signal \N__50581\ : std_logic;
signal \N__50578\ : std_logic;
signal \N__50575\ : std_logic;
signal \N__50572\ : std_logic;
signal \N__50565\ : std_logic;
signal \N__50562\ : std_logic;
signal \N__50559\ : std_logic;
signal \N__50558\ : std_logic;
signal \N__50555\ : std_logic;
signal \N__50552\ : std_logic;
signal \N__50551\ : std_logic;
signal \N__50546\ : std_logic;
signal \N__50545\ : std_logic;
signal \N__50544\ : std_logic;
signal \N__50543\ : std_logic;
signal \N__50540\ : std_logic;
signal \N__50539\ : std_logic;
signal \N__50538\ : std_logic;
signal \N__50537\ : std_logic;
signal \N__50536\ : std_logic;
signal \N__50533\ : std_logic;
signal \N__50530\ : std_logic;
signal \N__50525\ : std_logic;
signal \N__50522\ : std_logic;
signal \N__50517\ : std_logic;
signal \N__50512\ : std_logic;
signal \N__50509\ : std_logic;
signal \N__50506\ : std_logic;
signal \N__50493\ : std_logic;
signal \N__50490\ : std_logic;
signal \N__50487\ : std_logic;
signal \N__50484\ : std_logic;
signal \N__50481\ : std_logic;
signal \N__50478\ : std_logic;
signal \N__50475\ : std_logic;
signal \N__50472\ : std_logic;
signal \N__50469\ : std_logic;
signal \N__50466\ : std_logic;
signal \N__50463\ : std_logic;
signal \N__50460\ : std_logic;
signal \N__50457\ : std_logic;
signal \N__50456\ : std_logic;
signal \N__50453\ : std_logic;
signal \N__50450\ : std_logic;
signal \N__50449\ : std_logic;
signal \N__50446\ : std_logic;
signal \N__50443\ : std_logic;
signal \N__50440\ : std_logic;
signal \N__50437\ : std_logic;
signal \N__50434\ : std_logic;
signal \N__50427\ : std_logic;
signal \N__50424\ : std_logic;
signal \N__50421\ : std_logic;
signal \N__50418\ : std_logic;
signal \N__50415\ : std_logic;
signal \N__50412\ : std_logic;
signal \N__50409\ : std_logic;
signal \N__50408\ : std_logic;
signal \N__50407\ : std_logic;
signal \N__50406\ : std_logic;
signal \N__50405\ : std_logic;
signal \N__50404\ : std_logic;
signal \N__50403\ : std_logic;
signal \N__50402\ : std_logic;
signal \N__50401\ : std_logic;
signal \N__50398\ : std_logic;
signal \N__50397\ : std_logic;
signal \N__50396\ : std_logic;
signal \N__50395\ : std_logic;
signal \N__50394\ : std_logic;
signal \N__50393\ : std_logic;
signal \N__50392\ : std_logic;
signal \N__50391\ : std_logic;
signal \N__50390\ : std_logic;
signal \N__50389\ : std_logic;
signal \N__50388\ : std_logic;
signal \N__50387\ : std_logic;
signal \N__50386\ : std_logic;
signal \N__50381\ : std_logic;
signal \N__50380\ : std_logic;
signal \N__50379\ : std_logic;
signal \N__50368\ : std_logic;
signal \N__50359\ : std_logic;
signal \N__50356\ : std_logic;
signal \N__50355\ : std_logic;
signal \N__50354\ : std_logic;
signal \N__50353\ : std_logic;
signal \N__50352\ : std_logic;
signal \N__50351\ : std_logic;
signal \N__50350\ : std_logic;
signal \N__50349\ : std_logic;
signal \N__50348\ : std_logic;
signal \N__50347\ : std_logic;
signal \N__50334\ : std_logic;
signal \N__50329\ : std_logic;
signal \N__50326\ : std_logic;
signal \N__50323\ : std_logic;
signal \N__50318\ : std_logic;
signal \N__50313\ : std_logic;
signal \N__50308\ : std_logic;
signal \N__50301\ : std_logic;
signal \N__50290\ : std_logic;
signal \N__50285\ : std_logic;
signal \N__50282\ : std_logic;
signal \N__50277\ : std_logic;
signal \N__50274\ : std_logic;
signal \N__50265\ : std_logic;
signal \N__50262\ : std_logic;
signal \N__50257\ : std_logic;
signal \N__50254\ : std_logic;
signal \N__50251\ : std_logic;
signal \N__50248\ : std_logic;
signal \N__50245\ : std_logic;
signal \N__50244\ : std_logic;
signal \N__50239\ : std_logic;
signal \N__50236\ : std_logic;
signal \N__50233\ : std_logic;
signal \N__50226\ : std_logic;
signal \N__50223\ : std_logic;
signal \N__50220\ : std_logic;
signal \N__50219\ : std_logic;
signal \N__50218\ : std_logic;
signal \N__50215\ : std_logic;
signal \N__50208\ : std_logic;
signal \N__50205\ : std_logic;
signal \N__50202\ : std_logic;
signal \N__50199\ : std_logic;
signal \N__50196\ : std_logic;
signal \N__50193\ : std_logic;
signal \N__50192\ : std_logic;
signal \N__50191\ : std_logic;
signal \N__50188\ : std_logic;
signal \N__50185\ : std_logic;
signal \N__50182\ : std_logic;
signal \N__50175\ : std_logic;
signal \N__50172\ : std_logic;
signal \N__50169\ : std_logic;
signal \N__50166\ : std_logic;
signal \N__50163\ : std_logic;
signal \N__50160\ : std_logic;
signal \N__50157\ : std_logic;
signal \N__50154\ : std_logic;
signal \N__50151\ : std_logic;
signal \N__50148\ : std_logic;
signal \N__50145\ : std_logic;
signal \N__50142\ : std_logic;
signal \N__50141\ : std_logic;
signal \N__50140\ : std_logic;
signal \N__50139\ : std_logic;
signal \N__50138\ : std_logic;
signal \N__50137\ : std_logic;
signal \N__50134\ : std_logic;
signal \N__50131\ : std_logic;
signal \N__50126\ : std_logic;
signal \N__50121\ : std_logic;
signal \N__50114\ : std_logic;
signal \N__50113\ : std_logic;
signal \N__50112\ : std_logic;
signal \N__50109\ : std_logic;
signal \N__50106\ : std_logic;
signal \N__50103\ : std_logic;
signal \N__50100\ : std_logic;
signal \N__50091\ : std_logic;
signal \N__50088\ : std_logic;
signal \N__50087\ : std_logic;
signal \N__50084\ : std_logic;
signal \N__50081\ : std_logic;
signal \N__50080\ : std_logic;
signal \N__50077\ : std_logic;
signal \N__50076\ : std_logic;
signal \N__50073\ : std_logic;
signal \N__50070\ : std_logic;
signal \N__50067\ : std_logic;
signal \N__50064\ : std_logic;
signal \N__50061\ : std_logic;
signal \N__50058\ : std_logic;
signal \N__50053\ : std_logic;
signal \N__50052\ : std_logic;
signal \N__50051\ : std_logic;
signal \N__50050\ : std_logic;
signal \N__50049\ : std_logic;
signal \N__50046\ : std_logic;
signal \N__50043\ : std_logic;
signal \N__50040\ : std_logic;
signal \N__50037\ : std_logic;
signal \N__50030\ : std_logic;
signal \N__50019\ : std_logic;
signal \N__50016\ : std_logic;
signal \N__50015\ : std_logic;
signal \N__50012\ : std_logic;
signal \N__50009\ : std_logic;
signal \N__50004\ : std_logic;
signal \N__50001\ : std_logic;
signal \N__49998\ : std_logic;
signal \N__49997\ : std_logic;
signal \N__49994\ : std_logic;
signal \N__49991\ : std_logic;
signal \N__49986\ : std_logic;
signal \N__49983\ : std_logic;
signal \N__49980\ : std_logic;
signal \N__49977\ : std_logic;
signal \N__49974\ : std_logic;
signal \N__49971\ : std_logic;
signal \N__49968\ : std_logic;
signal \N__49965\ : std_logic;
signal \N__49962\ : std_logic;
signal \N__49961\ : std_logic;
signal \N__49958\ : std_logic;
signal \N__49955\ : std_logic;
signal \N__49952\ : std_logic;
signal \N__49949\ : std_logic;
signal \N__49948\ : std_logic;
signal \N__49943\ : std_logic;
signal \N__49940\ : std_logic;
signal \N__49935\ : std_logic;
signal \N__49932\ : std_logic;
signal \N__49929\ : std_logic;
signal \N__49926\ : std_logic;
signal \N__49923\ : std_logic;
signal \N__49920\ : std_logic;
signal \N__49917\ : std_logic;
signal \N__49914\ : std_logic;
signal \N__49911\ : std_logic;
signal \N__49908\ : std_logic;
signal \N__49905\ : std_logic;
signal \N__49902\ : std_logic;
signal \N__49899\ : std_logic;
signal \N__49896\ : std_logic;
signal \N__49893\ : std_logic;
signal \N__49890\ : std_logic;
signal \N__49887\ : std_logic;
signal \N__49884\ : std_logic;
signal \N__49881\ : std_logic;
signal \N__49878\ : std_logic;
signal \N__49875\ : std_logic;
signal \N__49872\ : std_logic;
signal \N__49869\ : std_logic;
signal \N__49866\ : std_logic;
signal \N__49863\ : std_logic;
signal \N__49860\ : std_logic;
signal \N__49857\ : std_logic;
signal \N__49854\ : std_logic;
signal \N__49851\ : std_logic;
signal \N__49848\ : std_logic;
signal \N__49845\ : std_logic;
signal \N__49842\ : std_logic;
signal \N__49839\ : std_logic;
signal \N__49836\ : std_logic;
signal \N__49833\ : std_logic;
signal \N__49832\ : std_logic;
signal \N__49829\ : std_logic;
signal \N__49826\ : std_logic;
signal \N__49823\ : std_logic;
signal \N__49820\ : std_logic;
signal \N__49819\ : std_logic;
signal \N__49816\ : std_logic;
signal \N__49813\ : std_logic;
signal \N__49810\ : std_logic;
signal \N__49803\ : std_logic;
signal \N__49800\ : std_logic;
signal \N__49797\ : std_logic;
signal \N__49794\ : std_logic;
signal \N__49791\ : std_logic;
signal \N__49788\ : std_logic;
signal \N__49785\ : std_logic;
signal \N__49782\ : std_logic;
signal \N__49779\ : std_logic;
signal \N__49776\ : std_logic;
signal \N__49773\ : std_logic;
signal \N__49770\ : std_logic;
signal \N__49767\ : std_logic;
signal \N__49764\ : std_logic;
signal \N__49761\ : std_logic;
signal \N__49758\ : std_logic;
signal \N__49755\ : std_logic;
signal \N__49752\ : std_logic;
signal \N__49751\ : std_logic;
signal \N__49748\ : std_logic;
signal \N__49747\ : std_logic;
signal \N__49744\ : std_logic;
signal \N__49741\ : std_logic;
signal \N__49738\ : std_logic;
signal \N__49735\ : std_logic;
signal \N__49732\ : std_logic;
signal \N__49729\ : std_logic;
signal \N__49726\ : std_logic;
signal \N__49719\ : std_logic;
signal \N__49718\ : std_logic;
signal \N__49715\ : std_logic;
signal \N__49712\ : std_logic;
signal \N__49709\ : std_logic;
signal \N__49706\ : std_logic;
signal \N__49703\ : std_logic;
signal \N__49700\ : std_logic;
signal \N__49697\ : std_logic;
signal \N__49694\ : std_logic;
signal \N__49693\ : std_logic;
signal \N__49690\ : std_logic;
signal \N__49687\ : std_logic;
signal \N__49684\ : std_logic;
signal \N__49677\ : std_logic;
signal \N__49676\ : std_logic;
signal \N__49673\ : std_logic;
signal \N__49670\ : std_logic;
signal \N__49669\ : std_logic;
signal \N__49666\ : std_logic;
signal \N__49663\ : std_logic;
signal \N__49660\ : std_logic;
signal \N__49657\ : std_logic;
signal \N__49654\ : std_logic;
signal \N__49651\ : std_logic;
signal \N__49648\ : std_logic;
signal \N__49641\ : std_logic;
signal \N__49638\ : std_logic;
signal \N__49637\ : std_logic;
signal \N__49636\ : std_logic;
signal \N__49633\ : std_logic;
signal \N__49630\ : std_logic;
signal \N__49627\ : std_logic;
signal \N__49624\ : std_logic;
signal \N__49621\ : std_logic;
signal \N__49618\ : std_logic;
signal \N__49615\ : std_logic;
signal \N__49612\ : std_logic;
signal \N__49609\ : std_logic;
signal \N__49602\ : std_logic;
signal \N__49599\ : std_logic;
signal \N__49596\ : std_logic;
signal \N__49593\ : std_logic;
signal \N__49590\ : std_logic;
signal \N__49587\ : std_logic;
signal \N__49584\ : std_logic;
signal \N__49581\ : std_logic;
signal \N__49578\ : std_logic;
signal \N__49575\ : std_logic;
signal \N__49572\ : std_logic;
signal \N__49569\ : std_logic;
signal \N__49566\ : std_logic;
signal \N__49563\ : std_logic;
signal \N__49560\ : std_logic;
signal \N__49557\ : std_logic;
signal \N__49554\ : std_logic;
signal \N__49551\ : std_logic;
signal \N__49548\ : std_logic;
signal \N__49545\ : std_logic;
signal \N__49542\ : std_logic;
signal \N__49539\ : std_logic;
signal \N__49536\ : std_logic;
signal \N__49533\ : std_logic;
signal \N__49530\ : std_logic;
signal \N__49527\ : std_logic;
signal \N__49524\ : std_logic;
signal \N__49521\ : std_logic;
signal \N__49518\ : std_logic;
signal \N__49515\ : std_logic;
signal \N__49512\ : std_logic;
signal \N__49509\ : std_logic;
signal \N__49506\ : std_logic;
signal \N__49503\ : std_logic;
signal \N__49500\ : std_logic;
signal \N__49497\ : std_logic;
signal \N__49494\ : std_logic;
signal \N__49493\ : std_logic;
signal \N__49490\ : std_logic;
signal \N__49487\ : std_logic;
signal \N__49484\ : std_logic;
signal \N__49481\ : std_logic;
signal \N__49480\ : std_logic;
signal \N__49477\ : std_logic;
signal \N__49474\ : std_logic;
signal \N__49471\ : std_logic;
signal \N__49464\ : std_logic;
signal \N__49461\ : std_logic;
signal \N__49458\ : std_logic;
signal \N__49455\ : std_logic;
signal \N__49454\ : std_logic;
signal \N__49453\ : std_logic;
signal \N__49450\ : std_logic;
signal \N__49447\ : std_logic;
signal \N__49444\ : std_logic;
signal \N__49437\ : std_logic;
signal \N__49434\ : std_logic;
signal \N__49431\ : std_logic;
signal \N__49428\ : std_logic;
signal \N__49427\ : std_logic;
signal \N__49424\ : std_logic;
signal \N__49423\ : std_logic;
signal \N__49420\ : std_logic;
signal \N__49417\ : std_logic;
signal \N__49414\ : std_logic;
signal \N__49411\ : std_logic;
signal \N__49408\ : std_logic;
signal \N__49405\ : std_logic;
signal \N__49402\ : std_logic;
signal \N__49399\ : std_logic;
signal \N__49394\ : std_logic;
signal \N__49391\ : std_logic;
signal \N__49386\ : std_logic;
signal \N__49383\ : std_logic;
signal \N__49382\ : std_logic;
signal \N__49379\ : std_logic;
signal \N__49378\ : std_logic;
signal \N__49375\ : std_logic;
signal \N__49372\ : std_logic;
signal \N__49369\ : std_logic;
signal \N__49366\ : std_logic;
signal \N__49363\ : std_logic;
signal \N__49360\ : std_logic;
signal \N__49357\ : std_logic;
signal \N__49354\ : std_logic;
signal \N__49349\ : std_logic;
signal \N__49344\ : std_logic;
signal \N__49341\ : std_logic;
signal \N__49340\ : std_logic;
signal \N__49339\ : std_logic;
signal \N__49336\ : std_logic;
signal \N__49333\ : std_logic;
signal \N__49330\ : std_logic;
signal \N__49327\ : std_logic;
signal \N__49324\ : std_logic;
signal \N__49321\ : std_logic;
signal \N__49318\ : std_logic;
signal \N__49313\ : std_logic;
signal \N__49308\ : std_logic;
signal \N__49307\ : std_logic;
signal \N__49304\ : std_logic;
signal \N__49301\ : std_logic;
signal \N__49298\ : std_logic;
signal \N__49295\ : std_logic;
signal \N__49292\ : std_logic;
signal \N__49289\ : std_logic;
signal \N__49286\ : std_logic;
signal \N__49285\ : std_logic;
signal \N__49282\ : std_logic;
signal \N__49279\ : std_logic;
signal \N__49276\ : std_logic;
signal \N__49269\ : std_logic;
signal \N__49268\ : std_logic;
signal \N__49265\ : std_logic;
signal \N__49262\ : std_logic;
signal \N__49259\ : std_logic;
signal \N__49256\ : std_logic;
signal \N__49255\ : std_logic;
signal \N__49252\ : std_logic;
signal \N__49249\ : std_logic;
signal \N__49246\ : std_logic;
signal \N__49241\ : std_logic;
signal \N__49238\ : std_logic;
signal \N__49233\ : std_logic;
signal \N__49230\ : std_logic;
signal \N__49227\ : std_logic;
signal \N__49224\ : std_logic;
signal \N__49221\ : std_logic;
signal \N__49218\ : std_logic;
signal \N__49215\ : std_logic;
signal \N__49212\ : std_logic;
signal \N__49209\ : std_logic;
signal \N__49206\ : std_logic;
signal \N__49203\ : std_logic;
signal \N__49200\ : std_logic;
signal \N__49197\ : std_logic;
signal \N__49194\ : std_logic;
signal \N__49191\ : std_logic;
signal \N__49188\ : std_logic;
signal \N__49185\ : std_logic;
signal \N__49182\ : std_logic;
signal \N__49179\ : std_logic;
signal \N__49176\ : std_logic;
signal \N__49173\ : std_logic;
signal \N__49170\ : std_logic;
signal \N__49167\ : std_logic;
signal \N__49164\ : std_logic;
signal \N__49163\ : std_logic;
signal \N__49160\ : std_logic;
signal \N__49157\ : std_logic;
signal \N__49156\ : std_logic;
signal \N__49153\ : std_logic;
signal \N__49148\ : std_logic;
signal \N__49143\ : std_logic;
signal \N__49140\ : std_logic;
signal \N__49137\ : std_logic;
signal \N__49134\ : std_logic;
signal \N__49131\ : std_logic;
signal \N__49128\ : std_logic;
signal \N__49125\ : std_logic;
signal \N__49122\ : std_logic;
signal \N__49119\ : std_logic;
signal \N__49116\ : std_logic;
signal \N__49113\ : std_logic;
signal \N__49110\ : std_logic;
signal \N__49107\ : std_logic;
signal \N__49104\ : std_logic;
signal \N__49101\ : std_logic;
signal \N__49098\ : std_logic;
signal \N__49095\ : std_logic;
signal \N__49094\ : std_logic;
signal \N__49093\ : std_logic;
signal \N__49090\ : std_logic;
signal \N__49087\ : std_logic;
signal \N__49084\ : std_logic;
signal \N__49083\ : std_logic;
signal \N__49080\ : std_logic;
signal \N__49075\ : std_logic;
signal \N__49072\ : std_logic;
signal \N__49071\ : std_logic;
signal \N__49064\ : std_logic;
signal \N__49063\ : std_logic;
signal \N__49060\ : std_logic;
signal \N__49059\ : std_logic;
signal \N__49056\ : std_logic;
signal \N__49053\ : std_logic;
signal \N__49050\ : std_logic;
signal \N__49047\ : std_logic;
signal \N__49044\ : std_logic;
signal \N__49041\ : std_logic;
signal \N__49038\ : std_logic;
signal \N__49035\ : std_logic;
signal \N__49034\ : std_logic;
signal \N__49033\ : std_logic;
signal \N__49028\ : std_logic;
signal \N__49023\ : std_logic;
signal \N__49020\ : std_logic;
signal \N__49017\ : std_logic;
signal \N__49008\ : std_logic;
signal \N__49005\ : std_logic;
signal \N__49004\ : std_logic;
signal \N__49003\ : std_logic;
signal \N__49000\ : std_logic;
signal \N__48997\ : std_logic;
signal \N__48994\ : std_logic;
signal \N__48991\ : std_logic;
signal \N__48988\ : std_logic;
signal \N__48985\ : std_logic;
signal \N__48982\ : std_logic;
signal \N__48975\ : std_logic;
signal \N__48974\ : std_logic;
signal \N__48971\ : std_logic;
signal \N__48968\ : std_logic;
signal \N__48965\ : std_logic;
signal \N__48964\ : std_logic;
signal \N__48961\ : std_logic;
signal \N__48958\ : std_logic;
signal \N__48955\ : std_logic;
signal \N__48950\ : std_logic;
signal \N__48945\ : std_logic;
signal \N__48942\ : std_logic;
signal \N__48939\ : std_logic;
signal \N__48936\ : std_logic;
signal \N__48935\ : std_logic;
signal \N__48934\ : std_logic;
signal \N__48931\ : std_logic;
signal \N__48926\ : std_logic;
signal \N__48921\ : std_logic;
signal \N__48918\ : std_logic;
signal \N__48915\ : std_logic;
signal \N__48914\ : std_logic;
signal \N__48911\ : std_logic;
signal \N__48910\ : std_logic;
signal \N__48907\ : std_logic;
signal \N__48904\ : std_logic;
signal \N__48901\ : std_logic;
signal \N__48898\ : std_logic;
signal \N__48891\ : std_logic;
signal \N__48888\ : std_logic;
signal \N__48885\ : std_logic;
signal \N__48882\ : std_logic;
signal \N__48879\ : std_logic;
signal \N__48878\ : std_logic;
signal \N__48875\ : std_logic;
signal \N__48872\ : std_logic;
signal \N__48867\ : std_logic;
signal \N__48866\ : std_logic;
signal \N__48863\ : std_logic;
signal \N__48862\ : std_logic;
signal \N__48859\ : std_logic;
signal \N__48856\ : std_logic;
signal \N__48853\ : std_logic;
signal \N__48848\ : std_logic;
signal \N__48845\ : std_logic;
signal \N__48842\ : std_logic;
signal \N__48837\ : std_logic;
signal \N__48834\ : std_logic;
signal \N__48831\ : std_logic;
signal \N__48828\ : std_logic;
signal \N__48825\ : std_logic;
signal \N__48822\ : std_logic;
signal \N__48819\ : std_logic;
signal \N__48816\ : std_logic;
signal \N__48813\ : std_logic;
signal \N__48810\ : std_logic;
signal \N__48807\ : std_logic;
signal \N__48804\ : std_logic;
signal \N__48801\ : std_logic;
signal \N__48798\ : std_logic;
signal \N__48795\ : std_logic;
signal \N__48792\ : std_logic;
signal \N__48789\ : std_logic;
signal \N__48786\ : std_logic;
signal \N__48783\ : std_logic;
signal \N__48780\ : std_logic;
signal \N__48777\ : std_logic;
signal \N__48774\ : std_logic;
signal \N__48771\ : std_logic;
signal \N__48768\ : std_logic;
signal \N__48765\ : std_logic;
signal \N__48762\ : std_logic;
signal \N__48759\ : std_logic;
signal \N__48756\ : std_logic;
signal \N__48753\ : std_logic;
signal \N__48750\ : std_logic;
signal \N__48749\ : std_logic;
signal \N__48746\ : std_logic;
signal \N__48745\ : std_logic;
signal \N__48742\ : std_logic;
signal \N__48739\ : std_logic;
signal \N__48736\ : std_logic;
signal \N__48733\ : std_logic;
signal \N__48726\ : std_logic;
signal \N__48725\ : std_logic;
signal \N__48724\ : std_logic;
signal \N__48723\ : std_logic;
signal \N__48722\ : std_logic;
signal \N__48711\ : std_logic;
signal \N__48708\ : std_logic;
signal \N__48705\ : std_logic;
signal \N__48702\ : std_logic;
signal \N__48701\ : std_logic;
signal \N__48698\ : std_logic;
signal \N__48695\ : std_logic;
signal \N__48694\ : std_logic;
signal \N__48691\ : std_logic;
signal \N__48686\ : std_logic;
signal \N__48681\ : std_logic;
signal \N__48678\ : std_logic;
signal \N__48677\ : std_logic;
signal \N__48674\ : std_logic;
signal \N__48671\ : std_logic;
signal \N__48670\ : std_logic;
signal \N__48667\ : std_logic;
signal \N__48664\ : std_logic;
signal \N__48661\ : std_logic;
signal \N__48654\ : std_logic;
signal \N__48653\ : std_logic;
signal \N__48652\ : std_logic;
signal \N__48651\ : std_logic;
signal \N__48642\ : std_logic;
signal \N__48641\ : std_logic;
signal \N__48640\ : std_logic;
signal \N__48639\ : std_logic;
signal \N__48638\ : std_logic;
signal \N__48635\ : std_logic;
signal \N__48626\ : std_logic;
signal \N__48621\ : std_logic;
signal \N__48618\ : std_logic;
signal \N__48617\ : std_logic;
signal \N__48616\ : std_logic;
signal \N__48613\ : std_logic;
signal \N__48610\ : std_logic;
signal \N__48607\ : std_logic;
signal \N__48600\ : std_logic;
signal \N__48597\ : std_logic;
signal \N__48594\ : std_logic;
signal \N__48591\ : std_logic;
signal \N__48588\ : std_logic;
signal \N__48585\ : std_logic;
signal \N__48582\ : std_logic;
signal \N__48581\ : std_logic;
signal \N__48578\ : std_logic;
signal \N__48575\ : std_logic;
signal \N__48572\ : std_logic;
signal \N__48569\ : std_logic;
signal \N__48566\ : std_logic;
signal \N__48565\ : std_logic;
signal \N__48562\ : std_logic;
signal \N__48559\ : std_logic;
signal \N__48556\ : std_logic;
signal \N__48551\ : std_logic;
signal \N__48548\ : std_logic;
signal \N__48545\ : std_logic;
signal \N__48542\ : std_logic;
signal \N__48537\ : std_logic;
signal \N__48534\ : std_logic;
signal \N__48531\ : std_logic;
signal \N__48528\ : std_logic;
signal \N__48525\ : std_logic;
signal \N__48522\ : std_logic;
signal \N__48519\ : std_logic;
signal \N__48516\ : std_logic;
signal \N__48513\ : std_logic;
signal \N__48510\ : std_logic;
signal \N__48507\ : std_logic;
signal \N__48504\ : std_logic;
signal \N__48501\ : std_logic;
signal \N__48498\ : std_logic;
signal \N__48495\ : std_logic;
signal \N__48492\ : std_logic;
signal \N__48489\ : std_logic;
signal \N__48486\ : std_logic;
signal \N__48483\ : std_logic;
signal \N__48482\ : std_logic;
signal \N__48479\ : std_logic;
signal \N__48478\ : std_logic;
signal \N__48475\ : std_logic;
signal \N__48472\ : std_logic;
signal \N__48469\ : std_logic;
signal \N__48462\ : std_logic;
signal \N__48459\ : std_logic;
signal \N__48458\ : std_logic;
signal \N__48457\ : std_logic;
signal \N__48454\ : std_logic;
signal \N__48451\ : std_logic;
signal \N__48448\ : std_logic;
signal \N__48445\ : std_logic;
signal \N__48438\ : std_logic;
signal \N__48435\ : std_logic;
signal \N__48434\ : std_logic;
signal \N__48431\ : std_logic;
signal \N__48430\ : std_logic;
signal \N__48427\ : std_logic;
signal \N__48424\ : std_logic;
signal \N__48421\ : std_logic;
signal \N__48414\ : std_logic;
signal \N__48411\ : std_logic;
signal \N__48410\ : std_logic;
signal \N__48409\ : std_logic;
signal \N__48406\ : std_logic;
signal \N__48401\ : std_logic;
signal \N__48396\ : std_logic;
signal \N__48393\ : std_logic;
signal \N__48392\ : std_logic;
signal \N__48391\ : std_logic;
signal \N__48388\ : std_logic;
signal \N__48383\ : std_logic;
signal \N__48378\ : std_logic;
signal \N__48375\ : std_logic;
signal \N__48374\ : std_logic;
signal \N__48373\ : std_logic;
signal \N__48370\ : std_logic;
signal \N__48365\ : std_logic;
signal \N__48360\ : std_logic;
signal \N__48357\ : std_logic;
signal \N__48356\ : std_logic;
signal \N__48355\ : std_logic;
signal \N__48352\ : std_logic;
signal \N__48349\ : std_logic;
signal \N__48346\ : std_logic;
signal \N__48343\ : std_logic;
signal \N__48340\ : std_logic;
signal \N__48333\ : std_logic;
signal \N__48330\ : std_logic;
signal \N__48329\ : std_logic;
signal \N__48326\ : std_logic;
signal \N__48325\ : std_logic;
signal \N__48322\ : std_logic;
signal \N__48317\ : std_logic;
signal \N__48314\ : std_logic;
signal \N__48311\ : std_logic;
signal \N__48310\ : std_logic;
signal \N__48307\ : std_logic;
signal \N__48304\ : std_logic;
signal \N__48301\ : std_logic;
signal \N__48294\ : std_logic;
signal \N__48293\ : std_logic;
signal \N__48292\ : std_logic;
signal \N__48291\ : std_logic;
signal \N__48290\ : std_logic;
signal \N__48287\ : std_logic;
signal \N__48284\ : std_logic;
signal \N__48281\ : std_logic;
signal \N__48278\ : std_logic;
signal \N__48275\ : std_logic;
signal \N__48272\ : std_logic;
signal \N__48263\ : std_logic;
signal \N__48262\ : std_logic;
signal \N__48259\ : std_logic;
signal \N__48258\ : std_logic;
signal \N__48257\ : std_logic;
signal \N__48256\ : std_logic;
signal \N__48253\ : std_logic;
signal \N__48250\ : std_logic;
signal \N__48247\ : std_logic;
signal \N__48244\ : std_logic;
signal \N__48241\ : std_logic;
signal \N__48238\ : std_logic;
signal \N__48235\ : std_logic;
signal \N__48222\ : std_logic;
signal \N__48221\ : std_logic;
signal \N__48220\ : std_logic;
signal \N__48219\ : std_logic;
signal \N__48216\ : std_logic;
signal \N__48213\ : std_logic;
signal \N__48210\ : std_logic;
signal \N__48209\ : std_logic;
signal \N__48206\ : std_logic;
signal \N__48205\ : std_logic;
signal \N__48196\ : std_logic;
signal \N__48195\ : std_logic;
signal \N__48190\ : std_logic;
signal \N__48187\ : std_logic;
signal \N__48184\ : std_logic;
signal \N__48183\ : std_logic;
signal \N__48182\ : std_logic;
signal \N__48181\ : std_logic;
signal \N__48174\ : std_logic;
signal \N__48167\ : std_logic;
signal \N__48162\ : std_logic;
signal \N__48159\ : std_logic;
signal \N__48158\ : std_logic;
signal \N__48157\ : std_logic;
signal \N__48156\ : std_logic;
signal \N__48153\ : std_logic;
signal \N__48150\ : std_logic;
signal \N__48147\ : std_logic;
signal \N__48144\ : std_logic;
signal \N__48141\ : std_logic;
signal \N__48140\ : std_logic;
signal \N__48133\ : std_logic;
signal \N__48132\ : std_logic;
signal \N__48129\ : std_logic;
signal \N__48126\ : std_logic;
signal \N__48123\ : std_logic;
signal \N__48120\ : std_logic;
signal \N__48111\ : std_logic;
signal \N__48108\ : std_logic;
signal \N__48107\ : std_logic;
signal \N__48106\ : std_logic;
signal \N__48105\ : std_logic;
signal \N__48102\ : std_logic;
signal \N__48099\ : std_logic;
signal \N__48096\ : std_logic;
signal \N__48093\ : std_logic;
signal \N__48090\ : std_logic;
signal \N__48085\ : std_logic;
signal \N__48082\ : std_logic;
signal \N__48081\ : std_logic;
signal \N__48080\ : std_logic;
signal \N__48077\ : std_logic;
signal \N__48074\ : std_logic;
signal \N__48071\ : std_logic;
signal \N__48066\ : std_logic;
signal \N__48057\ : std_logic;
signal \N__48056\ : std_logic;
signal \N__48053\ : std_logic;
signal \N__48050\ : std_logic;
signal \N__48049\ : std_logic;
signal \N__48048\ : std_logic;
signal \N__48045\ : std_logic;
signal \N__48042\ : std_logic;
signal \N__48039\ : std_logic;
signal \N__48036\ : std_logic;
signal \N__48033\ : std_logic;
signal \N__48032\ : std_logic;
signal \N__48029\ : std_logic;
signal \N__48024\ : std_logic;
signal \N__48021\ : std_logic;
signal \N__48020\ : std_logic;
signal \N__48017\ : std_logic;
signal \N__48014\ : std_logic;
signal \N__48009\ : std_logic;
signal \N__48006\ : std_logic;
signal \N__47997\ : std_logic;
signal \N__47996\ : std_logic;
signal \N__47995\ : std_logic;
signal \N__47994\ : std_logic;
signal \N__47993\ : std_logic;
signal \N__47992\ : std_logic;
signal \N__47991\ : std_logic;
signal \N__47990\ : std_logic;
signal \N__47989\ : std_logic;
signal \N__47988\ : std_logic;
signal \N__47987\ : std_logic;
signal \N__47986\ : std_logic;
signal \N__47985\ : std_logic;
signal \N__47984\ : std_logic;
signal \N__47983\ : std_logic;
signal \N__47982\ : std_logic;
signal \N__47981\ : std_logic;
signal \N__47980\ : std_logic;
signal \N__47979\ : std_logic;
signal \N__47978\ : std_logic;
signal \N__47937\ : std_logic;
signal \N__47934\ : std_logic;
signal \N__47931\ : std_logic;
signal \N__47928\ : std_logic;
signal \N__47925\ : std_logic;
signal \N__47922\ : std_logic;
signal \N__47921\ : std_logic;
signal \N__47918\ : std_logic;
signal \N__47915\ : std_logic;
signal \N__47914\ : std_logic;
signal \N__47913\ : std_logic;
signal \N__47912\ : std_logic;
signal \N__47907\ : std_logic;
signal \N__47904\ : std_logic;
signal \N__47899\ : std_logic;
signal \N__47892\ : std_logic;
signal \N__47889\ : std_logic;
signal \N__47886\ : std_logic;
signal \N__47883\ : std_logic;
signal \N__47882\ : std_logic;
signal \N__47881\ : std_logic;
signal \N__47880\ : std_logic;
signal \N__47879\ : std_logic;
signal \N__47878\ : std_logic;
signal \N__47877\ : std_logic;
signal \N__47876\ : std_logic;
signal \N__47875\ : std_logic;
signal \N__47874\ : std_logic;
signal \N__47873\ : std_logic;
signal \N__47872\ : std_logic;
signal \N__47871\ : std_logic;
signal \N__47870\ : std_logic;
signal \N__47869\ : std_logic;
signal \N__47868\ : std_logic;
signal \N__47867\ : std_logic;
signal \N__47866\ : std_logic;
signal \N__47865\ : std_logic;
signal \N__47864\ : std_logic;
signal \N__47863\ : std_logic;
signal \N__47860\ : std_logic;
signal \N__47859\ : std_logic;
signal \N__47858\ : std_logic;
signal \N__47857\ : std_logic;
signal \N__47856\ : std_logic;
signal \N__47855\ : std_logic;
signal \N__47854\ : std_logic;
signal \N__47853\ : std_logic;
signal \N__47852\ : std_logic;
signal \N__47851\ : std_logic;
signal \N__47850\ : std_logic;
signal \N__47849\ : std_logic;
signal \N__47848\ : std_logic;
signal \N__47847\ : std_logic;
signal \N__47846\ : std_logic;
signal \N__47845\ : std_logic;
signal \N__47844\ : std_logic;
signal \N__47843\ : std_logic;
signal \N__47842\ : std_logic;
signal \N__47833\ : std_logic;
signal \N__47828\ : std_logic;
signal \N__47823\ : std_logic;
signal \N__47820\ : std_logic;
signal \N__47815\ : std_logic;
signal \N__47814\ : std_logic;
signal \N__47813\ : std_logic;
signal \N__47812\ : std_logic;
signal \N__47811\ : std_logic;
signal \N__47810\ : std_logic;
signal \N__47803\ : std_logic;
signal \N__47798\ : std_logic;
signal \N__47795\ : std_logic;
signal \N__47788\ : std_logic;
signal \N__47785\ : std_logic;
signal \N__47778\ : std_logic;
signal \N__47771\ : std_logic;
signal \N__47764\ : std_logic;
signal \N__47759\ : std_logic;
signal \N__47756\ : std_logic;
signal \N__47743\ : std_logic;
signal \N__47742\ : std_logic;
signal \N__47741\ : std_logic;
signal \N__47732\ : std_logic;
signal \N__47731\ : std_logic;
signal \N__47730\ : std_logic;
signal \N__47729\ : std_logic;
signal \N__47728\ : std_logic;
signal \N__47727\ : std_logic;
signal \N__47726\ : std_logic;
signal \N__47725\ : std_logic;
signal \N__47724\ : std_logic;
signal \N__47721\ : std_logic;
signal \N__47716\ : std_logic;
signal \N__47711\ : std_logic;
signal \N__47708\ : std_logic;
signal \N__47707\ : std_logic;
signal \N__47706\ : std_logic;
signal \N__47703\ : std_logic;
signal \N__47696\ : std_logic;
signal \N__47681\ : std_logic;
signal \N__47676\ : std_logic;
signal \N__47673\ : std_logic;
signal \N__47664\ : std_logic;
signal \N__47655\ : std_logic;
signal \N__47654\ : std_logic;
signal \N__47653\ : std_logic;
signal \N__47652\ : std_logic;
signal \N__47651\ : std_logic;
signal \N__47650\ : std_logic;
signal \N__47649\ : std_logic;
signal \N__47648\ : std_logic;
signal \N__47647\ : std_logic;
signal \N__47646\ : std_logic;
signal \N__47645\ : std_logic;
signal \N__47644\ : std_logic;
signal \N__47639\ : std_logic;
signal \N__47634\ : std_logic;
signal \N__47629\ : std_logic;
signal \N__47620\ : std_logic;
signal \N__47613\ : std_logic;
signal \N__47602\ : std_logic;
signal \N__47591\ : std_logic;
signal \N__47588\ : std_logic;
signal \N__47571\ : std_logic;
signal \N__47568\ : std_logic;
signal \N__47565\ : std_logic;
signal \N__47564\ : std_logic;
signal \N__47563\ : std_logic;
signal \N__47562\ : std_logic;
signal \N__47557\ : std_logic;
signal \N__47552\ : std_logic;
signal \N__47547\ : std_logic;
signal \N__47546\ : std_logic;
signal \N__47545\ : std_logic;
signal \N__47538\ : std_logic;
signal \N__47535\ : std_logic;
signal \N__47532\ : std_logic;
signal \N__47529\ : std_logic;
signal \N__47526\ : std_logic;
signal \N__47523\ : std_logic;
signal \N__47520\ : std_logic;
signal \N__47517\ : std_logic;
signal \N__47514\ : std_logic;
signal \N__47511\ : std_logic;
signal \N__47510\ : std_logic;
signal \N__47507\ : std_logic;
signal \N__47504\ : std_logic;
signal \N__47501\ : std_logic;
signal \N__47498\ : std_logic;
signal \N__47493\ : std_logic;
signal \N__47490\ : std_logic;
signal \N__47487\ : std_logic;
signal \N__47484\ : std_logic;
signal \N__47481\ : std_logic;
signal \N__47478\ : std_logic;
signal \N__47475\ : std_logic;
signal \N__47472\ : std_logic;
signal \N__47469\ : std_logic;
signal \N__47468\ : std_logic;
signal \N__47463\ : std_logic;
signal \N__47460\ : std_logic;
signal \N__47457\ : std_logic;
signal \N__47456\ : std_logic;
signal \N__47453\ : std_logic;
signal \N__47450\ : std_logic;
signal \N__47445\ : std_logic;
signal \N__47442\ : std_logic;
signal \N__47439\ : std_logic;
signal \N__47436\ : std_logic;
signal \N__47433\ : std_logic;
signal \N__47430\ : std_logic;
signal \N__47427\ : std_logic;
signal \N__47426\ : std_logic;
signal \N__47423\ : std_logic;
signal \N__47420\ : std_logic;
signal \N__47415\ : std_logic;
signal \N__47414\ : std_logic;
signal \N__47413\ : std_logic;
signal \N__47412\ : std_logic;
signal \N__47411\ : std_logic;
signal \N__47410\ : std_logic;
signal \N__47409\ : std_logic;
signal \N__47404\ : std_logic;
signal \N__47403\ : std_logic;
signal \N__47400\ : std_logic;
signal \N__47391\ : std_logic;
signal \N__47388\ : std_logic;
signal \N__47385\ : std_logic;
signal \N__47384\ : std_logic;
signal \N__47383\ : std_logic;
signal \N__47382\ : std_logic;
signal \N__47381\ : std_logic;
signal \N__47380\ : std_logic;
signal \N__47379\ : std_logic;
signal \N__47378\ : std_logic;
signal \N__47375\ : std_logic;
signal \N__47372\ : std_logic;
signal \N__47369\ : std_logic;
signal \N__47366\ : std_logic;
signal \N__47357\ : std_logic;
signal \N__47350\ : std_logic;
signal \N__47347\ : std_logic;
signal \N__47344\ : std_logic;
signal \N__47341\ : std_logic;
signal \N__47328\ : std_logic;
signal \N__47325\ : std_logic;
signal \N__47322\ : std_logic;
signal \N__47319\ : std_logic;
signal \N__47316\ : std_logic;
signal \N__47313\ : std_logic;
signal \N__47310\ : std_logic;
signal \N__47307\ : std_logic;
signal \N__47304\ : std_logic;
signal \N__47301\ : std_logic;
signal \N__47298\ : std_logic;
signal \N__47295\ : std_logic;
signal \N__47292\ : std_logic;
signal \N__47289\ : std_logic;
signal \N__47286\ : std_logic;
signal \N__47283\ : std_logic;
signal \N__47280\ : std_logic;
signal \N__47277\ : std_logic;
signal \N__47274\ : std_logic;
signal \N__47271\ : std_logic;
signal \N__47268\ : std_logic;
signal \N__47265\ : std_logic;
signal \N__47262\ : std_logic;
signal \N__47259\ : std_logic;
signal \N__47256\ : std_logic;
signal \N__47253\ : std_logic;
signal \N__47250\ : std_logic;
signal \N__47247\ : std_logic;
signal \N__47246\ : std_logic;
signal \N__47245\ : std_logic;
signal \N__47244\ : std_logic;
signal \N__47243\ : std_logic;
signal \N__47240\ : std_logic;
signal \N__47237\ : std_logic;
signal \N__47232\ : std_logic;
signal \N__47229\ : std_logic;
signal \N__47222\ : std_logic;
signal \N__47219\ : std_logic;
signal \N__47216\ : std_logic;
signal \N__47213\ : std_logic;
signal \N__47208\ : std_logic;
signal \N__47207\ : std_logic;
signal \N__47206\ : std_logic;
signal \N__47201\ : std_logic;
signal \N__47198\ : std_logic;
signal \N__47197\ : std_logic;
signal \N__47196\ : std_logic;
signal \N__47193\ : std_logic;
signal \N__47190\ : std_logic;
signal \N__47187\ : std_logic;
signal \N__47184\ : std_logic;
signal \N__47179\ : std_logic;
signal \N__47172\ : std_logic;
signal \N__47171\ : std_logic;
signal \N__47170\ : std_logic;
signal \N__47169\ : std_logic;
signal \N__47168\ : std_logic;
signal \N__47165\ : std_logic;
signal \N__47164\ : std_logic;
signal \N__47161\ : std_logic;
signal \N__47158\ : std_logic;
signal \N__47153\ : std_logic;
signal \N__47150\ : std_logic;
signal \N__47147\ : std_logic;
signal \N__47140\ : std_logic;
signal \N__47137\ : std_logic;
signal \N__47134\ : std_logic;
signal \N__47129\ : std_logic;
signal \N__47124\ : std_logic;
signal \N__47123\ : std_logic;
signal \N__47122\ : std_logic;
signal \N__47119\ : std_logic;
signal \N__47118\ : std_logic;
signal \N__47115\ : std_logic;
signal \N__47112\ : std_logic;
signal \N__47111\ : std_logic;
signal \N__47110\ : std_logic;
signal \N__47107\ : std_logic;
signal \N__47104\ : std_logic;
signal \N__47099\ : std_logic;
signal \N__47094\ : std_logic;
signal \N__47093\ : std_logic;
signal \N__47090\ : std_logic;
signal \N__47085\ : std_logic;
signal \N__47082\ : std_logic;
signal \N__47079\ : std_logic;
signal \N__47076\ : std_logic;
signal \N__47073\ : std_logic;
signal \N__47068\ : std_logic;
signal \N__47061\ : std_logic;
signal \N__47058\ : std_logic;
signal \N__47055\ : std_logic;
signal \N__47052\ : std_logic;
signal \N__47049\ : std_logic;
signal \N__47046\ : std_logic;
signal \N__47043\ : std_logic;
signal \N__47042\ : std_logic;
signal \N__47041\ : std_logic;
signal \N__47038\ : std_logic;
signal \N__47037\ : std_logic;
signal \N__47034\ : std_logic;
signal \N__47031\ : std_logic;
signal \N__47028\ : std_logic;
signal \N__47025\ : std_logic;
signal \N__47018\ : std_logic;
signal \N__47013\ : std_logic;
signal \N__47012\ : std_logic;
signal \N__47009\ : std_logic;
signal \N__47008\ : std_logic;
signal \N__47007\ : std_logic;
signal \N__47004\ : std_logic;
signal \N__47001\ : std_logic;
signal \N__46998\ : std_logic;
signal \N__46995\ : std_logic;
signal \N__46992\ : std_logic;
signal \N__46989\ : std_logic;
signal \N__46980\ : std_logic;
signal \N__46977\ : std_logic;
signal \N__46974\ : std_logic;
signal \N__46971\ : std_logic;
signal \N__46968\ : std_logic;
signal \N__46965\ : std_logic;
signal \N__46962\ : std_logic;
signal \N__46959\ : std_logic;
signal \N__46956\ : std_logic;
signal \N__46953\ : std_logic;
signal \N__46950\ : std_logic;
signal \N__46947\ : std_logic;
signal \N__46946\ : std_logic;
signal \N__46943\ : std_logic;
signal \N__46942\ : std_logic;
signal \N__46939\ : std_logic;
signal \N__46938\ : std_logic;
signal \N__46935\ : std_logic;
signal \N__46932\ : std_logic;
signal \N__46929\ : std_logic;
signal \N__46926\ : std_logic;
signal \N__46923\ : std_logic;
signal \N__46914\ : std_logic;
signal \N__46911\ : std_logic;
signal \N__46910\ : std_logic;
signal \N__46909\ : std_logic;
signal \N__46908\ : std_logic;
signal \N__46907\ : std_logic;
signal \N__46904\ : std_logic;
signal \N__46901\ : std_logic;
signal \N__46900\ : std_logic;
signal \N__46897\ : std_logic;
signal \N__46896\ : std_logic;
signal \N__46893\ : std_logic;
signal \N__46892\ : std_logic;
signal \N__46891\ : std_logic;
signal \N__46888\ : std_logic;
signal \N__46885\ : std_logic;
signal \N__46876\ : std_logic;
signal \N__46869\ : std_logic;
signal \N__46866\ : std_logic;
signal \N__46863\ : std_logic;
signal \N__46860\ : std_logic;
signal \N__46857\ : std_logic;
signal \N__46854\ : std_logic;
signal \N__46849\ : std_logic;
signal \N__46846\ : std_logic;
signal \N__46843\ : std_logic;
signal \N__46840\ : std_logic;
signal \N__46837\ : std_logic;
signal \N__46832\ : std_logic;
signal \N__46829\ : std_logic;
signal \N__46824\ : std_logic;
signal \N__46821\ : std_logic;
signal \N__46818\ : std_logic;
signal \N__46817\ : std_logic;
signal \N__46814\ : std_logic;
signal \N__46813\ : std_logic;
signal \N__46812\ : std_logic;
signal \N__46811\ : std_logic;
signal \N__46808\ : std_logic;
signal \N__46807\ : std_logic;
signal \N__46804\ : std_logic;
signal \N__46799\ : std_logic;
signal \N__46796\ : std_logic;
signal \N__46793\ : std_logic;
signal \N__46790\ : std_logic;
signal \N__46787\ : std_logic;
signal \N__46782\ : std_logic;
signal \N__46779\ : std_logic;
signal \N__46772\ : std_logic;
signal \N__46769\ : std_logic;
signal \N__46764\ : std_logic;
signal \N__46763\ : std_logic;
signal \N__46762\ : std_logic;
signal \N__46761\ : std_logic;
signal \N__46760\ : std_logic;
signal \N__46757\ : std_logic;
signal \N__46756\ : std_logic;
signal \N__46753\ : std_logic;
signal \N__46746\ : std_logic;
signal \N__46743\ : std_logic;
signal \N__46740\ : std_logic;
signal \N__46737\ : std_logic;
signal \N__46732\ : std_logic;
signal \N__46725\ : std_logic;
signal \N__46722\ : std_logic;
signal \N__46719\ : std_logic;
signal \N__46716\ : std_logic;
signal \N__46713\ : std_logic;
signal \N__46710\ : std_logic;
signal \N__46707\ : std_logic;
signal \N__46704\ : std_logic;
signal \N__46701\ : std_logic;
signal \N__46698\ : std_logic;
signal \N__46695\ : std_logic;
signal \N__46692\ : std_logic;
signal \N__46689\ : std_logic;
signal \N__46686\ : std_logic;
signal \N__46683\ : std_logic;
signal \N__46680\ : std_logic;
signal \N__46677\ : std_logic;
signal \N__46674\ : std_logic;
signal \N__46671\ : std_logic;
signal \N__46668\ : std_logic;
signal \N__46667\ : std_logic;
signal \N__46664\ : std_logic;
signal \N__46661\ : std_logic;
signal \N__46660\ : std_logic;
signal \N__46657\ : std_logic;
signal \N__46654\ : std_logic;
signal \N__46651\ : std_logic;
signal \N__46644\ : std_logic;
signal \N__46641\ : std_logic;
signal \N__46638\ : std_logic;
signal \N__46635\ : std_logic;
signal \N__46634\ : std_logic;
signal \N__46631\ : std_logic;
signal \N__46628\ : std_logic;
signal \N__46627\ : std_logic;
signal \N__46624\ : std_logic;
signal \N__46619\ : std_logic;
signal \N__46614\ : std_logic;
signal \N__46611\ : std_logic;
signal \N__46608\ : std_logic;
signal \N__46605\ : std_logic;
signal \N__46602\ : std_logic;
signal \N__46599\ : std_logic;
signal \N__46598\ : std_logic;
signal \N__46597\ : std_logic;
signal \N__46594\ : std_logic;
signal \N__46589\ : std_logic;
signal \N__46586\ : std_logic;
signal \N__46583\ : std_logic;
signal \N__46578\ : std_logic;
signal \N__46575\ : std_logic;
signal \N__46572\ : std_logic;
signal \N__46569\ : std_logic;
signal \N__46566\ : std_logic;
signal \N__46563\ : std_logic;
signal \N__46560\ : std_logic;
signal \N__46557\ : std_logic;
signal \N__46556\ : std_logic;
signal \N__46553\ : std_logic;
signal \N__46552\ : std_logic;
signal \N__46549\ : std_logic;
signal \N__46546\ : std_logic;
signal \N__46541\ : std_logic;
signal \N__46538\ : std_logic;
signal \N__46535\ : std_logic;
signal \N__46530\ : std_logic;
signal \N__46527\ : std_logic;
signal \N__46526\ : std_logic;
signal \N__46525\ : std_logic;
signal \N__46524\ : std_logic;
signal \N__46523\ : std_logic;
signal \N__46520\ : std_logic;
signal \N__46517\ : std_logic;
signal \N__46514\ : std_logic;
signal \N__46511\ : std_logic;
signal \N__46508\ : std_logic;
signal \N__46507\ : std_logic;
signal \N__46502\ : std_logic;
signal \N__46501\ : std_logic;
signal \N__46500\ : std_logic;
signal \N__46497\ : std_logic;
signal \N__46494\ : std_logic;
signal \N__46491\ : std_logic;
signal \N__46488\ : std_logic;
signal \N__46485\ : std_logic;
signal \N__46482\ : std_logic;
signal \N__46479\ : std_logic;
signal \N__46476\ : std_logic;
signal \N__46471\ : std_logic;
signal \N__46468\ : std_logic;
signal \N__46465\ : std_logic;
signal \N__46462\ : std_logic;
signal \N__46461\ : std_logic;
signal \N__46458\ : std_logic;
signal \N__46453\ : std_logic;
signal \N__46450\ : std_logic;
signal \N__46447\ : std_logic;
signal \N__46444\ : std_logic;
signal \N__46441\ : std_logic;
signal \N__46438\ : std_logic;
signal \N__46435\ : std_logic;
signal \N__46428\ : std_logic;
signal \N__46419\ : std_logic;
signal \N__46416\ : std_logic;
signal \N__46413\ : std_logic;
signal \N__46410\ : std_logic;
signal \N__46407\ : std_logic;
signal \N__46404\ : std_logic;
signal \N__46401\ : std_logic;
signal \N__46398\ : std_logic;
signal \N__46395\ : std_logic;
signal \N__46392\ : std_logic;
signal \N__46389\ : std_logic;
signal \N__46386\ : std_logic;
signal \N__46383\ : std_logic;
signal \N__46380\ : std_logic;
signal \N__46377\ : std_logic;
signal \N__46376\ : std_logic;
signal \N__46373\ : std_logic;
signal \N__46370\ : std_logic;
signal \N__46369\ : std_logic;
signal \N__46366\ : std_logic;
signal \N__46363\ : std_logic;
signal \N__46360\ : std_logic;
signal \N__46355\ : std_logic;
signal \N__46350\ : std_logic;
signal \N__46347\ : std_logic;
signal \N__46346\ : std_logic;
signal \N__46343\ : std_logic;
signal \N__46340\ : std_logic;
signal \N__46339\ : std_logic;
signal \N__46336\ : std_logic;
signal \N__46333\ : std_logic;
signal \N__46330\ : std_logic;
signal \N__46327\ : std_logic;
signal \N__46322\ : std_logic;
signal \N__46317\ : std_logic;
signal \N__46314\ : std_logic;
signal \N__46311\ : std_logic;
signal \N__46308\ : std_logic;
signal \N__46307\ : std_logic;
signal \N__46306\ : std_logic;
signal \N__46303\ : std_logic;
signal \N__46298\ : std_logic;
signal \N__46293\ : std_logic;
signal \N__46290\ : std_logic;
signal \N__46287\ : std_logic;
signal \N__46284\ : std_logic;
signal \N__46281\ : std_logic;
signal \N__46278\ : std_logic;
signal \N__46275\ : std_logic;
signal \N__46272\ : std_logic;
signal \N__46271\ : std_logic;
signal \N__46270\ : std_logic;
signal \N__46267\ : std_logic;
signal \N__46264\ : std_logic;
signal \N__46261\ : std_logic;
signal \N__46258\ : std_logic;
signal \N__46255\ : std_logic;
signal \N__46252\ : std_logic;
signal \N__46249\ : std_logic;
signal \N__46246\ : std_logic;
signal \N__46243\ : std_logic;
signal \N__46240\ : std_logic;
signal \N__46237\ : std_logic;
signal \N__46234\ : std_logic;
signal \N__46227\ : std_logic;
signal \N__46224\ : std_logic;
signal \N__46221\ : std_logic;
signal \N__46218\ : std_logic;
signal \N__46215\ : std_logic;
signal \N__46212\ : std_logic;
signal \N__46211\ : std_logic;
signal \N__46208\ : std_logic;
signal \N__46205\ : std_logic;
signal \N__46202\ : std_logic;
signal \N__46199\ : std_logic;
signal \N__46198\ : std_logic;
signal \N__46195\ : std_logic;
signal \N__46192\ : std_logic;
signal \N__46189\ : std_logic;
signal \N__46186\ : std_logic;
signal \N__46183\ : std_logic;
signal \N__46180\ : std_logic;
signal \N__46173\ : std_logic;
signal \N__46172\ : std_logic;
signal \N__46169\ : std_logic;
signal \N__46166\ : std_logic;
signal \N__46163\ : std_logic;
signal \N__46160\ : std_logic;
signal \N__46159\ : std_logic;
signal \N__46154\ : std_logic;
signal \N__46151\ : std_logic;
signal \N__46148\ : std_logic;
signal \N__46145\ : std_logic;
signal \N__46142\ : std_logic;
signal \N__46137\ : std_logic;
signal \N__46134\ : std_logic;
signal \N__46131\ : std_logic;
signal \N__46128\ : std_logic;
signal \N__46125\ : std_logic;
signal \N__46122\ : std_logic;
signal \N__46119\ : std_logic;
signal \N__46116\ : std_logic;
signal \N__46115\ : std_logic;
signal \N__46112\ : std_logic;
signal \N__46109\ : std_logic;
signal \N__46106\ : std_logic;
signal \N__46101\ : std_logic;
signal \N__46098\ : std_logic;
signal \N__46095\ : std_logic;
signal \N__46092\ : std_logic;
signal \N__46089\ : std_logic;
signal \N__46086\ : std_logic;
signal \N__46083\ : std_logic;
signal \N__46080\ : std_logic;
signal \N__46077\ : std_logic;
signal \N__46074\ : std_logic;
signal \N__46071\ : std_logic;
signal \N__46068\ : std_logic;
signal \N__46065\ : std_logic;
signal \N__46064\ : std_logic;
signal \N__46061\ : std_logic;
signal \N__46060\ : std_logic;
signal \N__46059\ : std_logic;
signal \N__46058\ : std_logic;
signal \N__46057\ : std_logic;
signal \N__46056\ : std_logic;
signal \N__46055\ : std_logic;
signal \N__46054\ : std_logic;
signal \N__46053\ : std_logic;
signal \N__46052\ : std_logic;
signal \N__46051\ : std_logic;
signal \N__46050\ : std_logic;
signal \N__46047\ : std_logic;
signal \N__46046\ : std_logic;
signal \N__46045\ : std_logic;
signal \N__46044\ : std_logic;
signal \N__46043\ : std_logic;
signal \N__46042\ : std_logic;
signal \N__46041\ : std_logic;
signal \N__46038\ : std_logic;
signal \N__46035\ : std_logic;
signal \N__46032\ : std_logic;
signal \N__46027\ : std_logic;
signal \N__46014\ : std_logic;
signal \N__46013\ : std_logic;
signal \N__46010\ : std_logic;
signal \N__46007\ : std_logic;
signal \N__45996\ : std_logic;
signal \N__45993\ : std_logic;
signal \N__45992\ : std_logic;
signal \N__45991\ : std_logic;
signal \N__45990\ : std_logic;
signal \N__45989\ : std_logic;
signal \N__45984\ : std_logic;
signal \N__45977\ : std_logic;
signal \N__45974\ : std_logic;
signal \N__45967\ : std_logic;
signal \N__45962\ : std_logic;
signal \N__45959\ : std_logic;
signal \N__45954\ : std_logic;
signal \N__45949\ : std_logic;
signal \N__45944\ : std_logic;
signal \N__45941\ : std_logic;
signal \N__45934\ : std_logic;
signal \N__45931\ : std_logic;
signal \N__45926\ : std_logic;
signal \N__45921\ : std_logic;
signal \N__45920\ : std_logic;
signal \N__45919\ : std_logic;
signal \N__45916\ : std_logic;
signal \N__45915\ : std_logic;
signal \N__45912\ : std_logic;
signal \N__45909\ : std_logic;
signal \N__45908\ : std_logic;
signal \N__45907\ : std_logic;
signal \N__45906\ : std_logic;
signal \N__45905\ : std_logic;
signal \N__45904\ : std_logic;
signal \N__45903\ : std_logic;
signal \N__45902\ : std_logic;
signal \N__45899\ : std_logic;
signal \N__45896\ : std_logic;
signal \N__45879\ : std_logic;
signal \N__45876\ : std_logic;
signal \N__45875\ : std_logic;
signal \N__45874\ : std_logic;
signal \N__45873\ : std_logic;
signal \N__45872\ : std_logic;
signal \N__45871\ : std_logic;
signal \N__45870\ : std_logic;
signal \N__45869\ : std_logic;
signal \N__45868\ : std_logic;
signal \N__45867\ : std_logic;
signal \N__45866\ : std_logic;
signal \N__45863\ : std_logic;
signal \N__45860\ : std_logic;
signal \N__45857\ : std_logic;
signal \N__45854\ : std_logic;
signal \N__45843\ : std_logic;
signal \N__45842\ : std_logic;
signal \N__45839\ : std_logic;
signal \N__45836\ : std_logic;
signal \N__45833\ : std_logic;
signal \N__45832\ : std_logic;
signal \N__45831\ : std_logic;
signal \N__45826\ : std_logic;
signal \N__45819\ : std_logic;
signal \N__45814\ : std_logic;
signal \N__45811\ : std_logic;
signal \N__45808\ : std_logic;
signal \N__45805\ : std_logic;
signal \N__45798\ : std_logic;
signal \N__45795\ : std_logic;
signal \N__45788\ : std_logic;
signal \N__45781\ : std_logic;
signal \N__45776\ : std_logic;
signal \N__45773\ : std_logic;
signal \N__45768\ : std_logic;
signal \N__45765\ : std_logic;
signal \N__45764\ : std_logic;
signal \N__45763\ : std_logic;
signal \N__45760\ : std_logic;
signal \N__45755\ : std_logic;
signal \N__45752\ : std_logic;
signal \N__45749\ : std_logic;
signal \N__45744\ : std_logic;
signal \N__45743\ : std_logic;
signal \N__45742\ : std_logic;
signal \N__45739\ : std_logic;
signal \N__45736\ : std_logic;
signal \N__45733\ : std_logic;
signal \N__45730\ : std_logic;
signal \N__45727\ : std_logic;
signal \N__45724\ : std_logic;
signal \N__45719\ : std_logic;
signal \N__45714\ : std_logic;
signal \N__45711\ : std_logic;
signal \N__45708\ : std_logic;
signal \N__45705\ : std_logic;
signal \N__45702\ : std_logic;
signal \N__45699\ : std_logic;
signal \N__45696\ : std_logic;
signal \N__45693\ : std_logic;
signal \N__45692\ : std_logic;
signal \N__45691\ : std_logic;
signal \N__45688\ : std_logic;
signal \N__45683\ : std_logic;
signal \N__45678\ : std_logic;
signal \N__45675\ : std_logic;
signal \N__45674\ : std_logic;
signal \N__45671\ : std_logic;
signal \N__45670\ : std_logic;
signal \N__45667\ : std_logic;
signal \N__45664\ : std_logic;
signal \N__45661\ : std_logic;
signal \N__45658\ : std_logic;
signal \N__45651\ : std_logic;
signal \N__45648\ : std_logic;
signal \N__45645\ : std_logic;
signal \N__45642\ : std_logic;
signal \N__45639\ : std_logic;
signal \N__45636\ : std_logic;
signal \N__45633\ : std_logic;
signal \N__45630\ : std_logic;
signal \N__45627\ : std_logic;
signal \N__45624\ : std_logic;
signal \N__45621\ : std_logic;
signal \N__45618\ : std_logic;
signal \N__45617\ : std_logic;
signal \N__45614\ : std_logic;
signal \N__45613\ : std_logic;
signal \N__45610\ : std_logic;
signal \N__45605\ : std_logic;
signal \N__45602\ : std_logic;
signal \N__45599\ : std_logic;
signal \N__45594\ : std_logic;
signal \N__45591\ : std_logic;
signal \N__45588\ : std_logic;
signal \N__45585\ : std_logic;
signal \N__45582\ : std_logic;
signal \N__45579\ : std_logic;
signal \N__45576\ : std_logic;
signal \N__45573\ : std_logic;
signal \N__45572\ : std_logic;
signal \N__45571\ : std_logic;
signal \N__45570\ : std_logic;
signal \N__45569\ : std_logic;
signal \N__45568\ : std_logic;
signal \N__45567\ : std_logic;
signal \N__45552\ : std_logic;
signal \N__45549\ : std_logic;
signal \N__45546\ : std_logic;
signal \N__45543\ : std_logic;
signal \N__45540\ : std_logic;
signal \N__45537\ : std_logic;
signal \N__45534\ : std_logic;
signal \N__45531\ : std_logic;
signal \N__45530\ : std_logic;
signal \N__45529\ : std_logic;
signal \N__45526\ : std_logic;
signal \N__45523\ : std_logic;
signal \N__45520\ : std_logic;
signal \N__45513\ : std_logic;
signal \N__45510\ : std_logic;
signal \N__45507\ : std_logic;
signal \N__45504\ : std_logic;
signal \N__45501\ : std_logic;
signal \N__45498\ : std_logic;
signal \N__45495\ : std_logic;
signal \N__45492\ : std_logic;
signal \N__45489\ : std_logic;
signal \N__45486\ : std_logic;
signal \N__45485\ : std_logic;
signal \N__45482\ : std_logic;
signal \N__45479\ : std_logic;
signal \N__45476\ : std_logic;
signal \N__45473\ : std_logic;
signal \N__45470\ : std_logic;
signal \N__45469\ : std_logic;
signal \N__45466\ : std_logic;
signal \N__45465\ : std_logic;
signal \N__45464\ : std_logic;
signal \N__45463\ : std_logic;
signal \N__45462\ : std_logic;
signal \N__45461\ : std_logic;
signal \N__45460\ : std_logic;
signal \N__45459\ : std_logic;
signal \N__45458\ : std_logic;
signal \N__45457\ : std_logic;
signal \N__45456\ : std_logic;
signal \N__45455\ : std_logic;
signal \N__45454\ : std_logic;
signal \N__45453\ : std_logic;
signal \N__45452\ : std_logic;
signal \N__45451\ : std_logic;
signal \N__45450\ : std_logic;
signal \N__45449\ : std_logic;
signal \N__45448\ : std_logic;
signal \N__45447\ : std_logic;
signal \N__45446\ : std_logic;
signal \N__45445\ : std_logic;
signal \N__45444\ : std_logic;
signal \N__45443\ : std_logic;
signal \N__45442\ : std_logic;
signal \N__45441\ : std_logic;
signal \N__45438\ : std_logic;
signal \N__45435\ : std_logic;
signal \N__45432\ : std_logic;
signal \N__45429\ : std_logic;
signal \N__45428\ : std_logic;
signal \N__45427\ : std_logic;
signal \N__45426\ : std_logic;
signal \N__45423\ : std_logic;
signal \N__45422\ : std_logic;
signal \N__45419\ : std_logic;
signal \N__45418\ : std_logic;
signal \N__45417\ : std_logic;
signal \N__45416\ : std_logic;
signal \N__45415\ : std_logic;
signal \N__45412\ : std_logic;
signal \N__45411\ : std_logic;
signal \N__45410\ : std_logic;
signal \N__45409\ : std_logic;
signal \N__45408\ : std_logic;
signal \N__45407\ : std_logic;
signal \N__45406\ : std_logic;
signal \N__45405\ : std_logic;
signal \N__45404\ : std_logic;
signal \N__45403\ : std_logic;
signal \N__45402\ : std_logic;
signal \N__45397\ : std_logic;
signal \N__45392\ : std_logic;
signal \N__45391\ : std_logic;
signal \N__45390\ : std_logic;
signal \N__45389\ : std_logic;
signal \N__45388\ : std_logic;
signal \N__45385\ : std_logic;
signal \N__45382\ : std_logic;
signal \N__45373\ : std_logic;
signal \N__45364\ : std_logic;
signal \N__45361\ : std_logic;
signal \N__45360\ : std_logic;
signal \N__45359\ : std_logic;
signal \N__45358\ : std_logic;
signal \N__45357\ : std_logic;
signal \N__45354\ : std_logic;
signal \N__45349\ : std_logic;
signal \N__45346\ : std_logic;
signal \N__45341\ : std_logic;
signal \N__45336\ : std_logic;
signal \N__45333\ : std_logic;
signal \N__45326\ : std_logic;
signal \N__45319\ : std_logic;
signal \N__45310\ : std_logic;
signal \N__45303\ : std_logic;
signal \N__45294\ : std_logic;
signal \N__45285\ : std_logic;
signal \N__45282\ : std_logic;
signal \N__45277\ : std_logic;
signal \N__45274\ : std_logic;
signal \N__45271\ : std_logic;
signal \N__45266\ : std_logic;
signal \N__45263\ : std_logic;
signal \N__45254\ : std_logic;
signal \N__45251\ : std_logic;
signal \N__45248\ : std_logic;
signal \N__45247\ : std_logic;
signal \N__45246\ : std_logic;
signal \N__45245\ : std_logic;
signal \N__45244\ : std_logic;
signal \N__45243\ : std_logic;
signal \N__45242\ : std_logic;
signal \N__45241\ : std_logic;
signal \N__45240\ : std_logic;
signal \N__45239\ : std_logic;
signal \N__45236\ : std_logic;
signal \N__45233\ : std_logic;
signal \N__45232\ : std_logic;
signal \N__45229\ : std_logic;
signal \N__45222\ : std_logic;
signal \N__45205\ : std_logic;
signal \N__45202\ : std_logic;
signal \N__45201\ : std_logic;
signal \N__45194\ : std_logic;
signal \N__45191\ : std_logic;
signal \N__45182\ : std_logic;
signal \N__45179\ : std_logic;
signal \N__45178\ : std_logic;
signal \N__45177\ : std_logic;
signal \N__45176\ : std_logic;
signal \N__45175\ : std_logic;
signal \N__45174\ : std_logic;
signal \N__45169\ : std_logic;
signal \N__45162\ : std_logic;
signal \N__45155\ : std_logic;
signal \N__45148\ : std_logic;
signal \N__45139\ : std_logic;
signal \N__45136\ : std_logic;
signal \N__45127\ : std_logic;
signal \N__45120\ : std_logic;
signal \N__45117\ : std_logic;
signal \N__45114\ : std_logic;
signal \N__45101\ : std_logic;
signal \N__45090\ : std_logic;
signal \N__45089\ : std_logic;
signal \N__45088\ : std_logic;
signal \N__45087\ : std_logic;
signal \N__45086\ : std_logic;
signal \N__45085\ : std_logic;
signal \N__45084\ : std_logic;
signal \N__45083\ : std_logic;
signal \N__45082\ : std_logic;
signal \N__45081\ : std_logic;
signal \N__45080\ : std_logic;
signal \N__45079\ : std_logic;
signal \N__45078\ : std_logic;
signal \N__45077\ : std_logic;
signal \N__45076\ : std_logic;
signal \N__45075\ : std_logic;
signal \N__45074\ : std_logic;
signal \N__45073\ : std_logic;
signal \N__45072\ : std_logic;
signal \N__45071\ : std_logic;
signal \N__45070\ : std_logic;
signal \N__45069\ : std_logic;
signal \N__45068\ : std_logic;
signal \N__45067\ : std_logic;
signal \N__45066\ : std_logic;
signal \N__45065\ : std_logic;
signal \N__45064\ : std_logic;
signal \N__45061\ : std_logic;
signal \N__45060\ : std_logic;
signal \N__45059\ : std_logic;
signal \N__45058\ : std_logic;
signal \N__45057\ : std_logic;
signal \N__45054\ : std_logic;
signal \N__45053\ : std_logic;
signal \N__45052\ : std_logic;
signal \N__45051\ : std_logic;
signal \N__45050\ : std_logic;
signal \N__45049\ : std_logic;
signal \N__45048\ : std_logic;
signal \N__45047\ : std_logic;
signal \N__45046\ : std_logic;
signal \N__45045\ : std_logic;
signal \N__45044\ : std_logic;
signal \N__45043\ : std_logic;
signal \N__45042\ : std_logic;
signal \N__45041\ : std_logic;
signal \N__45040\ : std_logic;
signal \N__45039\ : std_logic;
signal \N__45036\ : std_logic;
signal \N__45035\ : std_logic;
signal \N__45034\ : std_logic;
signal \N__45033\ : std_logic;
signal \N__45032\ : std_logic;
signal \N__45031\ : std_logic;
signal \N__45030\ : std_logic;
signal \N__45029\ : std_logic;
signal \N__45028\ : std_logic;
signal \N__45027\ : std_logic;
signal \N__45026\ : std_logic;
signal \N__45023\ : std_logic;
signal \N__45020\ : std_logic;
signal \N__45013\ : std_logic;
signal \N__45010\ : std_logic;
signal \N__44999\ : std_logic;
signal \N__44992\ : std_logic;
signal \N__44983\ : std_logic;
signal \N__44974\ : std_logic;
signal \N__44971\ : std_logic;
signal \N__44968\ : std_logic;
signal \N__44965\ : std_logic;
signal \N__44964\ : std_logic;
signal \N__44961\ : std_logic;
signal \N__44956\ : std_logic;
signal \N__44953\ : std_logic;
signal \N__44950\ : std_logic;
signal \N__44949\ : std_logic;
signal \N__44948\ : std_logic;
signal \N__44943\ : std_logic;
signal \N__44936\ : std_logic;
signal \N__44931\ : std_logic;
signal \N__44930\ : std_logic;
signal \N__44929\ : std_logic;
signal \N__44926\ : std_logic;
signal \N__44923\ : std_logic;
signal \N__44914\ : std_logic;
signal \N__44909\ : std_logic;
signal \N__44906\ : std_logic;
signal \N__44903\ : std_logic;
signal \N__44902\ : std_logic;
signal \N__44901\ : std_logic;
signal \N__44900\ : std_logic;
signal \N__44899\ : std_logic;
signal \N__44898\ : std_logic;
signal \N__44897\ : std_logic;
signal \N__44896\ : std_logic;
signal \N__44895\ : std_logic;
signal \N__44894\ : std_logic;
signal \N__44889\ : std_logic;
signal \N__44882\ : std_logic;
signal \N__44873\ : std_logic;
signal \N__44870\ : std_logic;
signal \N__44853\ : std_logic;
signal \N__44850\ : std_logic;
signal \N__44847\ : std_logic;
signal \N__44844\ : std_logic;
signal \N__44835\ : std_logic;
signal \N__44832\ : std_logic;
signal \N__44829\ : std_logic;
signal \N__44822\ : std_logic;
signal \N__44817\ : std_logic;
signal \N__44804\ : std_logic;
signal \N__44801\ : std_logic;
signal \N__44796\ : std_logic;
signal \N__44793\ : std_logic;
signal \N__44788\ : std_logic;
signal \N__44781\ : std_logic;
signal \N__44776\ : std_logic;
signal \N__44771\ : std_logic;
signal \N__44766\ : std_logic;
signal \N__44763\ : std_logic;
signal \N__44758\ : std_logic;
signal \N__44751\ : std_logic;
signal \N__44746\ : std_logic;
signal \N__44721\ : std_logic;
signal \N__44718\ : std_logic;
signal \N__44715\ : std_logic;
signal \N__44712\ : std_logic;
signal \N__44709\ : std_logic;
signal \N__44706\ : std_logic;
signal \N__44703\ : std_logic;
signal \N__44700\ : std_logic;
signal \N__44697\ : std_logic;
signal \N__44694\ : std_logic;
signal \N__44691\ : std_logic;
signal \N__44688\ : std_logic;
signal \N__44685\ : std_logic;
signal \N__44682\ : std_logic;
signal \N__44679\ : std_logic;
signal \N__44676\ : std_logic;
signal \N__44675\ : std_logic;
signal \N__44672\ : std_logic;
signal \N__44669\ : std_logic;
signal \N__44666\ : std_logic;
signal \N__44665\ : std_logic;
signal \N__44664\ : std_logic;
signal \N__44663\ : std_logic;
signal \N__44662\ : std_logic;
signal \N__44661\ : std_logic;
signal \N__44660\ : std_logic;
signal \N__44659\ : std_logic;
signal \N__44658\ : std_logic;
signal \N__44657\ : std_logic;
signal \N__44654\ : std_logic;
signal \N__44651\ : std_logic;
signal \N__44648\ : std_logic;
signal \N__44647\ : std_logic;
signal \N__44644\ : std_logic;
signal \N__44641\ : std_logic;
signal \N__44640\ : std_logic;
signal \N__44639\ : std_logic;
signal \N__44636\ : std_logic;
signal \N__44635\ : std_logic;
signal \N__44632\ : std_logic;
signal \N__44629\ : std_logic;
signal \N__44628\ : std_logic;
signal \N__44625\ : std_logic;
signal \N__44624\ : std_logic;
signal \N__44621\ : std_logic;
signal \N__44618\ : std_logic;
signal \N__44617\ : std_logic;
signal \N__44616\ : std_logic;
signal \N__44615\ : std_logic;
signal \N__44614\ : std_logic;
signal \N__44609\ : std_logic;
signal \N__44606\ : std_logic;
signal \N__44603\ : std_logic;
signal \N__44598\ : std_logic;
signal \N__44593\ : std_logic;
signal \N__44592\ : std_logic;
signal \N__44591\ : std_logic;
signal \N__44590\ : std_logic;
signal \N__44585\ : std_logic;
signal \N__44582\ : std_logic;
signal \N__44577\ : std_logic;
signal \N__44572\ : std_logic;
signal \N__44567\ : std_logic;
signal \N__44564\ : std_logic;
signal \N__44557\ : std_logic;
signal \N__44552\ : std_logic;
signal \N__44549\ : std_logic;
signal \N__44548\ : std_logic;
signal \N__44547\ : std_logic;
signal \N__44542\ : std_logic;
signal \N__44541\ : std_logic;
signal \N__44538\ : std_logic;
signal \N__44535\ : std_logic;
signal \N__44534\ : std_logic;
signal \N__44533\ : std_logic;
signal \N__44530\ : std_logic;
signal \N__44527\ : std_logic;
signal \N__44518\ : std_logic;
signal \N__44515\ : std_logic;
signal \N__44510\ : std_logic;
signal \N__44509\ : std_logic;
signal \N__44508\ : std_logic;
signal \N__44505\ : std_logic;
signal \N__44500\ : std_logic;
signal \N__44497\ : std_logic;
signal \N__44486\ : std_logic;
signal \N__44479\ : std_logic;
signal \N__44474\ : std_logic;
signal \N__44469\ : std_logic;
signal \N__44454\ : std_logic;
signal \N__44451\ : std_logic;
signal \N__44448\ : std_logic;
signal \N__44445\ : std_logic;
signal \N__44442\ : std_logic;
signal \N__44439\ : std_logic;
signal \N__44436\ : std_logic;
signal \N__44433\ : std_logic;
signal \N__44432\ : std_logic;
signal \N__44431\ : std_logic;
signal \N__44428\ : std_logic;
signal \N__44427\ : std_logic;
signal \N__44422\ : std_logic;
signal \N__44419\ : std_logic;
signal \N__44418\ : std_logic;
signal \N__44415\ : std_logic;
signal \N__44414\ : std_logic;
signal \N__44413\ : std_logic;
signal \N__44410\ : std_logic;
signal \N__44409\ : std_logic;
signal \N__44408\ : std_logic;
signal \N__44407\ : std_logic;
signal \N__44406\ : std_logic;
signal \N__44403\ : std_logic;
signal \N__44400\ : std_logic;
signal \N__44397\ : std_logic;
signal \N__44394\ : std_logic;
signal \N__44391\ : std_logic;
signal \N__44388\ : std_logic;
signal \N__44383\ : std_logic;
signal \N__44378\ : std_logic;
signal \N__44373\ : std_logic;
signal \N__44372\ : std_logic;
signal \N__44371\ : std_logic;
signal \N__44370\ : std_logic;
signal \N__44369\ : std_logic;
signal \N__44368\ : std_logic;
signal \N__44367\ : std_logic;
signal \N__44360\ : std_logic;
signal \N__44355\ : std_logic;
signal \N__44350\ : std_logic;
signal \N__44343\ : std_logic;
signal \N__44340\ : std_logic;
signal \N__44335\ : std_logic;
signal \N__44334\ : std_logic;
signal \N__44333\ : std_logic;
signal \N__44332\ : std_logic;
signal \N__44331\ : std_logic;
signal \N__44330\ : std_logic;
signal \N__44329\ : std_logic;
signal \N__44328\ : std_logic;
signal \N__44327\ : std_logic;
signal \N__44326\ : std_logic;
signal \N__44323\ : std_logic;
signal \N__44320\ : std_logic;
signal \N__44315\ : std_logic;
signal \N__44310\ : std_logic;
signal \N__44305\ : std_logic;
signal \N__44300\ : std_logic;
signal \N__44289\ : std_logic;
signal \N__44274\ : std_logic;
signal \N__44271\ : std_logic;
signal \N__44268\ : std_logic;
signal \N__44265\ : std_logic;
signal \N__44262\ : std_logic;
signal \N__44259\ : std_logic;
signal \N__44256\ : std_logic;
signal \N__44253\ : std_logic;
signal \N__44250\ : std_logic;
signal \N__44247\ : std_logic;
signal \N__44244\ : std_logic;
signal \N__44241\ : std_logic;
signal \N__44238\ : std_logic;
signal \N__44235\ : std_logic;
signal \N__44232\ : std_logic;
signal \N__44229\ : std_logic;
signal \N__44226\ : std_logic;
signal \N__44223\ : std_logic;
signal \N__44220\ : std_logic;
signal \N__44217\ : std_logic;
signal \N__44214\ : std_logic;
signal \N__44211\ : std_logic;
signal \N__44208\ : std_logic;
signal \N__44205\ : std_logic;
signal \N__44202\ : std_logic;
signal \N__44199\ : std_logic;
signal \N__44196\ : std_logic;
signal \N__44193\ : std_logic;
signal \N__44190\ : std_logic;
signal \N__44187\ : std_logic;
signal \N__44184\ : std_logic;
signal \N__44181\ : std_logic;
signal \N__44178\ : std_logic;
signal \N__44175\ : std_logic;
signal \N__44172\ : std_logic;
signal \N__44169\ : std_logic;
signal \N__44166\ : std_logic;
signal \N__44163\ : std_logic;
signal \N__44160\ : std_logic;
signal \N__44157\ : std_logic;
signal \N__44154\ : std_logic;
signal \N__44151\ : std_logic;
signal \N__44148\ : std_logic;
signal \N__44145\ : std_logic;
signal \N__44142\ : std_logic;
signal \N__44141\ : std_logic;
signal \N__44140\ : std_logic;
signal \N__44135\ : std_logic;
signal \N__44132\ : std_logic;
signal \N__44127\ : std_logic;
signal \N__44124\ : std_logic;
signal \N__44121\ : std_logic;
signal \N__44118\ : std_logic;
signal \N__44115\ : std_logic;
signal \N__44112\ : std_logic;
signal \N__44109\ : std_logic;
signal \N__44106\ : std_logic;
signal \N__44105\ : std_logic;
signal \N__44102\ : std_logic;
signal \N__44099\ : std_logic;
signal \N__44096\ : std_logic;
signal \N__44093\ : std_logic;
signal \N__44092\ : std_logic;
signal \N__44089\ : std_logic;
signal \N__44088\ : std_logic;
signal \N__44085\ : std_logic;
signal \N__44082\ : std_logic;
signal \N__44079\ : std_logic;
signal \N__44076\ : std_logic;
signal \N__44071\ : std_logic;
signal \N__44068\ : std_logic;
signal \N__44065\ : std_logic;
signal \N__44062\ : std_logic;
signal \N__44061\ : std_logic;
signal \N__44058\ : std_logic;
signal \N__44055\ : std_logic;
signal \N__44052\ : std_logic;
signal \N__44049\ : std_logic;
signal \N__44046\ : std_logic;
signal \N__44043\ : std_logic;
signal \N__44040\ : std_logic;
signal \N__44035\ : std_logic;
signal \N__44030\ : std_logic;
signal \N__44025\ : std_logic;
signal \N__44022\ : std_logic;
signal \N__44019\ : std_logic;
signal \N__44016\ : std_logic;
signal \N__44013\ : std_logic;
signal \N__44010\ : std_logic;
signal \N__44007\ : std_logic;
signal \N__44004\ : std_logic;
signal \N__44003\ : std_logic;
signal \N__44000\ : std_logic;
signal \N__43997\ : std_logic;
signal \N__43994\ : std_logic;
signal \N__43991\ : std_logic;
signal \N__43988\ : std_logic;
signal \N__43985\ : std_logic;
signal \N__43982\ : std_logic;
signal \N__43979\ : std_logic;
signal \N__43974\ : std_logic;
signal \N__43971\ : std_logic;
signal \N__43968\ : std_logic;
signal \N__43965\ : std_logic;
signal \N__43962\ : std_logic;
signal \N__43959\ : std_logic;
signal \N__43956\ : std_logic;
signal \N__43955\ : std_logic;
signal \N__43954\ : std_logic;
signal \N__43951\ : std_logic;
signal \N__43948\ : std_logic;
signal \N__43945\ : std_logic;
signal \N__43942\ : std_logic;
signal \N__43939\ : std_logic;
signal \N__43938\ : std_logic;
signal \N__43933\ : std_logic;
signal \N__43932\ : std_logic;
signal \N__43931\ : std_logic;
signal \N__43928\ : std_logic;
signal \N__43925\ : std_logic;
signal \N__43922\ : std_logic;
signal \N__43917\ : std_logic;
signal \N__43914\ : std_logic;
signal \N__43905\ : std_logic;
signal \N__43904\ : std_logic;
signal \N__43903\ : std_logic;
signal \N__43902\ : std_logic;
signal \N__43901\ : std_logic;
signal \N__43898\ : std_logic;
signal \N__43891\ : std_logic;
signal \N__43888\ : std_logic;
signal \N__43887\ : std_logic;
signal \N__43886\ : std_logic;
signal \N__43885\ : std_logic;
signal \N__43882\ : std_logic;
signal \N__43879\ : std_logic;
signal \N__43874\ : std_logic;
signal \N__43869\ : std_logic;
signal \N__43866\ : std_logic;
signal \N__43857\ : std_logic;
signal \N__43854\ : std_logic;
signal \N__43853\ : std_logic;
signal \N__43852\ : std_logic;
signal \N__43849\ : std_logic;
signal \N__43844\ : std_logic;
signal \N__43841\ : std_logic;
signal \N__43836\ : std_logic;
signal \N__43833\ : std_logic;
signal \N__43830\ : std_logic;
signal \N__43829\ : std_logic;
signal \N__43828\ : std_logic;
signal \N__43825\ : std_logic;
signal \N__43822\ : std_logic;
signal \N__43819\ : std_logic;
signal \N__43814\ : std_logic;
signal \N__43813\ : std_logic;
signal \N__43810\ : std_logic;
signal \N__43807\ : std_logic;
signal \N__43804\ : std_logic;
signal \N__43799\ : std_logic;
signal \N__43794\ : std_logic;
signal \N__43791\ : std_logic;
signal \N__43790\ : std_logic;
signal \N__43789\ : std_logic;
signal \N__43786\ : std_logic;
signal \N__43781\ : std_logic;
signal \N__43778\ : std_logic;
signal \N__43773\ : std_logic;
signal \N__43770\ : std_logic;
signal \N__43767\ : std_logic;
signal \N__43764\ : std_logic;
signal \N__43761\ : std_logic;
signal \N__43758\ : std_logic;
signal \N__43755\ : std_logic;
signal \N__43752\ : std_logic;
signal \N__43749\ : std_logic;
signal \N__43748\ : std_logic;
signal \N__43747\ : std_logic;
signal \N__43746\ : std_logic;
signal \N__43743\ : std_logic;
signal \N__43740\ : std_logic;
signal \N__43739\ : std_logic;
signal \N__43734\ : std_logic;
signal \N__43733\ : std_logic;
signal \N__43728\ : std_logic;
signal \N__43725\ : std_logic;
signal \N__43722\ : std_logic;
signal \N__43721\ : std_logic;
signal \N__43720\ : std_logic;
signal \N__43717\ : std_logic;
signal \N__43712\ : std_logic;
signal \N__43709\ : std_logic;
signal \N__43704\ : std_logic;
signal \N__43701\ : std_logic;
signal \N__43698\ : std_logic;
signal \N__43695\ : std_logic;
signal \N__43686\ : std_logic;
signal \N__43683\ : std_logic;
signal \N__43680\ : std_logic;
signal \N__43677\ : std_logic;
signal \N__43674\ : std_logic;
signal \N__43671\ : std_logic;
signal \N__43670\ : std_logic;
signal \N__43669\ : std_logic;
signal \N__43666\ : std_logic;
signal \N__43665\ : std_logic;
signal \N__43664\ : std_logic;
signal \N__43659\ : std_logic;
signal \N__43656\ : std_logic;
signal \N__43651\ : std_logic;
signal \N__43648\ : std_logic;
signal \N__43645\ : std_logic;
signal \N__43638\ : std_logic;
signal \N__43635\ : std_logic;
signal \N__43632\ : std_logic;
signal \N__43629\ : std_logic;
signal \N__43626\ : std_logic;
signal \N__43623\ : std_logic;
signal \N__43620\ : std_logic;
signal \N__43619\ : std_logic;
signal \N__43616\ : std_logic;
signal \N__43613\ : std_logic;
signal \N__43612\ : std_logic;
signal \N__43609\ : std_logic;
signal \N__43606\ : std_logic;
signal \N__43603\ : std_logic;
signal \N__43600\ : std_logic;
signal \N__43597\ : std_logic;
signal \N__43594\ : std_logic;
signal \N__43587\ : std_logic;
signal \N__43584\ : std_logic;
signal \N__43583\ : std_logic;
signal \N__43582\ : std_logic;
signal \N__43581\ : std_logic;
signal \N__43580\ : std_logic;
signal \N__43579\ : std_logic;
signal \N__43578\ : std_logic;
signal \N__43577\ : std_logic;
signal \N__43576\ : std_logic;
signal \N__43575\ : std_logic;
signal \N__43574\ : std_logic;
signal \N__43573\ : std_logic;
signal \N__43572\ : std_logic;
signal \N__43571\ : std_logic;
signal \N__43570\ : std_logic;
signal \N__43569\ : std_logic;
signal \N__43566\ : std_logic;
signal \N__43563\ : std_logic;
signal \N__43562\ : std_logic;
signal \N__43561\ : std_logic;
signal \N__43560\ : std_logic;
signal \N__43559\ : std_logic;
signal \N__43556\ : std_logic;
signal \N__43553\ : std_logic;
signal \N__43550\ : std_logic;
signal \N__43549\ : std_logic;
signal \N__43546\ : std_logic;
signal \N__43545\ : std_logic;
signal \N__43542\ : std_logic;
signal \N__43541\ : std_logic;
signal \N__43540\ : std_logic;
signal \N__43537\ : std_logic;
signal \N__43534\ : std_logic;
signal \N__43533\ : std_logic;
signal \N__43530\ : std_logic;
signal \N__43529\ : std_logic;
signal \N__43526\ : std_logic;
signal \N__43523\ : std_logic;
signal \N__43520\ : std_logic;
signal \N__43519\ : std_logic;
signal \N__43518\ : std_logic;
signal \N__43515\ : std_logic;
signal \N__43514\ : std_logic;
signal \N__43513\ : std_logic;
signal \N__43512\ : std_logic;
signal \N__43511\ : std_logic;
signal \N__43508\ : std_logic;
signal \N__43505\ : std_logic;
signal \N__43502\ : std_logic;
signal \N__43499\ : std_logic;
signal \N__43496\ : std_logic;
signal \N__43493\ : std_logic;
signal \N__43492\ : std_logic;
signal \N__43491\ : std_logic;
signal \N__43488\ : std_logic;
signal \N__43487\ : std_logic;
signal \N__43484\ : std_logic;
signal \N__43481\ : std_logic;
signal \N__43478\ : std_logic;
signal \N__43463\ : std_logic;
signal \N__43460\ : std_logic;
signal \N__43455\ : std_logic;
signal \N__43452\ : std_logic;
signal \N__43437\ : std_logic;
signal \N__43436\ : std_logic;
signal \N__43435\ : std_logic;
signal \N__43432\ : std_logic;
signal \N__43431\ : std_logic;
signal \N__43428\ : std_logic;
signal \N__43423\ : std_logic;
signal \N__43420\ : std_logic;
signal \N__43417\ : std_logic;
signal \N__43412\ : std_logic;
signal \N__43397\ : std_logic;
signal \N__43392\ : std_logic;
signal \N__43389\ : std_logic;
signal \N__43384\ : std_logic;
signal \N__43381\ : std_logic;
signal \N__43378\ : std_logic;
signal \N__43371\ : std_logic;
signal \N__43370\ : std_logic;
signal \N__43367\ : std_logic;
signal \N__43366\ : std_logic;
signal \N__43365\ : std_logic;
signal \N__43362\ : std_logic;
signal \N__43359\ : std_logic;
signal \N__43356\ : std_logic;
signal \N__43351\ : std_logic;
signal \N__43342\ : std_logic;
signal \N__43335\ : std_logic;
signal \N__43330\ : std_logic;
signal \N__43325\ : std_logic;
signal \N__43322\ : std_logic;
signal \N__43315\ : std_logic;
signal \N__43310\ : std_logic;
signal \N__43299\ : std_logic;
signal \N__43296\ : std_logic;
signal \N__43293\ : std_logic;
signal \N__43290\ : std_logic;
signal \N__43287\ : std_logic;
signal \N__43284\ : std_logic;
signal \N__43281\ : std_logic;
signal \N__43278\ : std_logic;
signal \N__43275\ : std_logic;
signal \N__43272\ : std_logic;
signal \N__43269\ : std_logic;
signal \N__43268\ : std_logic;
signal \N__43265\ : std_logic;
signal \N__43262\ : std_logic;
signal \N__43257\ : std_logic;
signal \N__43254\ : std_logic;
signal \N__43251\ : std_logic;
signal \N__43248\ : std_logic;
signal \N__43245\ : std_logic;
signal \N__43242\ : std_logic;
signal \N__43239\ : std_logic;
signal \N__43236\ : std_logic;
signal \N__43235\ : std_logic;
signal \N__43232\ : std_logic;
signal \N__43229\ : std_logic;
signal \N__43224\ : std_logic;
signal \N__43221\ : std_logic;
signal \N__43218\ : std_logic;
signal \N__43215\ : std_logic;
signal \N__43212\ : std_logic;
signal \N__43209\ : std_logic;
signal \N__43206\ : std_logic;
signal \N__43205\ : std_logic;
signal \N__43202\ : std_logic;
signal \N__43199\ : std_logic;
signal \N__43196\ : std_logic;
signal \N__43193\ : std_logic;
signal \N__43188\ : std_logic;
signal \N__43185\ : std_logic;
signal \N__43182\ : std_logic;
signal \N__43179\ : std_logic;
signal \N__43176\ : std_logic;
signal \N__43173\ : std_logic;
signal \N__43170\ : std_logic;
signal \N__43167\ : std_logic;
signal \N__43164\ : std_logic;
signal \N__43161\ : std_logic;
signal \N__43158\ : std_logic;
signal \N__43155\ : std_logic;
signal \N__43152\ : std_logic;
signal \N__43149\ : std_logic;
signal \N__43146\ : std_logic;
signal \N__43143\ : std_logic;
signal \N__43142\ : std_logic;
signal \N__43139\ : std_logic;
signal \N__43136\ : std_logic;
signal \N__43135\ : std_logic;
signal \N__43134\ : std_logic;
signal \N__43131\ : std_logic;
signal \N__43124\ : std_logic;
signal \N__43119\ : std_logic;
signal \N__43116\ : std_logic;
signal \N__43113\ : std_logic;
signal \N__43110\ : std_logic;
signal \N__43107\ : std_logic;
signal \N__43104\ : std_logic;
signal \N__43101\ : std_logic;
signal \N__43098\ : std_logic;
signal \N__43095\ : std_logic;
signal \N__43092\ : std_logic;
signal \N__43089\ : std_logic;
signal \N__43086\ : std_logic;
signal \N__43083\ : std_logic;
signal \N__43080\ : std_logic;
signal \N__43077\ : std_logic;
signal \N__43074\ : std_logic;
signal \N__43071\ : std_logic;
signal \N__43068\ : std_logic;
signal \N__43065\ : std_logic;
signal \N__43062\ : std_logic;
signal \N__43059\ : std_logic;
signal \N__43056\ : std_logic;
signal \N__43053\ : std_logic;
signal \N__43050\ : std_logic;
signal \N__43047\ : std_logic;
signal \N__43044\ : std_logic;
signal \N__43041\ : std_logic;
signal \N__43038\ : std_logic;
signal \N__43035\ : std_logic;
signal \N__43034\ : std_logic;
signal \N__43031\ : std_logic;
signal \N__43028\ : std_logic;
signal \N__43023\ : std_logic;
signal \N__43020\ : std_logic;
signal \N__43017\ : std_logic;
signal \N__43014\ : std_logic;
signal \N__43011\ : std_logic;
signal \N__43008\ : std_logic;
signal \N__43005\ : std_logic;
signal \N__43004\ : std_logic;
signal \N__43003\ : std_logic;
signal \N__43000\ : std_logic;
signal \N__42997\ : std_logic;
signal \N__42994\ : std_logic;
signal \N__42991\ : std_logic;
signal \N__42986\ : std_logic;
signal \N__42983\ : std_logic;
signal \N__42980\ : std_logic;
signal \N__42975\ : std_logic;
signal \N__42972\ : std_logic;
signal \N__42969\ : std_logic;
signal \N__42966\ : std_logic;
signal \N__42965\ : std_logic;
signal \N__42964\ : std_logic;
signal \N__42961\ : std_logic;
signal \N__42956\ : std_logic;
signal \N__42951\ : std_logic;
signal \N__42948\ : std_logic;
signal \N__42945\ : std_logic;
signal \N__42944\ : std_logic;
signal \N__42941\ : std_logic;
signal \N__42940\ : std_logic;
signal \N__42937\ : std_logic;
signal \N__42934\ : std_logic;
signal \N__42931\ : std_logic;
signal \N__42928\ : std_logic;
signal \N__42921\ : std_logic;
signal \N__42918\ : std_logic;
signal \N__42915\ : std_logic;
signal \N__42912\ : std_logic;
signal \N__42909\ : std_logic;
signal \N__42906\ : std_logic;
signal \N__42905\ : std_logic;
signal \N__42904\ : std_logic;
signal \N__42901\ : std_logic;
signal \N__42898\ : std_logic;
signal \N__42895\ : std_logic;
signal \N__42888\ : std_logic;
signal \N__42885\ : std_logic;
signal \N__42882\ : std_logic;
signal \N__42879\ : std_logic;
signal \N__42876\ : std_logic;
signal \N__42873\ : std_logic;
signal \N__42870\ : std_logic;
signal \N__42867\ : std_logic;
signal \N__42864\ : std_logic;
signal \N__42861\ : std_logic;
signal \N__42858\ : std_logic;
signal \N__42855\ : std_logic;
signal \N__42852\ : std_logic;
signal \N__42849\ : std_logic;
signal \N__42846\ : std_logic;
signal \N__42843\ : std_logic;
signal \N__42840\ : std_logic;
signal \N__42837\ : std_logic;
signal \N__42834\ : std_logic;
signal \N__42831\ : std_logic;
signal \N__42828\ : std_logic;
signal \N__42825\ : std_logic;
signal \N__42822\ : std_logic;
signal \N__42819\ : std_logic;
signal \N__42816\ : std_logic;
signal \N__42813\ : std_logic;
signal \N__42812\ : std_logic;
signal \N__42809\ : std_logic;
signal \N__42806\ : std_logic;
signal \N__42803\ : std_logic;
signal \N__42800\ : std_logic;
signal \N__42797\ : std_logic;
signal \N__42794\ : std_logic;
signal \N__42793\ : std_logic;
signal \N__42790\ : std_logic;
signal \N__42787\ : std_logic;
signal \N__42784\ : std_logic;
signal \N__42777\ : std_logic;
signal \N__42774\ : std_logic;
signal \N__42771\ : std_logic;
signal \N__42768\ : std_logic;
signal \N__42765\ : std_logic;
signal \N__42762\ : std_logic;
signal \N__42759\ : std_logic;
signal \N__42758\ : std_logic;
signal \N__42755\ : std_logic;
signal \N__42752\ : std_logic;
signal \N__42751\ : std_logic;
signal \N__42748\ : std_logic;
signal \N__42743\ : std_logic;
signal \N__42738\ : std_logic;
signal \N__42735\ : std_logic;
signal \N__42732\ : std_logic;
signal \N__42729\ : std_logic;
signal \N__42728\ : std_logic;
signal \N__42725\ : std_logic;
signal \N__42724\ : std_logic;
signal \N__42721\ : std_logic;
signal \N__42718\ : std_logic;
signal \N__42715\ : std_logic;
signal \N__42712\ : std_logic;
signal \N__42705\ : std_logic;
signal \N__42702\ : std_logic;
signal \N__42701\ : std_logic;
signal \N__42698\ : std_logic;
signal \N__42697\ : std_logic;
signal \N__42694\ : std_logic;
signal \N__42691\ : std_logic;
signal \N__42686\ : std_logic;
signal \N__42681\ : std_logic;
signal \N__42678\ : std_logic;
signal \N__42675\ : std_logic;
signal \N__42674\ : std_logic;
signal \N__42671\ : std_logic;
signal \N__42670\ : std_logic;
signal \N__42667\ : std_logic;
signal \N__42664\ : std_logic;
signal \N__42661\ : std_logic;
signal \N__42658\ : std_logic;
signal \N__42655\ : std_logic;
signal \N__42650\ : std_logic;
signal \N__42645\ : std_logic;
signal \N__42644\ : std_logic;
signal \N__42643\ : std_logic;
signal \N__42640\ : std_logic;
signal \N__42637\ : std_logic;
signal \N__42634\ : std_logic;
signal \N__42629\ : std_logic;
signal \N__42626\ : std_logic;
signal \N__42623\ : std_logic;
signal \N__42620\ : std_logic;
signal \N__42617\ : std_logic;
signal \N__42612\ : std_logic;
signal \N__42609\ : std_logic;
signal \N__42608\ : std_logic;
signal \N__42605\ : std_logic;
signal \N__42604\ : std_logic;
signal \N__42601\ : std_logic;
signal \N__42598\ : std_logic;
signal \N__42593\ : std_logic;
signal \N__42590\ : std_logic;
signal \N__42587\ : std_logic;
signal \N__42582\ : std_logic;
signal \N__42579\ : std_logic;
signal \N__42578\ : std_logic;
signal \N__42577\ : std_logic;
signal \N__42574\ : std_logic;
signal \N__42569\ : std_logic;
signal \N__42566\ : std_logic;
signal \N__42563\ : std_logic;
signal \N__42558\ : std_logic;
signal \N__42555\ : std_logic;
signal \N__42554\ : std_logic;
signal \N__42551\ : std_logic;
signal \N__42550\ : std_logic;
signal \N__42547\ : std_logic;
signal \N__42544\ : std_logic;
signal \N__42541\ : std_logic;
signal \N__42538\ : std_logic;
signal \N__42531\ : std_logic;
signal \N__42528\ : std_logic;
signal \N__42527\ : std_logic;
signal \N__42524\ : std_logic;
signal \N__42521\ : std_logic;
signal \N__42518\ : std_logic;
signal \N__42515\ : std_logic;
signal \N__42514\ : std_logic;
signal \N__42511\ : std_logic;
signal \N__42508\ : std_logic;
signal \N__42505\ : std_logic;
signal \N__42502\ : std_logic;
signal \N__42497\ : std_logic;
signal \N__42494\ : std_logic;
signal \N__42489\ : std_logic;
signal \N__42486\ : std_logic;
signal \N__42483\ : std_logic;
signal \N__42482\ : std_logic;
signal \N__42481\ : std_logic;
signal \N__42478\ : std_logic;
signal \N__42475\ : std_logic;
signal \N__42472\ : std_logic;
signal \N__42467\ : std_logic;
signal \N__42464\ : std_logic;
signal \N__42461\ : std_logic;
signal \N__42458\ : std_logic;
signal \N__42455\ : std_logic;
signal \N__42452\ : std_logic;
signal \N__42447\ : std_logic;
signal \N__42446\ : std_logic;
signal \N__42445\ : std_logic;
signal \N__42440\ : std_logic;
signal \N__42437\ : std_logic;
signal \N__42434\ : std_logic;
signal \N__42431\ : std_logic;
signal \N__42428\ : std_logic;
signal \N__42423\ : std_logic;
signal \N__42420\ : std_logic;
signal \N__42419\ : std_logic;
signal \N__42416\ : std_logic;
signal \N__42413\ : std_logic;
signal \N__42412\ : std_logic;
signal \N__42409\ : std_logic;
signal \N__42404\ : std_logic;
signal \N__42399\ : std_logic;
signal \N__42396\ : std_logic;
signal \N__42393\ : std_logic;
signal \N__42390\ : std_logic;
signal \N__42387\ : std_logic;
signal \N__42384\ : std_logic;
signal \N__42381\ : std_logic;
signal \N__42378\ : std_logic;
signal \N__42375\ : std_logic;
signal \N__42372\ : std_logic;
signal \N__42369\ : std_logic;
signal \N__42366\ : std_logic;
signal \N__42363\ : std_logic;
signal \N__42360\ : std_logic;
signal \N__42357\ : std_logic;
signal \N__42354\ : std_logic;
signal \N__42351\ : std_logic;
signal \N__42348\ : std_logic;
signal \N__42345\ : std_logic;
signal \N__42342\ : std_logic;
signal \N__42339\ : std_logic;
signal \N__42336\ : std_logic;
signal \N__42333\ : std_logic;
signal \N__42330\ : std_logic;
signal \N__42327\ : std_logic;
signal \N__42324\ : std_logic;
signal \N__42321\ : std_logic;
signal \N__42318\ : std_logic;
signal \N__42315\ : std_logic;
signal \N__42312\ : std_logic;
signal \N__42309\ : std_logic;
signal \N__42306\ : std_logic;
signal \N__42303\ : std_logic;
signal \N__42300\ : std_logic;
signal \N__42297\ : std_logic;
signal \N__42294\ : std_logic;
signal \N__42291\ : std_logic;
signal \N__42288\ : std_logic;
signal \N__42285\ : std_logic;
signal \N__42282\ : std_logic;
signal \N__42279\ : std_logic;
signal \N__42278\ : std_logic;
signal \N__42277\ : std_logic;
signal \N__42274\ : std_logic;
signal \N__42269\ : std_logic;
signal \N__42266\ : std_logic;
signal \N__42263\ : std_logic;
signal \N__42260\ : std_logic;
signal \N__42257\ : std_logic;
signal \N__42252\ : std_logic;
signal \N__42249\ : std_logic;
signal \N__42248\ : std_logic;
signal \N__42247\ : std_logic;
signal \N__42244\ : std_logic;
signal \N__42239\ : std_logic;
signal \N__42236\ : std_logic;
signal \N__42233\ : std_logic;
signal \N__42230\ : std_logic;
signal \N__42227\ : std_logic;
signal \N__42224\ : std_logic;
signal \N__42221\ : std_logic;
signal \N__42216\ : std_logic;
signal \N__42213\ : std_logic;
signal \N__42212\ : std_logic;
signal \N__42209\ : std_logic;
signal \N__42208\ : std_logic;
signal \N__42205\ : std_logic;
signal \N__42202\ : std_logic;
signal \N__42199\ : std_logic;
signal \N__42196\ : std_logic;
signal \N__42191\ : std_logic;
signal \N__42188\ : std_logic;
signal \N__42185\ : std_logic;
signal \N__42182\ : std_logic;
signal \N__42177\ : std_logic;
signal \N__42176\ : std_logic;
signal \N__42175\ : std_logic;
signal \N__42172\ : std_logic;
signal \N__42169\ : std_logic;
signal \N__42166\ : std_logic;
signal \N__42163\ : std_logic;
signal \N__42160\ : std_logic;
signal \N__42153\ : std_logic;
signal \N__42150\ : std_logic;
signal \N__42147\ : std_logic;
signal \N__42144\ : std_logic;
signal \N__42141\ : std_logic;
signal \N__42138\ : std_logic;
signal \N__42135\ : std_logic;
signal \N__42132\ : std_logic;
signal \N__42129\ : std_logic;
signal \N__42126\ : std_logic;
signal \N__42123\ : std_logic;
signal \N__42120\ : std_logic;
signal \N__42117\ : std_logic;
signal \N__42114\ : std_logic;
signal \N__42111\ : std_logic;
signal \N__42108\ : std_logic;
signal \N__42105\ : std_logic;
signal \N__42102\ : std_logic;
signal \N__42099\ : std_logic;
signal \N__42096\ : std_logic;
signal \N__42093\ : std_logic;
signal \N__42090\ : std_logic;
signal \N__42087\ : std_logic;
signal \N__42084\ : std_logic;
signal \N__42081\ : std_logic;
signal \N__42078\ : std_logic;
signal \N__42075\ : std_logic;
signal \N__42072\ : std_logic;
signal \N__42069\ : std_logic;
signal \N__42066\ : std_logic;
signal \N__42063\ : std_logic;
signal \N__42060\ : std_logic;
signal \N__42057\ : std_logic;
signal \N__42054\ : std_logic;
signal \N__42051\ : std_logic;
signal \N__42048\ : std_logic;
signal \N__42045\ : std_logic;
signal \N__42042\ : std_logic;
signal \N__42039\ : std_logic;
signal \N__42036\ : std_logic;
signal \N__42033\ : std_logic;
signal \N__42030\ : std_logic;
signal \N__42027\ : std_logic;
signal \N__42024\ : std_logic;
signal \N__42021\ : std_logic;
signal \N__42018\ : std_logic;
signal \N__42015\ : std_logic;
signal \N__42012\ : std_logic;
signal \N__42011\ : std_logic;
signal \N__42010\ : std_logic;
signal \N__42007\ : std_logic;
signal \N__42004\ : std_logic;
signal \N__42001\ : std_logic;
signal \N__41998\ : std_logic;
signal \N__41993\ : std_logic;
signal \N__41988\ : std_logic;
signal \N__41985\ : std_logic;
signal \N__41982\ : std_logic;
signal \N__41979\ : std_logic;
signal \N__41976\ : std_logic;
signal \N__41973\ : std_logic;
signal \N__41970\ : std_logic;
signal \N__41967\ : std_logic;
signal \N__41964\ : std_logic;
signal \N__41961\ : std_logic;
signal \N__41958\ : std_logic;
signal \N__41955\ : std_logic;
signal \N__41952\ : std_logic;
signal \N__41949\ : std_logic;
signal \N__41946\ : std_logic;
signal \N__41943\ : std_logic;
signal \N__41940\ : std_logic;
signal \N__41937\ : std_logic;
signal \N__41934\ : std_logic;
signal \N__41931\ : std_logic;
signal \N__41928\ : std_logic;
signal \N__41925\ : std_logic;
signal \N__41922\ : std_logic;
signal \N__41919\ : std_logic;
signal \N__41916\ : std_logic;
signal \N__41913\ : std_logic;
signal \N__41910\ : std_logic;
signal \N__41907\ : std_logic;
signal \N__41904\ : std_logic;
signal \N__41901\ : std_logic;
signal \N__41898\ : std_logic;
signal \N__41895\ : std_logic;
signal \N__41892\ : std_logic;
signal \N__41889\ : std_logic;
signal \N__41886\ : std_logic;
signal \N__41883\ : std_logic;
signal \N__41880\ : std_logic;
signal \N__41877\ : std_logic;
signal \N__41874\ : std_logic;
signal \N__41871\ : std_logic;
signal \N__41868\ : std_logic;
signal \N__41865\ : std_logic;
signal \N__41862\ : std_logic;
signal \N__41859\ : std_logic;
signal \N__41856\ : std_logic;
signal \N__41853\ : std_logic;
signal \N__41850\ : std_logic;
signal \N__41847\ : std_logic;
signal \N__41844\ : std_logic;
signal \N__41841\ : std_logic;
signal \N__41838\ : std_logic;
signal \N__41835\ : std_logic;
signal \N__41832\ : std_logic;
signal \N__41829\ : std_logic;
signal \N__41826\ : std_logic;
signal \N__41823\ : std_logic;
signal \N__41820\ : std_logic;
signal \N__41817\ : std_logic;
signal \N__41814\ : std_logic;
signal \N__41811\ : std_logic;
signal \N__41808\ : std_logic;
signal \N__41807\ : std_logic;
signal \N__41806\ : std_logic;
signal \N__41803\ : std_logic;
signal \N__41800\ : std_logic;
signal \N__41797\ : std_logic;
signal \N__41796\ : std_logic;
signal \N__41791\ : std_logic;
signal \N__41788\ : std_logic;
signal \N__41787\ : std_logic;
signal \N__41786\ : std_logic;
signal \N__41783\ : std_logic;
signal \N__41778\ : std_logic;
signal \N__41773\ : std_logic;
signal \N__41766\ : std_logic;
signal \N__41763\ : std_logic;
signal \N__41760\ : std_logic;
signal \N__41757\ : std_logic;
signal \N__41754\ : std_logic;
signal \N__41753\ : std_logic;
signal \N__41752\ : std_logic;
signal \N__41749\ : std_logic;
signal \N__41746\ : std_logic;
signal \N__41743\ : std_logic;
signal \N__41740\ : std_logic;
signal \N__41735\ : std_logic;
signal \N__41734\ : std_logic;
signal \N__41733\ : std_logic;
signal \N__41730\ : std_logic;
signal \N__41729\ : std_logic;
signal \N__41726\ : std_logic;
signal \N__41723\ : std_logic;
signal \N__41720\ : std_logic;
signal \N__41717\ : std_logic;
signal \N__41714\ : std_logic;
signal \N__41703\ : std_logic;
signal \N__41700\ : std_logic;
signal \N__41697\ : std_logic;
signal \N__41694\ : std_logic;
signal \N__41691\ : std_logic;
signal \N__41690\ : std_logic;
signal \N__41689\ : std_logic;
signal \N__41688\ : std_logic;
signal \N__41685\ : std_logic;
signal \N__41682\ : std_logic;
signal \N__41679\ : std_logic;
signal \N__41676\ : std_logic;
signal \N__41671\ : std_logic;
signal \N__41668\ : std_logic;
signal \N__41665\ : std_logic;
signal \N__41662\ : std_logic;
signal \N__41659\ : std_logic;
signal \N__41658\ : std_logic;
signal \N__41655\ : std_logic;
signal \N__41652\ : std_logic;
signal \N__41649\ : std_logic;
signal \N__41646\ : std_logic;
signal \N__41643\ : std_logic;
signal \N__41638\ : std_logic;
signal \N__41635\ : std_logic;
signal \N__41628\ : std_logic;
signal \N__41625\ : std_logic;
signal \N__41622\ : std_logic;
signal \N__41619\ : std_logic;
signal \N__41616\ : std_logic;
signal \N__41613\ : std_logic;
signal \N__41610\ : std_logic;
signal \N__41609\ : std_logic;
signal \N__41606\ : std_logic;
signal \N__41603\ : std_logic;
signal \N__41598\ : std_logic;
signal \N__41595\ : std_logic;
signal \N__41592\ : std_logic;
signal \N__41589\ : std_logic;
signal \N__41586\ : std_logic;
signal \N__41583\ : std_logic;
signal \N__41580\ : std_logic;
signal \N__41577\ : std_logic;
signal \N__41576\ : std_logic;
signal \N__41575\ : std_logic;
signal \N__41574\ : std_logic;
signal \N__41571\ : std_logic;
signal \N__41564\ : std_logic;
signal \N__41563\ : std_logic;
signal \N__41560\ : std_logic;
signal \N__41557\ : std_logic;
signal \N__41554\ : std_logic;
signal \N__41551\ : std_logic;
signal \N__41548\ : std_logic;
signal \N__41541\ : std_logic;
signal \N__41538\ : std_logic;
signal \N__41535\ : std_logic;
signal \N__41532\ : std_logic;
signal \N__41529\ : std_logic;
signal \N__41526\ : std_logic;
signal \N__41523\ : std_logic;
signal \N__41522\ : std_logic;
signal \N__41521\ : std_logic;
signal \N__41518\ : std_logic;
signal \N__41517\ : std_logic;
signal \N__41512\ : std_logic;
signal \N__41509\ : std_logic;
signal \N__41506\ : std_logic;
signal \N__41503\ : std_logic;
signal \N__41500\ : std_logic;
signal \N__41497\ : std_logic;
signal \N__41494\ : std_logic;
signal \N__41487\ : std_logic;
signal \N__41484\ : std_logic;
signal \N__41481\ : std_logic;
signal \N__41478\ : std_logic;
signal \N__41475\ : std_logic;
signal \N__41472\ : std_logic;
signal \N__41469\ : std_logic;
signal \N__41466\ : std_logic;
signal \N__41463\ : std_logic;
signal \N__41460\ : std_logic;
signal \N__41457\ : std_logic;
signal \N__41454\ : std_logic;
signal \N__41451\ : std_logic;
signal \N__41448\ : std_logic;
signal \N__41445\ : std_logic;
signal \N__41442\ : std_logic;
signal \N__41439\ : std_logic;
signal \N__41436\ : std_logic;
signal \N__41433\ : std_logic;
signal \N__41430\ : std_logic;
signal \N__41427\ : std_logic;
signal \N__41424\ : std_logic;
signal \N__41421\ : std_logic;
signal \N__41420\ : std_logic;
signal \N__41417\ : std_logic;
signal \N__41414\ : std_logic;
signal \N__41413\ : std_logic;
signal \N__41410\ : std_logic;
signal \N__41407\ : std_logic;
signal \N__41406\ : std_logic;
signal \N__41403\ : std_logic;
signal \N__41400\ : std_logic;
signal \N__41397\ : std_logic;
signal \N__41394\ : std_logic;
signal \N__41385\ : std_logic;
signal \N__41382\ : std_logic;
signal \N__41379\ : std_logic;
signal \N__41378\ : std_logic;
signal \N__41377\ : std_logic;
signal \N__41376\ : std_logic;
signal \N__41375\ : std_logic;
signal \N__41372\ : std_logic;
signal \N__41369\ : std_logic;
signal \N__41366\ : std_logic;
signal \N__41363\ : std_logic;
signal \N__41360\ : std_logic;
signal \N__41355\ : std_logic;
signal \N__41352\ : std_logic;
signal \N__41349\ : std_logic;
signal \N__41348\ : std_logic;
signal \N__41343\ : std_logic;
signal \N__41338\ : std_logic;
signal \N__41335\ : std_logic;
signal \N__41328\ : std_logic;
signal \N__41325\ : std_logic;
signal \N__41322\ : std_logic;
signal \N__41319\ : std_logic;
signal \N__41316\ : std_logic;
signal \N__41313\ : std_logic;
signal \N__41310\ : std_logic;
signal \N__41307\ : std_logic;
signal \N__41304\ : std_logic;
signal \N__41301\ : std_logic;
signal \N__41298\ : std_logic;
signal \N__41295\ : std_logic;
signal \N__41292\ : std_logic;
signal \N__41289\ : std_logic;
signal \N__41286\ : std_logic;
signal \N__41283\ : std_logic;
signal \N__41280\ : std_logic;
signal \N__41277\ : std_logic;
signal \N__41274\ : std_logic;
signal \N__41271\ : std_logic;
signal \N__41268\ : std_logic;
signal \N__41265\ : std_logic;
signal \N__41262\ : std_logic;
signal \N__41259\ : std_logic;
signal \N__41256\ : std_logic;
signal \N__41253\ : std_logic;
signal \N__41250\ : std_logic;
signal \N__41247\ : std_logic;
signal \N__41244\ : std_logic;
signal \N__41241\ : std_logic;
signal \N__41238\ : std_logic;
signal \N__41235\ : std_logic;
signal \N__41234\ : std_logic;
signal \N__41231\ : std_logic;
signal \N__41228\ : std_logic;
signal \N__41225\ : std_logic;
signal \N__41222\ : std_logic;
signal \N__41221\ : std_logic;
signal \N__41218\ : std_logic;
signal \N__41215\ : std_logic;
signal \N__41212\ : std_logic;
signal \N__41209\ : std_logic;
signal \N__41202\ : std_logic;
signal \N__41201\ : std_logic;
signal \N__41198\ : std_logic;
signal \N__41197\ : std_logic;
signal \N__41194\ : std_logic;
signal \N__41191\ : std_logic;
signal \N__41188\ : std_logic;
signal \N__41185\ : std_logic;
signal \N__41182\ : std_logic;
signal \N__41179\ : std_logic;
signal \N__41176\ : std_logic;
signal \N__41169\ : std_logic;
signal \N__41166\ : std_logic;
signal \N__41163\ : std_logic;
signal \N__41160\ : std_logic;
signal \N__41157\ : std_logic;
signal \N__41154\ : std_logic;
signal \N__41151\ : std_logic;
signal \N__41148\ : std_logic;
signal \N__41145\ : std_logic;
signal \N__41142\ : std_logic;
signal \N__41139\ : std_logic;
signal \N__41136\ : std_logic;
signal \N__41133\ : std_logic;
signal \N__41130\ : std_logic;
signal \N__41127\ : std_logic;
signal \N__41126\ : std_logic;
signal \N__41125\ : std_logic;
signal \N__41122\ : std_logic;
signal \N__41119\ : std_logic;
signal \N__41116\ : std_logic;
signal \N__41113\ : std_logic;
signal \N__41110\ : std_logic;
signal \N__41107\ : std_logic;
signal \N__41104\ : std_logic;
signal \N__41101\ : std_logic;
signal \N__41098\ : std_logic;
signal \N__41093\ : std_logic;
signal \N__41088\ : std_logic;
signal \N__41087\ : std_logic;
signal \N__41084\ : std_logic;
signal \N__41083\ : std_logic;
signal \N__41078\ : std_logic;
signal \N__41075\ : std_logic;
signal \N__41072\ : std_logic;
signal \N__41067\ : std_logic;
signal \N__41064\ : std_logic;
signal \N__41061\ : std_logic;
signal \N__41058\ : std_logic;
signal \N__41055\ : std_logic;
signal \N__41054\ : std_logic;
signal \N__41053\ : std_logic;
signal \N__41050\ : std_logic;
signal \N__41047\ : std_logic;
signal \N__41044\ : std_logic;
signal \N__41041\ : std_logic;
signal \N__41038\ : std_logic;
signal \N__41035\ : std_logic;
signal \N__41028\ : std_logic;
signal \N__41025\ : std_logic;
signal \N__41022\ : std_logic;
signal \N__41021\ : std_logic;
signal \N__41020\ : std_logic;
signal \N__41017\ : std_logic;
signal \N__41014\ : std_logic;
signal \N__41011\ : std_logic;
signal \N__41008\ : std_logic;
signal \N__41005\ : std_logic;
signal \N__41002\ : std_logic;
signal \N__40997\ : std_logic;
signal \N__40994\ : std_logic;
signal \N__40991\ : std_logic;
signal \N__40986\ : std_logic;
signal \N__40985\ : std_logic;
signal \N__40982\ : std_logic;
signal \N__40979\ : std_logic;
signal \N__40974\ : std_logic;
signal \N__40973\ : std_logic;
signal \N__40970\ : std_logic;
signal \N__40967\ : std_logic;
signal \N__40962\ : std_logic;
signal \N__40961\ : std_logic;
signal \N__40958\ : std_logic;
signal \N__40957\ : std_logic;
signal \N__40954\ : std_logic;
signal \N__40949\ : std_logic;
signal \N__40946\ : std_logic;
signal \N__40943\ : std_logic;
signal \N__40938\ : std_logic;
signal \N__40935\ : std_logic;
signal \N__40932\ : std_logic;
signal \N__40929\ : std_logic;
signal \N__40926\ : std_logic;
signal \N__40923\ : std_logic;
signal \N__40920\ : std_logic;
signal \N__40917\ : std_logic;
signal \N__40914\ : std_logic;
signal \N__40911\ : std_logic;
signal \N__40908\ : std_logic;
signal \N__40905\ : std_logic;
signal \N__40902\ : std_logic;
signal \N__40899\ : std_logic;
signal \N__40896\ : std_logic;
signal \N__40893\ : std_logic;
signal \N__40892\ : std_logic;
signal \N__40889\ : std_logic;
signal \N__40888\ : std_logic;
signal \N__40885\ : std_logic;
signal \N__40882\ : std_logic;
signal \N__40879\ : std_logic;
signal \N__40876\ : std_logic;
signal \N__40871\ : std_logic;
signal \N__40868\ : std_logic;
signal \N__40865\ : std_logic;
signal \N__40860\ : std_logic;
signal \N__40857\ : std_logic;
signal \N__40854\ : std_logic;
signal \N__40851\ : std_logic;
signal \N__40848\ : std_logic;
signal \N__40845\ : std_logic;
signal \N__40842\ : std_logic;
signal \N__40839\ : std_logic;
signal \N__40836\ : std_logic;
signal \N__40833\ : std_logic;
signal \N__40830\ : std_logic;
signal \N__40827\ : std_logic;
signal \N__40824\ : std_logic;
signal \N__40823\ : std_logic;
signal \N__40822\ : std_logic;
signal \N__40819\ : std_logic;
signal \N__40816\ : std_logic;
signal \N__40813\ : std_logic;
signal \N__40806\ : std_logic;
signal \N__40803\ : std_logic;
signal \N__40800\ : std_logic;
signal \N__40797\ : std_logic;
signal \N__40794\ : std_logic;
signal \N__40791\ : std_logic;
signal \N__40788\ : std_logic;
signal \N__40785\ : std_logic;
signal \N__40782\ : std_logic;
signal \N__40779\ : std_logic;
signal \N__40776\ : std_logic;
signal \N__40773\ : std_logic;
signal \N__40770\ : std_logic;
signal \N__40767\ : std_logic;
signal \N__40766\ : std_logic;
signal \N__40763\ : std_logic;
signal \N__40760\ : std_logic;
signal \N__40759\ : std_logic;
signal \N__40754\ : std_logic;
signal \N__40751\ : std_logic;
signal \N__40748\ : std_logic;
signal \N__40745\ : std_logic;
signal \N__40742\ : std_logic;
signal \N__40739\ : std_logic;
signal \N__40736\ : std_logic;
signal \N__40731\ : std_logic;
signal \N__40728\ : std_logic;
signal \N__40725\ : std_logic;
signal \N__40722\ : std_logic;
signal \N__40721\ : std_logic;
signal \N__40718\ : std_logic;
signal \N__40717\ : std_logic;
signal \N__40714\ : std_logic;
signal \N__40711\ : std_logic;
signal \N__40708\ : std_logic;
signal \N__40705\ : std_logic;
signal \N__40698\ : std_logic;
signal \N__40697\ : std_logic;
signal \N__40696\ : std_logic;
signal \N__40693\ : std_logic;
signal \N__40690\ : std_logic;
signal \N__40687\ : std_logic;
signal \N__40684\ : std_logic;
signal \N__40681\ : std_logic;
signal \N__40678\ : std_logic;
signal \N__40675\ : std_logic;
signal \N__40672\ : std_logic;
signal \N__40669\ : std_logic;
signal \N__40666\ : std_logic;
signal \N__40663\ : std_logic;
signal \N__40660\ : std_logic;
signal \N__40653\ : std_logic;
signal \N__40650\ : std_logic;
signal \N__40647\ : std_logic;
signal \N__40644\ : std_logic;
signal \N__40641\ : std_logic;
signal \N__40638\ : std_logic;
signal \N__40635\ : std_logic;
signal \N__40632\ : std_logic;
signal \N__40629\ : std_logic;
signal \N__40626\ : std_logic;
signal \N__40623\ : std_logic;
signal \N__40620\ : std_logic;
signal \N__40617\ : std_logic;
signal \N__40614\ : std_logic;
signal \N__40611\ : std_logic;
signal \N__40608\ : std_logic;
signal \N__40605\ : std_logic;
signal \N__40602\ : std_logic;
signal \N__40599\ : std_logic;
signal \N__40596\ : std_logic;
signal \N__40593\ : std_logic;
signal \N__40590\ : std_logic;
signal \N__40587\ : std_logic;
signal \N__40584\ : std_logic;
signal \N__40581\ : std_logic;
signal \N__40578\ : std_logic;
signal \N__40575\ : std_logic;
signal \N__40572\ : std_logic;
signal \N__40569\ : std_logic;
signal \N__40566\ : std_logic;
signal \N__40563\ : std_logic;
signal \N__40560\ : std_logic;
signal \N__40557\ : std_logic;
signal \N__40554\ : std_logic;
signal \N__40551\ : std_logic;
signal \N__40548\ : std_logic;
signal \N__40545\ : std_logic;
signal \N__40544\ : std_logic;
signal \N__40543\ : std_logic;
signal \N__40540\ : std_logic;
signal \N__40535\ : std_logic;
signal \N__40530\ : std_logic;
signal \N__40529\ : std_logic;
signal \N__40526\ : std_logic;
signal \N__40523\ : std_logic;
signal \N__40520\ : std_logic;
signal \N__40517\ : std_logic;
signal \N__40514\ : std_logic;
signal \N__40511\ : std_logic;
signal \N__40510\ : std_logic;
signal \N__40507\ : std_logic;
signal \N__40504\ : std_logic;
signal \N__40501\ : std_logic;
signal \N__40498\ : std_logic;
signal \N__40491\ : std_logic;
signal \N__40488\ : std_logic;
signal \N__40485\ : std_logic;
signal \N__40482\ : std_logic;
signal \N__40479\ : std_logic;
signal \N__40476\ : std_logic;
signal \N__40473\ : std_logic;
signal \N__40470\ : std_logic;
signal \N__40467\ : std_logic;
signal \N__40464\ : std_logic;
signal \N__40461\ : std_logic;
signal \N__40458\ : std_logic;
signal \N__40455\ : std_logic;
signal \N__40452\ : std_logic;
signal \N__40449\ : std_logic;
signal \N__40446\ : std_logic;
signal \N__40443\ : std_logic;
signal \N__40440\ : std_logic;
signal \N__40437\ : std_logic;
signal \N__40434\ : std_logic;
signal \N__40431\ : std_logic;
signal \N__40428\ : std_logic;
signal \N__40425\ : std_logic;
signal \N__40422\ : std_logic;
signal \N__40419\ : std_logic;
signal \N__40416\ : std_logic;
signal \N__40413\ : std_logic;
signal \N__40410\ : std_logic;
signal \N__40407\ : std_logic;
signal \N__40404\ : std_logic;
signal \N__40401\ : std_logic;
signal \N__40398\ : std_logic;
signal \N__40395\ : std_logic;
signal \N__40392\ : std_logic;
signal \N__40389\ : std_logic;
signal \N__40386\ : std_logic;
signal \N__40383\ : std_logic;
signal \N__40380\ : std_logic;
signal \N__40377\ : std_logic;
signal \N__40374\ : std_logic;
signal \N__40371\ : std_logic;
signal \N__40368\ : std_logic;
signal \N__40365\ : std_logic;
signal \N__40362\ : std_logic;
signal \N__40359\ : std_logic;
signal \N__40356\ : std_logic;
signal \N__40353\ : std_logic;
signal \N__40350\ : std_logic;
signal \N__40347\ : std_logic;
signal \N__40344\ : std_logic;
signal \N__40341\ : std_logic;
signal \N__40338\ : std_logic;
signal \N__40335\ : std_logic;
signal \N__40332\ : std_logic;
signal \N__40329\ : std_logic;
signal \N__40326\ : std_logic;
signal \N__40323\ : std_logic;
signal \N__40320\ : std_logic;
signal \N__40317\ : std_logic;
signal \N__40314\ : std_logic;
signal \N__40311\ : std_logic;
signal \N__40308\ : std_logic;
signal \N__40305\ : std_logic;
signal \N__40302\ : std_logic;
signal \N__40299\ : std_logic;
signal \N__40296\ : std_logic;
signal \N__40293\ : std_logic;
signal \N__40290\ : std_logic;
signal \N__40287\ : std_logic;
signal \N__40284\ : std_logic;
signal \N__40281\ : std_logic;
signal \N__40278\ : std_logic;
signal \N__40275\ : std_logic;
signal \N__40272\ : std_logic;
signal \N__40269\ : std_logic;
signal \N__40266\ : std_logic;
signal \N__40263\ : std_logic;
signal \N__40260\ : std_logic;
signal \N__40257\ : std_logic;
signal \N__40254\ : std_logic;
signal \N__40251\ : std_logic;
signal \N__40248\ : std_logic;
signal \N__40245\ : std_logic;
signal \N__40242\ : std_logic;
signal \N__40239\ : std_logic;
signal \N__40236\ : std_logic;
signal \N__40233\ : std_logic;
signal \N__40230\ : std_logic;
signal \N__40227\ : std_logic;
signal \N__40224\ : std_logic;
signal \N__40221\ : std_logic;
signal \N__40218\ : std_logic;
signal \N__40215\ : std_logic;
signal \N__40212\ : std_logic;
signal \N__40209\ : std_logic;
signal \N__40206\ : std_logic;
signal \N__40203\ : std_logic;
signal \N__40200\ : std_logic;
signal \N__40197\ : std_logic;
signal \N__40194\ : std_logic;
signal \N__40191\ : std_logic;
signal \N__40188\ : std_logic;
signal \N__40185\ : std_logic;
signal \N__40182\ : std_logic;
signal \N__40179\ : std_logic;
signal \N__40176\ : std_logic;
signal \N__40173\ : std_logic;
signal \N__40170\ : std_logic;
signal \N__40167\ : std_logic;
signal \N__40164\ : std_logic;
signal \N__40161\ : std_logic;
signal \N__40158\ : std_logic;
signal \N__40155\ : std_logic;
signal \N__40152\ : std_logic;
signal \N__40149\ : std_logic;
signal \N__40146\ : std_logic;
signal \N__40143\ : std_logic;
signal \N__40140\ : std_logic;
signal \N__40137\ : std_logic;
signal \N__40134\ : std_logic;
signal \N__40131\ : std_logic;
signal \N__40128\ : std_logic;
signal \N__40125\ : std_logic;
signal \N__40122\ : std_logic;
signal \N__40119\ : std_logic;
signal \N__40116\ : std_logic;
signal \N__40113\ : std_logic;
signal \N__40112\ : std_logic;
signal \N__40111\ : std_logic;
signal \N__40108\ : std_logic;
signal \N__40105\ : std_logic;
signal \N__40102\ : std_logic;
signal \N__40099\ : std_logic;
signal \N__40098\ : std_logic;
signal \N__40097\ : std_logic;
signal \N__40096\ : std_logic;
signal \N__40093\ : std_logic;
signal \N__40090\ : std_logic;
signal \N__40087\ : std_logic;
signal \N__40080\ : std_logic;
signal \N__40077\ : std_logic;
signal \N__40074\ : std_logic;
signal \N__40069\ : std_logic;
signal \N__40064\ : std_logic;
signal \N__40061\ : std_logic;
signal \N__40060\ : std_logic;
signal \N__40059\ : std_logic;
signal \N__40056\ : std_logic;
signal \N__40053\ : std_logic;
signal \N__40048\ : std_logic;
signal \N__40041\ : std_logic;
signal \N__40038\ : std_logic;
signal \N__40037\ : std_logic;
signal \N__40034\ : std_logic;
signal \N__40033\ : std_logic;
signal \N__40030\ : std_logic;
signal \N__40027\ : std_logic;
signal \N__40024\ : std_logic;
signal \N__40021\ : std_logic;
signal \N__40018\ : std_logic;
signal \N__40015\ : std_logic;
signal \N__40012\ : std_logic;
signal \N__40009\ : std_logic;
signal \N__40002\ : std_logic;
signal \N__40001\ : std_logic;
signal \N__40000\ : std_logic;
signal \N__39997\ : std_logic;
signal \N__39994\ : std_logic;
signal \N__39991\ : std_logic;
signal \N__39988\ : std_logic;
signal \N__39985\ : std_logic;
signal \N__39982\ : std_logic;
signal \N__39979\ : std_logic;
signal \N__39976\ : std_logic;
signal \N__39971\ : std_logic;
signal \N__39966\ : std_logic;
signal \N__39963\ : std_logic;
signal \N__39960\ : std_logic;
signal \N__39957\ : std_logic;
signal \N__39954\ : std_logic;
signal \N__39951\ : std_logic;
signal \N__39948\ : std_logic;
signal \N__39945\ : std_logic;
signal \N__39942\ : std_logic;
signal \N__39939\ : std_logic;
signal \N__39936\ : std_logic;
signal \N__39933\ : std_logic;
signal \N__39930\ : std_logic;
signal \N__39927\ : std_logic;
signal \N__39924\ : std_logic;
signal \N__39921\ : std_logic;
signal \N__39918\ : std_logic;
signal \N__39915\ : std_logic;
signal \N__39912\ : std_logic;
signal \N__39909\ : std_logic;
signal \N__39908\ : std_logic;
signal \N__39905\ : std_logic;
signal \N__39902\ : std_logic;
signal \N__39897\ : std_logic;
signal \N__39894\ : std_logic;
signal \N__39893\ : std_logic;
signal \N__39890\ : std_logic;
signal \N__39887\ : std_logic;
signal \N__39882\ : std_logic;
signal \N__39879\ : std_logic;
signal \N__39878\ : std_logic;
signal \N__39875\ : std_logic;
signal \N__39872\ : std_logic;
signal \N__39867\ : std_logic;
signal \N__39864\ : std_logic;
signal \N__39863\ : std_logic;
signal \N__39860\ : std_logic;
signal \N__39857\ : std_logic;
signal \N__39852\ : std_logic;
signal \N__39849\ : std_logic;
signal \N__39848\ : std_logic;
signal \N__39845\ : std_logic;
signal \N__39842\ : std_logic;
signal \N__39837\ : std_logic;
signal \N__39834\ : std_logic;
signal \N__39833\ : std_logic;
signal \N__39830\ : std_logic;
signal \N__39827\ : std_logic;
signal \N__39824\ : std_logic;
signal \N__39819\ : std_logic;
signal \N__39816\ : std_logic;
signal \N__39815\ : std_logic;
signal \N__39814\ : std_logic;
signal \N__39813\ : std_logic;
signal \N__39812\ : std_logic;
signal \N__39811\ : std_logic;
signal \N__39810\ : std_logic;
signal \N__39809\ : std_logic;
signal \N__39800\ : std_logic;
signal \N__39799\ : std_logic;
signal \N__39798\ : std_logic;
signal \N__39797\ : std_logic;
signal \N__39796\ : std_logic;
signal \N__39795\ : std_logic;
signal \N__39794\ : std_logic;
signal \N__39793\ : std_logic;
signal \N__39792\ : std_logic;
signal \N__39791\ : std_logic;
signal \N__39782\ : std_logic;
signal \N__39779\ : std_logic;
signal \N__39770\ : std_logic;
signal \N__39761\ : std_logic;
signal \N__39758\ : std_logic;
signal \N__39757\ : std_logic;
signal \N__39754\ : std_logic;
signal \N__39747\ : std_logic;
signal \N__39744\ : std_logic;
signal \N__39743\ : std_logic;
signal \N__39742\ : std_logic;
signal \N__39739\ : std_logic;
signal \N__39736\ : std_logic;
signal \N__39733\ : std_logic;
signal \N__39730\ : std_logic;
signal \N__39725\ : std_logic;
signal \N__39714\ : std_logic;
signal \N__39711\ : std_logic;
signal \N__39710\ : std_logic;
signal \N__39707\ : std_logic;
signal \N__39704\ : std_logic;
signal \N__39701\ : std_logic;
signal \N__39696\ : std_logic;
signal \N__39695\ : std_logic;
signal \N__39692\ : std_logic;
signal \N__39689\ : std_logic;
signal \N__39686\ : std_logic;
signal \N__39683\ : std_logic;
signal \N__39680\ : std_logic;
signal \N__39677\ : std_logic;
signal \N__39674\ : std_logic;
signal \N__39671\ : std_logic;
signal \N__39666\ : std_logic;
signal \N__39663\ : std_logic;
signal \N__39660\ : std_logic;
signal \N__39657\ : std_logic;
signal \N__39654\ : std_logic;
signal \N__39653\ : std_logic;
signal \N__39650\ : std_logic;
signal \N__39647\ : std_logic;
signal \N__39646\ : std_logic;
signal \N__39643\ : std_logic;
signal \N__39640\ : std_logic;
signal \N__39637\ : std_logic;
signal \N__39634\ : std_logic;
signal \N__39631\ : std_logic;
signal \N__39624\ : std_logic;
signal \N__39621\ : std_logic;
signal \N__39618\ : std_logic;
signal \N__39617\ : std_logic;
signal \N__39614\ : std_logic;
signal \N__39613\ : std_logic;
signal \N__39612\ : std_logic;
signal \N__39611\ : std_logic;
signal \N__39608\ : std_logic;
signal \N__39605\ : std_logic;
signal \N__39596\ : std_logic;
signal \N__39595\ : std_logic;
signal \N__39590\ : std_logic;
signal \N__39587\ : std_logic;
signal \N__39584\ : std_logic;
signal \N__39579\ : std_logic;
signal \N__39576\ : std_logic;
signal \N__39573\ : std_logic;
signal \N__39570\ : std_logic;
signal \N__39567\ : std_logic;
signal \N__39566\ : std_logic;
signal \N__39565\ : std_logic;
signal \N__39564\ : std_logic;
signal \N__39561\ : std_logic;
signal \N__39558\ : std_logic;
signal \N__39555\ : std_logic;
signal \N__39552\ : std_logic;
signal \N__39547\ : std_logic;
signal \N__39540\ : std_logic;
signal \N__39537\ : std_logic;
signal \N__39536\ : std_logic;
signal \N__39535\ : std_logic;
signal \N__39532\ : std_logic;
signal \N__39529\ : std_logic;
signal \N__39526\ : std_logic;
signal \N__39521\ : std_logic;
signal \N__39516\ : std_logic;
signal \N__39513\ : std_logic;
signal \N__39512\ : std_logic;
signal \N__39509\ : std_logic;
signal \N__39506\ : std_logic;
signal \N__39505\ : std_logic;
signal \N__39500\ : std_logic;
signal \N__39497\ : std_logic;
signal \N__39494\ : std_logic;
signal \N__39489\ : std_logic;
signal \N__39486\ : std_logic;
signal \N__39485\ : std_logic;
signal \N__39482\ : std_logic;
signal \N__39479\ : std_logic;
signal \N__39476\ : std_logic;
signal \N__39475\ : std_logic;
signal \N__39470\ : std_logic;
signal \N__39467\ : std_logic;
signal \N__39464\ : std_logic;
signal \N__39459\ : std_logic;
signal \N__39456\ : std_logic;
signal \N__39455\ : std_logic;
signal \N__39452\ : std_logic;
signal \N__39449\ : std_logic;
signal \N__39448\ : std_logic;
signal \N__39445\ : std_logic;
signal \N__39442\ : std_logic;
signal \N__39439\ : std_logic;
signal \N__39434\ : std_logic;
signal \N__39429\ : std_logic;
signal \N__39426\ : std_logic;
signal \N__39425\ : std_logic;
signal \N__39422\ : std_logic;
signal \N__39421\ : std_logic;
signal \N__39418\ : std_logic;
signal \N__39415\ : std_logic;
signal \N__39412\ : std_logic;
signal \N__39405\ : std_logic;
signal \N__39402\ : std_logic;
signal \N__39401\ : std_logic;
signal \N__39400\ : std_logic;
signal \N__39397\ : std_logic;
signal \N__39396\ : std_logic;
signal \N__39393\ : std_logic;
signal \N__39392\ : std_logic;
signal \N__39389\ : std_logic;
signal \N__39386\ : std_logic;
signal \N__39383\ : std_logic;
signal \N__39382\ : std_logic;
signal \N__39381\ : std_logic;
signal \N__39378\ : std_logic;
signal \N__39375\ : std_logic;
signal \N__39374\ : std_logic;
signal \N__39373\ : std_logic;
signal \N__39366\ : std_logic;
signal \N__39363\ : std_logic;
signal \N__39362\ : std_logic;
signal \N__39359\ : std_logic;
signal \N__39354\ : std_logic;
signal \N__39351\ : std_logic;
signal \N__39350\ : std_logic;
signal \N__39347\ : std_logic;
signal \N__39346\ : std_logic;
signal \N__39345\ : std_logic;
signal \N__39340\ : std_logic;
signal \N__39337\ : std_logic;
signal \N__39336\ : std_logic;
signal \N__39329\ : std_logic;
signal \N__39326\ : std_logic;
signal \N__39325\ : std_logic;
signal \N__39322\ : std_logic;
signal \N__39319\ : std_logic;
signal \N__39316\ : std_logic;
signal \N__39315\ : std_logic;
signal \N__39314\ : std_logic;
signal \N__39309\ : std_logic;
signal \N__39306\ : std_logic;
signal \N__39305\ : std_logic;
signal \N__39300\ : std_logic;
signal \N__39297\ : std_logic;
signal \N__39296\ : std_logic;
signal \N__39293\ : std_logic;
signal \N__39290\ : std_logic;
signal \N__39287\ : std_logic;
signal \N__39286\ : std_logic;
signal \N__39283\ : std_logic;
signal \N__39282\ : std_logic;
signal \N__39281\ : std_logic;
signal \N__39278\ : std_logic;
signal \N__39273\ : std_logic;
signal \N__39270\ : std_logic;
signal \N__39265\ : std_logic;
signal \N__39262\ : std_logic;
signal \N__39259\ : std_logic;
signal \N__39254\ : std_logic;
signal \N__39253\ : std_logic;
signal \N__39244\ : std_logic;
signal \N__39241\ : std_logic;
signal \N__39236\ : std_logic;
signal \N__39231\ : std_logic;
signal \N__39226\ : std_logic;
signal \N__39223\ : std_logic;
signal \N__39220\ : std_logic;
signal \N__39217\ : std_logic;
signal \N__39212\ : std_logic;
signal \N__39207\ : std_logic;
signal \N__39204\ : std_logic;
signal \N__39199\ : std_logic;
signal \N__39196\ : std_logic;
signal \N__39193\ : std_logic;
signal \N__39186\ : std_logic;
signal \N__39183\ : std_logic;
signal \N__39180\ : std_logic;
signal \N__39177\ : std_logic;
signal \N__39174\ : std_logic;
signal \N__39171\ : std_logic;
signal \N__39168\ : std_logic;
signal \N__39165\ : std_logic;
signal \N__39162\ : std_logic;
signal \N__39159\ : std_logic;
signal \N__39156\ : std_logic;
signal \N__39153\ : std_logic;
signal \N__39150\ : std_logic;
signal \N__39147\ : std_logic;
signal \N__39146\ : std_logic;
signal \N__39145\ : std_logic;
signal \N__39144\ : std_logic;
signal \N__39143\ : std_logic;
signal \N__39142\ : std_logic;
signal \N__39141\ : std_logic;
signal \N__39140\ : std_logic;
signal \N__39137\ : std_logic;
signal \N__39134\ : std_logic;
signal \N__39133\ : std_logic;
signal \N__39132\ : std_logic;
signal \N__39125\ : std_logic;
signal \N__39120\ : std_logic;
signal \N__39117\ : std_logic;
signal \N__39116\ : std_logic;
signal \N__39115\ : std_logic;
signal \N__39114\ : std_logic;
signal \N__39113\ : std_logic;
signal \N__39110\ : std_logic;
signal \N__39109\ : std_logic;
signal \N__39108\ : std_logic;
signal \N__39107\ : std_logic;
signal \N__39106\ : std_logic;
signal \N__39105\ : std_logic;
signal \N__39102\ : std_logic;
signal \N__39099\ : std_logic;
signal \N__39096\ : std_logic;
signal \N__39093\ : std_logic;
signal \N__39088\ : std_logic;
signal \N__39079\ : std_logic;
signal \N__39076\ : std_logic;
signal \N__39073\ : std_logic;
signal \N__39064\ : std_logic;
signal \N__39059\ : std_logic;
signal \N__39042\ : std_logic;
signal \N__39039\ : std_logic;
signal \N__39036\ : std_logic;
signal \N__39033\ : std_logic;
signal \N__39032\ : std_logic;
signal \N__39029\ : std_logic;
signal \N__39026\ : std_logic;
signal \N__39023\ : std_logic;
signal \N__39018\ : std_logic;
signal \N__39015\ : std_logic;
signal \N__39012\ : std_logic;
signal \N__39011\ : std_logic;
signal \N__39008\ : std_logic;
signal \N__39005\ : std_logic;
signal \N__39002\ : std_logic;
signal \N__38999\ : std_logic;
signal \N__38994\ : std_logic;
signal \N__38991\ : std_logic;
signal \N__38988\ : std_logic;
signal \N__38985\ : std_logic;
signal \N__38982\ : std_logic;
signal \N__38979\ : std_logic;
signal \N__38976\ : std_logic;
signal \N__38973\ : std_logic;
signal \N__38970\ : std_logic;
signal \N__38967\ : std_logic;
signal \N__38964\ : std_logic;
signal \N__38961\ : std_logic;
signal \N__38960\ : std_logic;
signal \N__38957\ : std_logic;
signal \N__38954\ : std_logic;
signal \N__38949\ : std_logic;
signal \N__38946\ : std_logic;
signal \N__38943\ : std_logic;
signal \N__38940\ : std_logic;
signal \N__38937\ : std_logic;
signal \N__38934\ : std_logic;
signal \N__38931\ : std_logic;
signal \N__38928\ : std_logic;
signal \N__38925\ : std_logic;
signal \N__38922\ : std_logic;
signal \N__38919\ : std_logic;
signal \N__38916\ : std_logic;
signal \N__38913\ : std_logic;
signal \N__38912\ : std_logic;
signal \N__38909\ : std_logic;
signal \N__38906\ : std_logic;
signal \N__38905\ : std_logic;
signal \N__38904\ : std_logic;
signal \N__38903\ : std_logic;
signal \N__38900\ : std_logic;
signal \N__38897\ : std_logic;
signal \N__38894\ : std_logic;
signal \N__38893\ : std_logic;
signal \N__38892\ : std_logic;
signal \N__38891\ : std_logic;
signal \N__38886\ : std_logic;
signal \N__38881\ : std_logic;
signal \N__38878\ : std_logic;
signal \N__38873\ : std_logic;
signal \N__38870\ : std_logic;
signal \N__38867\ : std_logic;
signal \N__38862\ : std_logic;
signal \N__38859\ : std_logic;
signal \N__38856\ : std_logic;
signal \N__38851\ : std_logic;
signal \N__38848\ : std_logic;
signal \N__38845\ : std_logic;
signal \N__38842\ : std_logic;
signal \N__38835\ : std_logic;
signal \N__38832\ : std_logic;
signal \N__38829\ : std_logic;
signal \N__38826\ : std_logic;
signal \N__38823\ : std_logic;
signal \N__38822\ : std_logic;
signal \N__38821\ : std_logic;
signal \N__38820\ : std_logic;
signal \N__38817\ : std_logic;
signal \N__38814\ : std_logic;
signal \N__38809\ : std_logic;
signal \N__38808\ : std_logic;
signal \N__38807\ : std_logic;
signal \N__38806\ : std_logic;
signal \N__38803\ : std_logic;
signal \N__38802\ : std_logic;
signal \N__38799\ : std_logic;
signal \N__38796\ : std_logic;
signal \N__38791\ : std_logic;
signal \N__38788\ : std_logic;
signal \N__38785\ : std_logic;
signal \N__38782\ : std_logic;
signal \N__38779\ : std_logic;
signal \N__38774\ : std_logic;
signal \N__38771\ : std_logic;
signal \N__38766\ : std_logic;
signal \N__38763\ : std_logic;
signal \N__38760\ : std_logic;
signal \N__38757\ : std_logic;
signal \N__38754\ : std_logic;
signal \N__38751\ : std_logic;
signal \N__38742\ : std_logic;
signal \N__38739\ : std_logic;
signal \N__38736\ : std_logic;
signal \N__38733\ : std_logic;
signal \N__38730\ : std_logic;
signal \N__38727\ : std_logic;
signal \N__38726\ : std_logic;
signal \N__38723\ : std_logic;
signal \N__38720\ : std_logic;
signal \N__38715\ : std_logic;
signal \N__38712\ : std_logic;
signal \N__38709\ : std_logic;
signal \N__38706\ : std_logic;
signal \N__38703\ : std_logic;
signal \N__38700\ : std_logic;
signal \N__38699\ : std_logic;
signal \N__38696\ : std_logic;
signal \N__38693\ : std_logic;
signal \N__38690\ : std_logic;
signal \N__38687\ : std_logic;
signal \N__38682\ : std_logic;
signal \N__38679\ : std_logic;
signal \N__38676\ : std_logic;
signal \N__38675\ : std_logic;
signal \N__38674\ : std_logic;
signal \N__38673\ : std_logic;
signal \N__38670\ : std_logic;
signal \N__38667\ : std_logic;
signal \N__38666\ : std_logic;
signal \N__38665\ : std_logic;
signal \N__38664\ : std_logic;
signal \N__38661\ : std_logic;
signal \N__38658\ : std_logic;
signal \N__38657\ : std_logic;
signal \N__38656\ : std_logic;
signal \N__38653\ : std_logic;
signal \N__38650\ : std_logic;
signal \N__38643\ : std_logic;
signal \N__38638\ : std_logic;
signal \N__38637\ : std_logic;
signal \N__38634\ : std_logic;
signal \N__38631\ : std_logic;
signal \N__38626\ : std_logic;
signal \N__38621\ : std_logic;
signal \N__38618\ : std_logic;
signal \N__38607\ : std_logic;
signal \N__38604\ : std_logic;
signal \N__38601\ : std_logic;
signal \N__38598\ : std_logic;
signal \N__38597\ : std_logic;
signal \N__38596\ : std_logic;
signal \N__38593\ : std_logic;
signal \N__38588\ : std_logic;
signal \N__38583\ : std_logic;
signal \N__38580\ : std_logic;
signal \N__38577\ : std_logic;
signal \N__38576\ : std_logic;
signal \N__38573\ : std_logic;
signal \N__38570\ : std_logic;
signal \N__38567\ : std_logic;
signal \N__38566\ : std_logic;
signal \N__38561\ : std_logic;
signal \N__38558\ : std_logic;
signal \N__38555\ : std_logic;
signal \N__38550\ : std_logic;
signal \N__38547\ : std_logic;
signal \N__38544\ : std_logic;
signal \N__38541\ : std_logic;
signal \N__38538\ : std_logic;
signal \N__38535\ : std_logic;
signal \N__38532\ : std_logic;
signal \N__38529\ : std_logic;
signal \N__38526\ : std_logic;
signal \N__38523\ : std_logic;
signal \N__38520\ : std_logic;
signal \N__38519\ : std_logic;
signal \N__38518\ : std_logic;
signal \N__38515\ : std_logic;
signal \N__38510\ : std_logic;
signal \N__38505\ : std_logic;
signal \N__38502\ : std_logic;
signal \N__38499\ : std_logic;
signal \N__38496\ : std_logic;
signal \N__38493\ : std_logic;
signal \N__38490\ : std_logic;
signal \N__38487\ : std_logic;
signal \N__38484\ : std_logic;
signal \N__38481\ : std_logic;
signal \N__38480\ : std_logic;
signal \N__38479\ : std_logic;
signal \N__38476\ : std_logic;
signal \N__38473\ : std_logic;
signal \N__38470\ : std_logic;
signal \N__38467\ : std_logic;
signal \N__38464\ : std_logic;
signal \N__38461\ : std_logic;
signal \N__38458\ : std_logic;
signal \N__38455\ : std_logic;
signal \N__38452\ : std_logic;
signal \N__38445\ : std_logic;
signal \N__38442\ : std_logic;
signal \N__38439\ : std_logic;
signal \N__38436\ : std_logic;
signal \N__38433\ : std_logic;
signal \N__38430\ : std_logic;
signal \N__38429\ : std_logic;
signal \N__38426\ : std_logic;
signal \N__38425\ : std_logic;
signal \N__38422\ : std_logic;
signal \N__38419\ : std_logic;
signal \N__38416\ : std_logic;
signal \N__38413\ : std_logic;
signal \N__38406\ : std_logic;
signal \N__38403\ : std_logic;
signal \N__38400\ : std_logic;
signal \N__38397\ : std_logic;
signal \N__38394\ : std_logic;
signal \N__38391\ : std_logic;
signal \N__38388\ : std_logic;
signal \N__38385\ : std_logic;
signal \N__38382\ : std_logic;
signal \N__38379\ : std_logic;
signal \N__38376\ : std_logic;
signal \N__38375\ : std_logic;
signal \N__38374\ : std_logic;
signal \N__38373\ : std_logic;
signal \N__38372\ : std_logic;
signal \N__38369\ : std_logic;
signal \N__38366\ : std_logic;
signal \N__38363\ : std_logic;
signal \N__38360\ : std_logic;
signal \N__38357\ : std_logic;
signal \N__38352\ : std_logic;
signal \N__38347\ : std_logic;
signal \N__38344\ : std_logic;
signal \N__38339\ : std_logic;
signal \N__38336\ : std_logic;
signal \N__38333\ : std_logic;
signal \N__38328\ : std_logic;
signal \N__38325\ : std_logic;
signal \N__38322\ : std_logic;
signal \N__38319\ : std_logic;
signal \N__38318\ : std_logic;
signal \N__38317\ : std_logic;
signal \N__38316\ : std_logic;
signal \N__38315\ : std_logic;
signal \N__38312\ : std_logic;
signal \N__38311\ : std_logic;
signal \N__38308\ : std_logic;
signal \N__38305\ : std_logic;
signal \N__38304\ : std_logic;
signal \N__38303\ : std_logic;
signal \N__38302\ : std_logic;
signal \N__38301\ : std_logic;
signal \N__38298\ : std_logic;
signal \N__38295\ : std_logic;
signal \N__38292\ : std_logic;
signal \N__38285\ : std_logic;
signal \N__38282\ : std_logic;
signal \N__38279\ : std_logic;
signal \N__38278\ : std_logic;
signal \N__38277\ : std_logic;
signal \N__38276\ : std_logic;
signal \N__38273\ : std_logic;
signal \N__38270\ : std_logic;
signal \N__38269\ : std_logic;
signal \N__38268\ : std_logic;
signal \N__38263\ : std_logic;
signal \N__38260\ : std_logic;
signal \N__38257\ : std_logic;
signal \N__38254\ : std_logic;
signal \N__38251\ : std_logic;
signal \N__38248\ : std_logic;
signal \N__38243\ : std_logic;
signal \N__38240\ : std_logic;
signal \N__38239\ : std_logic;
signal \N__38238\ : std_logic;
signal \N__38237\ : std_logic;
signal \N__38234\ : std_logic;
signal \N__38231\ : std_logic;
signal \N__38228\ : std_logic;
signal \N__38223\ : std_logic;
signal \N__38222\ : std_logic;
signal \N__38221\ : std_logic;
signal \N__38220\ : std_logic;
signal \N__38219\ : std_logic;
signal \N__38218\ : std_logic;
signal \N__38217\ : std_logic;
signal \N__38216\ : std_logic;
signal \N__38215\ : std_logic;
signal \N__38214\ : std_logic;
signal \N__38213\ : std_logic;
signal \N__38212\ : std_logic;
signal \N__38211\ : std_logic;
signal \N__38208\ : std_logic;
signal \N__38203\ : std_logic;
signal \N__38196\ : std_logic;
signal \N__38189\ : std_logic;
signal \N__38184\ : std_logic;
signal \N__38179\ : std_logic;
signal \N__38176\ : std_logic;
signal \N__38161\ : std_logic;
signal \N__38152\ : std_logic;
signal \N__38147\ : std_logic;
signal \N__38138\ : std_logic;
signal \N__38127\ : std_logic;
signal \N__38124\ : std_logic;
signal \N__38121\ : std_logic;
signal \N__38118\ : std_logic;
signal \N__38115\ : std_logic;
signal \N__38112\ : std_logic;
signal \N__38109\ : std_logic;
signal \N__38106\ : std_logic;
signal \N__38103\ : std_logic;
signal \N__38100\ : std_logic;
signal \N__38097\ : std_logic;
signal \N__38094\ : std_logic;
signal \N__38091\ : std_logic;
signal \N__38088\ : std_logic;
signal \N__38085\ : std_logic;
signal \N__38082\ : std_logic;
signal \N__38079\ : std_logic;
signal \N__38078\ : std_logic;
signal \N__38077\ : std_logic;
signal \N__38074\ : std_logic;
signal \N__38071\ : std_logic;
signal \N__38068\ : std_logic;
signal \N__38065\ : std_logic;
signal \N__38062\ : std_logic;
signal \N__38059\ : std_logic;
signal \N__38056\ : std_logic;
signal \N__38053\ : std_logic;
signal \N__38050\ : std_logic;
signal \N__38047\ : std_logic;
signal \N__38044\ : std_logic;
signal \N__38041\ : std_logic;
signal \N__38034\ : std_logic;
signal \N__38031\ : std_logic;
signal \N__38028\ : std_logic;
signal \N__38025\ : std_logic;
signal \N__38022\ : std_logic;
signal \N__38019\ : std_logic;
signal \N__38016\ : std_logic;
signal \N__38013\ : std_logic;
signal \N__38010\ : std_logic;
signal \N__38007\ : std_logic;
signal \N__38004\ : std_logic;
signal \N__38001\ : std_logic;
signal \N__37998\ : std_logic;
signal \N__37995\ : std_logic;
signal \N__37992\ : std_logic;
signal \N__37989\ : std_logic;
signal \N__37986\ : std_logic;
signal \N__37983\ : std_logic;
signal \N__37980\ : std_logic;
signal \N__37977\ : std_logic;
signal \N__37974\ : std_logic;
signal \N__37971\ : std_logic;
signal \N__37968\ : std_logic;
signal \N__37965\ : std_logic;
signal \N__37962\ : std_logic;
signal \N__37959\ : std_logic;
signal \N__37956\ : std_logic;
signal \N__37953\ : std_logic;
signal \N__37950\ : std_logic;
signal \N__37947\ : std_logic;
signal \N__37944\ : std_logic;
signal \N__37941\ : std_logic;
signal \N__37938\ : std_logic;
signal \N__37935\ : std_logic;
signal \N__37934\ : std_logic;
signal \N__37931\ : std_logic;
signal \N__37928\ : std_logic;
signal \N__37925\ : std_logic;
signal \N__37922\ : std_logic;
signal \N__37919\ : std_logic;
signal \N__37914\ : std_logic;
signal \N__37911\ : std_logic;
signal \N__37908\ : std_logic;
signal \N__37905\ : std_logic;
signal \N__37904\ : std_logic;
signal \N__37901\ : std_logic;
signal \N__37898\ : std_logic;
signal \N__37895\ : std_logic;
signal \N__37890\ : std_logic;
signal \N__37887\ : std_logic;
signal \N__37884\ : std_logic;
signal \N__37881\ : std_logic;
signal \N__37880\ : std_logic;
signal \N__37879\ : std_logic;
signal \N__37878\ : std_logic;
signal \N__37877\ : std_logic;
signal \N__37876\ : std_logic;
signal \N__37875\ : std_logic;
signal \N__37874\ : std_logic;
signal \N__37873\ : std_logic;
signal \N__37870\ : std_logic;
signal \N__37869\ : std_logic;
signal \N__37868\ : std_logic;
signal \N__37867\ : std_logic;
signal \N__37866\ : std_logic;
signal \N__37865\ : std_logic;
signal \N__37864\ : std_logic;
signal \N__37863\ : std_logic;
signal \N__37848\ : std_logic;
signal \N__37845\ : std_logic;
signal \N__37844\ : std_logic;
signal \N__37843\ : std_logic;
signal \N__37840\ : std_logic;
signal \N__37825\ : std_logic;
signal \N__37824\ : std_logic;
signal \N__37823\ : std_logic;
signal \N__37820\ : std_logic;
signal \N__37817\ : std_logic;
signal \N__37814\ : std_logic;
signal \N__37811\ : std_logic;
signal \N__37810\ : std_logic;
signal \N__37809\ : std_logic;
signal \N__37808\ : std_logic;
signal \N__37807\ : std_logic;
signal \N__37806\ : std_logic;
signal \N__37805\ : std_logic;
signal \N__37804\ : std_logic;
signal \N__37803\ : std_logic;
signal \N__37798\ : std_logic;
signal \N__37795\ : std_logic;
signal \N__37792\ : std_logic;
signal \N__37789\ : std_logic;
signal \N__37784\ : std_logic;
signal \N__37781\ : std_logic;
signal \N__37768\ : std_logic;
signal \N__37765\ : std_logic;
signal \N__37762\ : std_logic;
signal \N__37759\ : std_logic;
signal \N__37754\ : std_logic;
signal \N__37749\ : std_logic;
signal \N__37742\ : std_logic;
signal \N__37731\ : std_logic;
signal \N__37728\ : std_logic;
signal \N__37725\ : std_logic;
signal \N__37722\ : std_logic;
signal \N__37719\ : std_logic;
signal \N__37716\ : std_logic;
signal \N__37713\ : std_logic;
signal \N__37710\ : std_logic;
signal \N__37707\ : std_logic;
signal \N__37706\ : std_logic;
signal \N__37705\ : std_logic;
signal \N__37702\ : std_logic;
signal \N__37701\ : std_logic;
signal \N__37700\ : std_logic;
signal \N__37699\ : std_logic;
signal \N__37698\ : std_logic;
signal \N__37695\ : std_logic;
signal \N__37694\ : std_logic;
signal \N__37691\ : std_logic;
signal \N__37690\ : std_logic;
signal \N__37689\ : std_logic;
signal \N__37688\ : std_logic;
signal \N__37685\ : std_logic;
signal \N__37682\ : std_logic;
signal \N__37675\ : std_logic;
signal \N__37672\ : std_logic;
signal \N__37669\ : std_logic;
signal \N__37666\ : std_logic;
signal \N__37659\ : std_logic;
signal \N__37658\ : std_logic;
signal \N__37657\ : std_logic;
signal \N__37656\ : std_logic;
signal \N__37655\ : std_logic;
signal \N__37654\ : std_logic;
signal \N__37653\ : std_logic;
signal \N__37652\ : std_logic;
signal \N__37651\ : std_logic;
signal \N__37650\ : std_logic;
signal \N__37649\ : std_logic;
signal \N__37648\ : std_logic;
signal \N__37647\ : std_logic;
signal \N__37646\ : std_logic;
signal \N__37645\ : std_logic;
signal \N__37644\ : std_logic;
signal \N__37643\ : std_logic;
signal \N__37642\ : std_logic;
signal \N__37641\ : std_logic;
signal \N__37640\ : std_logic;
signal \N__37635\ : std_logic;
signal \N__37632\ : std_logic;
signal \N__37627\ : std_logic;
signal \N__37622\ : std_logic;
signal \N__37613\ : std_logic;
signal \N__37604\ : std_logic;
signal \N__37589\ : std_logic;
signal \N__37580\ : std_logic;
signal \N__37575\ : std_logic;
signal \N__37570\ : std_logic;
signal \N__37557\ : std_logic;
signal \N__37554\ : std_logic;
signal \N__37551\ : std_logic;
signal \N__37548\ : std_logic;
signal \N__37545\ : std_logic;
signal \N__37542\ : std_logic;
signal \N__37539\ : std_logic;
signal \N__37536\ : std_logic;
signal \N__37533\ : std_logic;
signal \N__37530\ : std_logic;
signal \N__37527\ : std_logic;
signal \N__37524\ : std_logic;
signal \N__37521\ : std_logic;
signal \N__37518\ : std_logic;
signal \N__37515\ : std_logic;
signal \N__37512\ : std_logic;
signal \N__37509\ : std_logic;
signal \N__37506\ : std_logic;
signal \N__37503\ : std_logic;
signal \N__37500\ : std_logic;
signal \N__37497\ : std_logic;
signal \N__37494\ : std_logic;
signal \N__37491\ : std_logic;
signal \N__37488\ : std_logic;
signal \N__37485\ : std_logic;
signal \N__37482\ : std_logic;
signal \N__37479\ : std_logic;
signal \N__37476\ : std_logic;
signal \N__37473\ : std_logic;
signal \N__37470\ : std_logic;
signal \N__37467\ : std_logic;
signal \N__37464\ : std_logic;
signal \N__37461\ : std_logic;
signal \N__37458\ : std_logic;
signal \N__37455\ : std_logic;
signal \N__37452\ : std_logic;
signal \N__37449\ : std_logic;
signal \N__37446\ : std_logic;
signal \N__37443\ : std_logic;
signal \N__37440\ : std_logic;
signal \N__37437\ : std_logic;
signal \N__37434\ : std_logic;
signal \N__37431\ : std_logic;
signal \N__37428\ : std_logic;
signal \N__37425\ : std_logic;
signal \N__37422\ : std_logic;
signal \N__37419\ : std_logic;
signal \N__37416\ : std_logic;
signal \N__37413\ : std_logic;
signal \N__37410\ : std_logic;
signal \N__37407\ : std_logic;
signal \N__37404\ : std_logic;
signal \N__37401\ : std_logic;
signal \N__37398\ : std_logic;
signal \N__37395\ : std_logic;
signal \N__37392\ : std_logic;
signal \N__37389\ : std_logic;
signal \N__37386\ : std_logic;
signal \N__37383\ : std_logic;
signal \N__37380\ : std_logic;
signal \N__37377\ : std_logic;
signal \N__37374\ : std_logic;
signal \N__37371\ : std_logic;
signal \N__37368\ : std_logic;
signal \N__37365\ : std_logic;
signal \N__37362\ : std_logic;
signal \N__37359\ : std_logic;
signal \N__37356\ : std_logic;
signal \N__37353\ : std_logic;
signal \N__37350\ : std_logic;
signal \N__37347\ : std_logic;
signal \N__37344\ : std_logic;
signal \N__37341\ : std_logic;
signal \N__37338\ : std_logic;
signal \N__37335\ : std_logic;
signal \N__37332\ : std_logic;
signal \N__37329\ : std_logic;
signal \N__37326\ : std_logic;
signal \N__37323\ : std_logic;
signal \N__37320\ : std_logic;
signal \N__37317\ : std_logic;
signal \N__37314\ : std_logic;
signal \N__37311\ : std_logic;
signal \N__37308\ : std_logic;
signal \N__37305\ : std_logic;
signal \N__37302\ : std_logic;
signal \N__37299\ : std_logic;
signal \N__37296\ : std_logic;
signal \N__37293\ : std_logic;
signal \N__37290\ : std_logic;
signal \N__37287\ : std_logic;
signal \N__37284\ : std_logic;
signal \N__37281\ : std_logic;
signal \N__37278\ : std_logic;
signal \N__37275\ : std_logic;
signal \N__37272\ : std_logic;
signal \N__37269\ : std_logic;
signal \N__37266\ : std_logic;
signal \N__37263\ : std_logic;
signal \N__37260\ : std_logic;
signal \N__37257\ : std_logic;
signal \N__37254\ : std_logic;
signal \N__37251\ : std_logic;
signal \N__37248\ : std_logic;
signal \N__37245\ : std_logic;
signal \N__37242\ : std_logic;
signal \N__37239\ : std_logic;
signal \N__37236\ : std_logic;
signal \N__37233\ : std_logic;
signal \N__37230\ : std_logic;
signal \N__37227\ : std_logic;
signal \N__37224\ : std_logic;
signal \N__37221\ : std_logic;
signal \N__37218\ : std_logic;
signal \N__37215\ : std_logic;
signal \N__37212\ : std_logic;
signal \N__37209\ : std_logic;
signal \N__37206\ : std_logic;
signal \N__37203\ : std_logic;
signal \N__37200\ : std_logic;
signal \N__37197\ : std_logic;
signal \N__37194\ : std_logic;
signal \N__37191\ : std_logic;
signal \N__37188\ : std_logic;
signal \N__37185\ : std_logic;
signal \N__37182\ : std_logic;
signal \N__37179\ : std_logic;
signal \N__37176\ : std_logic;
signal \N__37173\ : std_logic;
signal \N__37170\ : std_logic;
signal \N__37169\ : std_logic;
signal \N__37168\ : std_logic;
signal \N__37165\ : std_logic;
signal \N__37162\ : std_logic;
signal \N__37161\ : std_logic;
signal \N__37160\ : std_logic;
signal \N__37159\ : std_logic;
signal \N__37156\ : std_logic;
signal \N__37153\ : std_logic;
signal \N__37150\ : std_logic;
signal \N__37149\ : std_logic;
signal \N__37148\ : std_logic;
signal \N__37145\ : std_logic;
signal \N__37140\ : std_logic;
signal \N__37137\ : std_logic;
signal \N__37132\ : std_logic;
signal \N__37127\ : std_logic;
signal \N__37116\ : std_logic;
signal \N__37113\ : std_logic;
signal \N__37110\ : std_logic;
signal \N__37109\ : std_logic;
signal \N__37108\ : std_logic;
signal \N__37107\ : std_logic;
signal \N__37106\ : std_logic;
signal \N__37103\ : std_logic;
signal \N__37100\ : std_logic;
signal \N__37097\ : std_logic;
signal \N__37092\ : std_logic;
signal \N__37083\ : std_logic;
signal \N__37082\ : std_logic;
signal \N__37077\ : std_logic;
signal \N__37074\ : std_logic;
signal \N__37071\ : std_logic;
signal \N__37068\ : std_logic;
signal \N__37065\ : std_logic;
signal \N__37064\ : std_logic;
signal \N__37061\ : std_logic;
signal \N__37058\ : std_logic;
signal \N__37053\ : std_logic;
signal \N__37050\ : std_logic;
signal \N__37049\ : std_logic;
signal \N__37048\ : std_logic;
signal \N__37045\ : std_logic;
signal \N__37042\ : std_logic;
signal \N__37037\ : std_logic;
signal \N__37032\ : std_logic;
signal \N__37031\ : std_logic;
signal \N__37028\ : std_logic;
signal \N__37025\ : std_logic;
signal \N__37020\ : std_logic;
signal \N__37019\ : std_logic;
signal \N__37016\ : std_logic;
signal \N__37013\ : std_logic;
signal \N__37008\ : std_logic;
signal \N__37005\ : std_logic;
signal \N__37002\ : std_logic;
signal \N__36999\ : std_logic;
signal \N__36996\ : std_logic;
signal \N__36993\ : std_logic;
signal \N__36990\ : std_logic;
signal \N__36987\ : std_logic;
signal \N__36984\ : std_logic;
signal \N__36981\ : std_logic;
signal \N__36978\ : std_logic;
signal \N__36975\ : std_logic;
signal \N__36972\ : std_logic;
signal \N__36969\ : std_logic;
signal \N__36968\ : std_logic;
signal \N__36967\ : std_logic;
signal \N__36964\ : std_logic;
signal \N__36961\ : std_logic;
signal \N__36960\ : std_logic;
signal \N__36959\ : std_logic;
signal \N__36958\ : std_logic;
signal \N__36957\ : std_logic;
signal \N__36956\ : std_logic;
signal \N__36955\ : std_logic;
signal \N__36954\ : std_logic;
signal \N__36951\ : std_logic;
signal \N__36948\ : std_logic;
signal \N__36939\ : std_logic;
signal \N__36934\ : std_logic;
signal \N__36929\ : std_logic;
signal \N__36926\ : std_logic;
signal \N__36923\ : std_logic;
signal \N__36918\ : std_logic;
signal \N__36909\ : std_logic;
signal \N__36908\ : std_logic;
signal \N__36905\ : std_logic;
signal \N__36904\ : std_logic;
signal \N__36901\ : std_logic;
signal \N__36900\ : std_logic;
signal \N__36897\ : std_logic;
signal \N__36894\ : std_logic;
signal \N__36891\ : std_logic;
signal \N__36888\ : std_logic;
signal \N__36883\ : std_logic;
signal \N__36880\ : std_logic;
signal \N__36873\ : std_logic;
signal \N__36870\ : std_logic;
signal \N__36869\ : std_logic;
signal \N__36868\ : std_logic;
signal \N__36865\ : std_logic;
signal \N__36862\ : std_logic;
signal \N__36859\ : std_logic;
signal \N__36856\ : std_logic;
signal \N__36851\ : std_logic;
signal \N__36846\ : std_logic;
signal \N__36843\ : std_logic;
signal \N__36840\ : std_logic;
signal \N__36839\ : std_logic;
signal \N__36838\ : std_logic;
signal \N__36837\ : std_logic;
signal \N__36836\ : std_logic;
signal \N__36831\ : std_logic;
signal \N__36828\ : std_logic;
signal \N__36825\ : std_logic;
signal \N__36822\ : std_logic;
signal \N__36819\ : std_logic;
signal \N__36816\ : std_logic;
signal \N__36807\ : std_logic;
signal \N__36804\ : std_logic;
signal \N__36801\ : std_logic;
signal \N__36798\ : std_logic;
signal \N__36795\ : std_logic;
signal \N__36792\ : std_logic;
signal \N__36789\ : std_logic;
signal \N__36786\ : std_logic;
signal \N__36785\ : std_logic;
signal \N__36780\ : std_logic;
signal \N__36777\ : std_logic;
signal \N__36774\ : std_logic;
signal \N__36771\ : std_logic;
signal \N__36770\ : std_logic;
signal \N__36767\ : std_logic;
signal \N__36764\ : std_logic;
signal \N__36759\ : std_logic;
signal \N__36756\ : std_logic;
signal \N__36753\ : std_logic;
signal \N__36750\ : std_logic;
signal \N__36747\ : std_logic;
signal \N__36744\ : std_logic;
signal \N__36741\ : std_logic;
signal \N__36738\ : std_logic;
signal \N__36737\ : std_logic;
signal \N__36736\ : std_logic;
signal \N__36735\ : std_logic;
signal \N__36734\ : std_logic;
signal \N__36731\ : std_logic;
signal \N__36722\ : std_logic;
signal \N__36717\ : std_logic;
signal \N__36716\ : std_logic;
signal \N__36715\ : std_logic;
signal \N__36714\ : std_logic;
signal \N__36711\ : std_logic;
signal \N__36708\ : std_logic;
signal \N__36703\ : std_logic;
signal \N__36696\ : std_logic;
signal \N__36695\ : std_logic;
signal \N__36690\ : std_logic;
signal \N__36689\ : std_logic;
signal \N__36686\ : std_logic;
signal \N__36683\ : std_logic;
signal \N__36678\ : std_logic;
signal \N__36677\ : std_logic;
signal \N__36676\ : std_logic;
signal \N__36675\ : std_logic;
signal \N__36672\ : std_logic;
signal \N__36665\ : std_logic;
signal \N__36662\ : std_logic;
signal \N__36657\ : std_logic;
signal \N__36654\ : std_logic;
signal \N__36651\ : std_logic;
signal \N__36648\ : std_logic;
signal \N__36647\ : std_logic;
signal \N__36644\ : std_logic;
signal \N__36643\ : std_logic;
signal \N__36642\ : std_logic;
signal \N__36641\ : std_logic;
signal \N__36640\ : std_logic;
signal \N__36639\ : std_logic;
signal \N__36638\ : std_logic;
signal \N__36635\ : std_logic;
signal \N__36634\ : std_logic;
signal \N__36631\ : std_logic;
signal \N__36626\ : std_logic;
signal \N__36623\ : std_logic;
signal \N__36616\ : std_logic;
signal \N__36611\ : std_logic;
signal \N__36600\ : std_logic;
signal \N__36599\ : std_logic;
signal \N__36596\ : std_logic;
signal \N__36595\ : std_logic;
signal \N__36592\ : std_logic;
signal \N__36589\ : std_logic;
signal \N__36586\ : std_logic;
signal \N__36579\ : std_logic;
signal \N__36576\ : std_logic;
signal \N__36573\ : std_logic;
signal \N__36570\ : std_logic;
signal \N__36567\ : std_logic;
signal \N__36564\ : std_logic;
signal \N__36561\ : std_logic;
signal \N__36558\ : std_logic;
signal \N__36555\ : std_logic;
signal \N__36552\ : std_logic;
signal \N__36549\ : std_logic;
signal \N__36546\ : std_logic;
signal \N__36543\ : std_logic;
signal \N__36540\ : std_logic;
signal \N__36537\ : std_logic;
signal \N__36534\ : std_logic;
signal \N__36531\ : std_logic;
signal \N__36530\ : std_logic;
signal \N__36527\ : std_logic;
signal \N__36524\ : std_logic;
signal \N__36519\ : std_logic;
signal \N__36516\ : std_logic;
signal \N__36513\ : std_logic;
signal \N__36510\ : std_logic;
signal \N__36507\ : std_logic;
signal \N__36504\ : std_logic;
signal \N__36503\ : std_logic;
signal \N__36500\ : std_logic;
signal \N__36497\ : std_logic;
signal \N__36494\ : std_logic;
signal \N__36491\ : std_logic;
signal \N__36486\ : std_logic;
signal \N__36483\ : std_logic;
signal \N__36480\ : std_logic;
signal \N__36477\ : std_logic;
signal \N__36474\ : std_logic;
signal \N__36473\ : std_logic;
signal \N__36472\ : std_logic;
signal \N__36469\ : std_logic;
signal \N__36466\ : std_logic;
signal \N__36463\ : std_logic;
signal \N__36460\ : std_logic;
signal \N__36453\ : std_logic;
signal \N__36450\ : std_logic;
signal \N__36449\ : std_logic;
signal \N__36444\ : std_logic;
signal \N__36441\ : std_logic;
signal \N__36438\ : std_logic;
signal \N__36435\ : std_logic;
signal \N__36432\ : std_logic;
signal \N__36431\ : std_logic;
signal \N__36428\ : std_logic;
signal \N__36425\ : std_logic;
signal \N__36422\ : std_logic;
signal \N__36417\ : std_logic;
signal \N__36414\ : std_logic;
signal \N__36411\ : std_logic;
signal \N__36408\ : std_logic;
signal \N__36405\ : std_logic;
signal \N__36402\ : std_logic;
signal \N__36399\ : std_logic;
signal \N__36396\ : std_logic;
signal \N__36393\ : std_logic;
signal \N__36390\ : std_logic;
signal \N__36387\ : std_logic;
signal \N__36384\ : std_logic;
signal \N__36381\ : std_logic;
signal \N__36378\ : std_logic;
signal \N__36375\ : std_logic;
signal \N__36372\ : std_logic;
signal \N__36369\ : std_logic;
signal \N__36366\ : std_logic;
signal \N__36363\ : std_logic;
signal \N__36362\ : std_logic;
signal \N__36359\ : std_logic;
signal \N__36356\ : std_logic;
signal \N__36355\ : std_logic;
signal \N__36354\ : std_logic;
signal \N__36351\ : std_logic;
signal \N__36348\ : std_logic;
signal \N__36345\ : std_logic;
signal \N__36342\ : std_logic;
signal \N__36339\ : std_logic;
signal \N__36336\ : std_logic;
signal \N__36333\ : std_logic;
signal \N__36324\ : std_logic;
signal \N__36321\ : std_logic;
signal \N__36318\ : std_logic;
signal \N__36317\ : std_logic;
signal \N__36314\ : std_logic;
signal \N__36311\ : std_logic;
signal \N__36306\ : std_logic;
signal \N__36305\ : std_logic;
signal \N__36302\ : std_logic;
signal \N__36299\ : std_logic;
signal \N__36296\ : std_logic;
signal \N__36295\ : std_logic;
signal \N__36294\ : std_logic;
signal \N__36291\ : std_logic;
signal \N__36288\ : std_logic;
signal \N__36283\ : std_logic;
signal \N__36280\ : std_logic;
signal \N__36273\ : std_logic;
signal \N__36272\ : std_logic;
signal \N__36269\ : std_logic;
signal \N__36268\ : std_logic;
signal \N__36265\ : std_logic;
signal \N__36260\ : std_logic;
signal \N__36259\ : std_logic;
signal \N__36256\ : std_logic;
signal \N__36253\ : std_logic;
signal \N__36250\ : std_logic;
signal \N__36247\ : std_logic;
signal \N__36244\ : std_logic;
signal \N__36237\ : std_logic;
signal \N__36236\ : std_logic;
signal \N__36235\ : std_logic;
signal \N__36228\ : std_logic;
signal \N__36225\ : std_logic;
signal \N__36222\ : std_logic;
signal \N__36221\ : std_logic;
signal \N__36220\ : std_logic;
signal \N__36219\ : std_logic;
signal \N__36218\ : std_logic;
signal \N__36215\ : std_logic;
signal \N__36206\ : std_logic;
signal \N__36201\ : std_logic;
signal \N__36198\ : std_logic;
signal \N__36195\ : std_logic;
signal \N__36192\ : std_logic;
signal \N__36189\ : std_logic;
signal \N__36186\ : std_logic;
signal \N__36183\ : std_logic;
signal \N__36182\ : std_logic;
signal \N__36179\ : std_logic;
signal \N__36176\ : std_logic;
signal \N__36171\ : std_logic;
signal \N__36168\ : std_logic;
signal \N__36165\ : std_logic;
signal \N__36162\ : std_logic;
signal \N__36159\ : std_logic;
signal \N__36158\ : std_logic;
signal \N__36155\ : std_logic;
signal \N__36152\ : std_logic;
signal \N__36147\ : std_logic;
signal \N__36144\ : std_logic;
signal \N__36141\ : std_logic;
signal \N__36140\ : std_logic;
signal \N__36137\ : std_logic;
signal \N__36134\ : std_logic;
signal \N__36129\ : std_logic;
signal \N__36126\ : std_logic;
signal \N__36123\ : std_logic;
signal \N__36120\ : std_logic;
signal \N__36117\ : std_logic;
signal \N__36114\ : std_logic;
signal \N__36113\ : std_logic;
signal \N__36110\ : std_logic;
signal \N__36107\ : std_logic;
signal \N__36104\ : std_logic;
signal \N__36101\ : std_logic;
signal \N__36098\ : std_logic;
signal \N__36095\ : std_logic;
signal \N__36092\ : std_logic;
signal \N__36089\ : std_logic;
signal \N__36086\ : std_logic;
signal \N__36083\ : std_logic;
signal \N__36080\ : std_logic;
signal \N__36077\ : std_logic;
signal \N__36074\ : std_logic;
signal \N__36071\ : std_logic;
signal \N__36068\ : std_logic;
signal \N__36065\ : std_logic;
signal \N__36062\ : std_logic;
signal \N__36059\ : std_logic;
signal \N__36056\ : std_logic;
signal \N__36053\ : std_logic;
signal \N__36050\ : std_logic;
signal \N__36047\ : std_logic;
signal \N__36044\ : std_logic;
signal \N__36041\ : std_logic;
signal \N__36038\ : std_logic;
signal \N__36035\ : std_logic;
signal \N__36032\ : std_logic;
signal \N__36029\ : std_logic;
signal \N__36026\ : std_logic;
signal \N__36023\ : std_logic;
signal \N__36020\ : std_logic;
signal \N__36017\ : std_logic;
signal \N__36014\ : std_logic;
signal \N__36011\ : std_logic;
signal \N__36006\ : std_logic;
signal \N__36003\ : std_logic;
signal \N__36000\ : std_logic;
signal \N__35997\ : std_logic;
signal \N__35996\ : std_logic;
signal \N__35993\ : std_logic;
signal \N__35992\ : std_logic;
signal \N__35991\ : std_logic;
signal \N__35990\ : std_logic;
signal \N__35989\ : std_logic;
signal \N__35988\ : std_logic;
signal \N__35987\ : std_logic;
signal \N__35986\ : std_logic;
signal \N__35983\ : std_logic;
signal \N__35974\ : std_logic;
signal \N__35973\ : std_logic;
signal \N__35968\ : std_logic;
signal \N__35963\ : std_logic;
signal \N__35960\ : std_logic;
signal \N__35957\ : std_logic;
signal \N__35954\ : std_logic;
signal \N__35949\ : std_logic;
signal \N__35944\ : std_logic;
signal \N__35941\ : std_logic;
signal \N__35938\ : std_logic;
signal \N__35935\ : std_logic;
signal \N__35930\ : std_logic;
signal \N__35925\ : std_logic;
signal \N__35922\ : std_logic;
signal \N__35919\ : std_logic;
signal \N__35916\ : std_logic;
signal \N__35915\ : std_logic;
signal \N__35912\ : std_logic;
signal \N__35909\ : std_logic;
signal \N__35906\ : std_logic;
signal \N__35903\ : std_logic;
signal \N__35900\ : std_logic;
signal \N__35897\ : std_logic;
signal \N__35892\ : std_logic;
signal \N__35889\ : std_logic;
signal \N__35888\ : std_logic;
signal \N__35885\ : std_logic;
signal \N__35882\ : std_logic;
signal \N__35881\ : std_logic;
signal \N__35878\ : std_logic;
signal \N__35875\ : std_logic;
signal \N__35872\ : std_logic;
signal \N__35869\ : std_logic;
signal \N__35862\ : std_logic;
signal \N__35861\ : std_logic;
signal \N__35860\ : std_logic;
signal \N__35857\ : std_logic;
signal \N__35856\ : std_logic;
signal \N__35855\ : std_logic;
signal \N__35854\ : std_logic;
signal \N__35853\ : std_logic;
signal \N__35848\ : std_logic;
signal \N__35845\ : std_logic;
signal \N__35838\ : std_logic;
signal \N__35835\ : std_logic;
signal \N__35832\ : std_logic;
signal \N__35829\ : std_logic;
signal \N__35826\ : std_logic;
signal \N__35823\ : std_logic;
signal \N__35820\ : std_logic;
signal \N__35819\ : std_logic;
signal \N__35818\ : std_logic;
signal \N__35813\ : std_logic;
signal \N__35808\ : std_logic;
signal \N__35803\ : std_logic;
signal \N__35796\ : std_logic;
signal \N__35795\ : std_logic;
signal \N__35792\ : std_logic;
signal \N__35789\ : std_logic;
signal \N__35786\ : std_logic;
signal \N__35783\ : std_logic;
signal \N__35780\ : std_logic;
signal \N__35777\ : std_logic;
signal \N__35774\ : std_logic;
signal \N__35771\ : std_logic;
signal \N__35768\ : std_logic;
signal \N__35763\ : std_logic;
signal \N__35762\ : std_logic;
signal \N__35761\ : std_logic;
signal \N__35758\ : std_logic;
signal \N__35757\ : std_logic;
signal \N__35756\ : std_logic;
signal \N__35755\ : std_logic;
signal \N__35752\ : std_logic;
signal \N__35749\ : std_logic;
signal \N__35748\ : std_logic;
signal \N__35743\ : std_logic;
signal \N__35738\ : std_logic;
signal \N__35735\ : std_logic;
signal \N__35732\ : std_logic;
signal \N__35729\ : std_logic;
signal \N__35726\ : std_logic;
signal \N__35725\ : std_logic;
signal \N__35724\ : std_logic;
signal \N__35719\ : std_logic;
signal \N__35716\ : std_logic;
signal \N__35711\ : std_logic;
signal \N__35708\ : std_logic;
signal \N__35705\ : std_logic;
signal \N__35700\ : std_logic;
signal \N__35691\ : std_logic;
signal \N__35688\ : std_logic;
signal \N__35685\ : std_logic;
signal \N__35682\ : std_logic;
signal \N__35681\ : std_logic;
signal \N__35680\ : std_logic;
signal \N__35677\ : std_logic;
signal \N__35672\ : std_logic;
signal \N__35667\ : std_logic;
signal \N__35664\ : std_logic;
signal \N__35661\ : std_logic;
signal \N__35658\ : std_logic;
signal \N__35655\ : std_logic;
signal \N__35652\ : std_logic;
signal \N__35651\ : std_logic;
signal \N__35648\ : std_logic;
signal \N__35645\ : std_logic;
signal \N__35642\ : std_logic;
signal \N__35639\ : std_logic;
signal \N__35636\ : std_logic;
signal \N__35631\ : std_logic;
signal \N__35628\ : std_logic;
signal \N__35625\ : std_logic;
signal \N__35622\ : std_logic;
signal \N__35619\ : std_logic;
signal \N__35616\ : std_logic;
signal \N__35613\ : std_logic;
signal \N__35610\ : std_logic;
signal \N__35607\ : std_logic;
signal \N__35604\ : std_logic;
signal \N__35603\ : std_logic;
signal \N__35600\ : std_logic;
signal \N__35597\ : std_logic;
signal \N__35594\ : std_logic;
signal \N__35589\ : std_logic;
signal \N__35586\ : std_logic;
signal \N__35583\ : std_logic;
signal \N__35580\ : std_logic;
signal \N__35577\ : std_logic;
signal \N__35574\ : std_logic;
signal \N__35573\ : std_logic;
signal \N__35570\ : std_logic;
signal \N__35567\ : std_logic;
signal \N__35564\ : std_logic;
signal \N__35561\ : std_logic;
signal \N__35558\ : std_logic;
signal \N__35553\ : std_logic;
signal \N__35550\ : std_logic;
signal \N__35547\ : std_logic;
signal \N__35544\ : std_logic;
signal \N__35541\ : std_logic;
signal \N__35538\ : std_logic;
signal \N__35537\ : std_logic;
signal \N__35534\ : std_logic;
signal \N__35533\ : std_logic;
signal \N__35530\ : std_logic;
signal \N__35527\ : std_logic;
signal \N__35524\ : std_logic;
signal \N__35519\ : std_logic;
signal \N__35516\ : std_logic;
signal \N__35513\ : std_logic;
signal \N__35508\ : std_logic;
signal \N__35505\ : std_logic;
signal \N__35502\ : std_logic;
signal \N__35499\ : std_logic;
signal \N__35496\ : std_logic;
signal \N__35493\ : std_logic;
signal \N__35490\ : std_logic;
signal \N__35487\ : std_logic;
signal \N__35484\ : std_logic;
signal \N__35483\ : std_logic;
signal \N__35482\ : std_logic;
signal \N__35481\ : std_logic;
signal \N__35474\ : std_logic;
signal \N__35471\ : std_logic;
signal \N__35468\ : std_logic;
signal \N__35465\ : std_logic;
signal \N__35464\ : std_logic;
signal \N__35461\ : std_logic;
signal \N__35458\ : std_logic;
signal \N__35457\ : std_logic;
signal \N__35454\ : std_logic;
signal \N__35451\ : std_logic;
signal \N__35448\ : std_logic;
signal \N__35445\ : std_logic;
signal \N__35442\ : std_logic;
signal \N__35439\ : std_logic;
signal \N__35436\ : std_logic;
signal \N__35433\ : std_logic;
signal \N__35430\ : std_logic;
signal \N__35427\ : std_logic;
signal \N__35424\ : std_logic;
signal \N__35421\ : std_logic;
signal \N__35418\ : std_logic;
signal \N__35415\ : std_logic;
signal \N__35410\ : std_logic;
signal \N__35407\ : std_logic;
signal \N__35400\ : std_logic;
signal \N__35397\ : std_logic;
signal \N__35396\ : std_logic;
signal \N__35395\ : std_logic;
signal \N__35394\ : std_logic;
signal \N__35391\ : std_logic;
signal \N__35388\ : std_logic;
signal \N__35383\ : std_logic;
signal \N__35380\ : std_logic;
signal \N__35375\ : std_logic;
signal \N__35370\ : std_logic;
signal \N__35367\ : std_logic;
signal \N__35364\ : std_logic;
signal \N__35361\ : std_logic;
signal \N__35360\ : std_logic;
signal \N__35357\ : std_logic;
signal \N__35354\ : std_logic;
signal \N__35351\ : std_logic;
signal \N__35348\ : std_logic;
signal \N__35343\ : std_logic;
signal \N__35340\ : std_logic;
signal \N__35337\ : std_logic;
signal \N__35334\ : std_logic;
signal \N__35331\ : std_logic;
signal \N__35330\ : std_logic;
signal \N__35327\ : std_logic;
signal \N__35324\ : std_logic;
signal \N__35321\ : std_logic;
signal \N__35316\ : std_logic;
signal \N__35313\ : std_logic;
signal \N__35310\ : std_logic;
signal \N__35307\ : std_logic;
signal \N__35304\ : std_logic;
signal \N__35303\ : std_logic;
signal \N__35300\ : std_logic;
signal \N__35297\ : std_logic;
signal \N__35294\ : std_logic;
signal \N__35291\ : std_logic;
signal \N__35288\ : std_logic;
signal \N__35283\ : std_logic;
signal \N__35280\ : std_logic;
signal \N__35277\ : std_logic;
signal \N__35274\ : std_logic;
signal \N__35271\ : std_logic;
signal \N__35268\ : std_logic;
signal \N__35265\ : std_logic;
signal \N__35264\ : std_logic;
signal \N__35261\ : std_logic;
signal \N__35258\ : std_logic;
signal \N__35255\ : std_logic;
signal \N__35250\ : std_logic;
signal \N__35247\ : std_logic;
signal \N__35244\ : std_logic;
signal \N__35241\ : std_logic;
signal \N__35238\ : std_logic;
signal \N__35235\ : std_logic;
signal \N__35234\ : std_logic;
signal \N__35231\ : std_logic;
signal \N__35228\ : std_logic;
signal \N__35225\ : std_logic;
signal \N__35220\ : std_logic;
signal \N__35217\ : std_logic;
signal \N__35214\ : std_logic;
signal \N__35211\ : std_logic;
signal \N__35208\ : std_logic;
signal \N__35205\ : std_logic;
signal \N__35202\ : std_logic;
signal \N__35199\ : std_logic;
signal \N__35198\ : std_logic;
signal \N__35195\ : std_logic;
signal \N__35192\ : std_logic;
signal \N__35189\ : std_logic;
signal \N__35184\ : std_logic;
signal \N__35181\ : std_logic;
signal \N__35178\ : std_logic;
signal \N__35177\ : std_logic;
signal \N__35174\ : std_logic;
signal \N__35171\ : std_logic;
signal \N__35168\ : std_logic;
signal \N__35163\ : std_logic;
signal \N__35160\ : std_logic;
signal \N__35157\ : std_logic;
signal \N__35154\ : std_logic;
signal \N__35151\ : std_logic;
signal \N__35148\ : std_logic;
signal \N__35145\ : std_logic;
signal \N__35142\ : std_logic;
signal \N__35139\ : std_logic;
signal \N__35136\ : std_logic;
signal \N__35133\ : std_logic;
signal \N__35130\ : std_logic;
signal \N__35127\ : std_logic;
signal \N__35124\ : std_logic;
signal \N__35121\ : std_logic;
signal \N__35118\ : std_logic;
signal \N__35115\ : std_logic;
signal \N__35112\ : std_logic;
signal \N__35109\ : std_logic;
signal \N__35106\ : std_logic;
signal \N__35103\ : std_logic;
signal \N__35100\ : std_logic;
signal \N__35099\ : std_logic;
signal \N__35096\ : std_logic;
signal \N__35093\ : std_logic;
signal \N__35090\ : std_logic;
signal \N__35087\ : std_logic;
signal \N__35084\ : std_logic;
signal \N__35079\ : std_logic;
signal \N__35076\ : std_logic;
signal \N__35073\ : std_logic;
signal \N__35070\ : std_logic;
signal \N__35067\ : std_logic;
signal \N__35064\ : std_logic;
signal \N__35061\ : std_logic;
signal \N__35060\ : std_logic;
signal \N__35057\ : std_logic;
signal \N__35054\ : std_logic;
signal \N__35051\ : std_logic;
signal \N__35048\ : std_logic;
signal \N__35045\ : std_logic;
signal \N__35040\ : std_logic;
signal \N__35037\ : std_logic;
signal \N__35034\ : std_logic;
signal \N__35031\ : std_logic;
signal \N__35028\ : std_logic;
signal \N__35025\ : std_logic;
signal \N__35022\ : std_logic;
signal \N__35019\ : std_logic;
signal \N__35018\ : std_logic;
signal \N__35015\ : std_logic;
signal \N__35012\ : std_logic;
signal \N__35009\ : std_logic;
signal \N__35004\ : std_logic;
signal \N__35001\ : std_logic;
signal \N__34998\ : std_logic;
signal \N__34995\ : std_logic;
signal \N__34992\ : std_logic;
signal \N__34989\ : std_logic;
signal \N__34988\ : std_logic;
signal \N__34985\ : std_logic;
signal \N__34982\ : std_logic;
signal \N__34979\ : std_logic;
signal \N__34976\ : std_logic;
signal \N__34973\ : std_logic;
signal \N__34968\ : std_logic;
signal \N__34965\ : std_logic;
signal \N__34962\ : std_logic;
signal \N__34959\ : std_logic;
signal \N__34956\ : std_logic;
signal \N__34953\ : std_logic;
signal \N__34950\ : std_logic;
signal \N__34947\ : std_logic;
signal \N__34944\ : std_logic;
signal \N__34943\ : std_logic;
signal \N__34940\ : std_logic;
signal \N__34937\ : std_logic;
signal \N__34934\ : std_logic;
signal \N__34931\ : std_logic;
signal \N__34928\ : std_logic;
signal \N__34923\ : std_logic;
signal \N__34920\ : std_logic;
signal \N__34917\ : std_logic;
signal \N__34914\ : std_logic;
signal \N__34911\ : std_logic;
signal \N__34910\ : std_logic;
signal \N__34907\ : std_logic;
signal \N__34904\ : std_logic;
signal \N__34901\ : std_logic;
signal \N__34898\ : std_logic;
signal \N__34895\ : std_logic;
signal \N__34890\ : std_logic;
signal \N__34887\ : std_logic;
signal \N__34884\ : std_logic;
signal \N__34881\ : std_logic;
signal \N__34878\ : std_logic;
signal \N__34875\ : std_logic;
signal \N__34872\ : std_logic;
signal \N__34869\ : std_logic;
signal \N__34866\ : std_logic;
signal \N__34863\ : std_logic;
signal \N__34860\ : std_logic;
signal \N__34857\ : std_logic;
signal \N__34856\ : std_logic;
signal \N__34853\ : std_logic;
signal \N__34852\ : std_logic;
signal \N__34851\ : std_logic;
signal \N__34848\ : std_logic;
signal \N__34845\ : std_logic;
signal \N__34844\ : std_logic;
signal \N__34843\ : std_logic;
signal \N__34840\ : std_logic;
signal \N__34837\ : std_logic;
signal \N__34832\ : std_logic;
signal \N__34827\ : std_logic;
signal \N__34818\ : std_logic;
signal \N__34815\ : std_logic;
signal \N__34812\ : std_logic;
signal \N__34809\ : std_logic;
signal \N__34806\ : std_logic;
signal \N__34803\ : std_logic;
signal \N__34800\ : std_logic;
signal \N__34797\ : std_logic;
signal \N__34794\ : std_logic;
signal \N__34791\ : std_logic;
signal \N__34788\ : std_logic;
signal \N__34785\ : std_logic;
signal \N__34782\ : std_logic;
signal \N__34779\ : std_logic;
signal \N__34776\ : std_logic;
signal \N__34773\ : std_logic;
signal \N__34770\ : std_logic;
signal \N__34767\ : std_logic;
signal \N__34764\ : std_logic;
signal \N__34761\ : std_logic;
signal \N__34758\ : std_logic;
signal \N__34755\ : std_logic;
signal \N__34752\ : std_logic;
signal \N__34749\ : std_logic;
signal \N__34746\ : std_logic;
signal \N__34743\ : std_logic;
signal \N__34740\ : std_logic;
signal \N__34737\ : std_logic;
signal \N__34734\ : std_logic;
signal \N__34731\ : std_logic;
signal \N__34728\ : std_logic;
signal \N__34725\ : std_logic;
signal \N__34722\ : std_logic;
signal \N__34719\ : std_logic;
signal \N__34716\ : std_logic;
signal \N__34713\ : std_logic;
signal \N__34710\ : std_logic;
signal \N__34707\ : std_logic;
signal \N__34704\ : std_logic;
signal \N__34701\ : std_logic;
signal \N__34698\ : std_logic;
signal \N__34695\ : std_logic;
signal \N__34692\ : std_logic;
signal \N__34689\ : std_logic;
signal \N__34686\ : std_logic;
signal \N__34683\ : std_logic;
signal \N__34680\ : std_logic;
signal \N__34677\ : std_logic;
signal \N__34674\ : std_logic;
signal \N__34671\ : std_logic;
signal \N__34670\ : std_logic;
signal \N__34667\ : std_logic;
signal \N__34662\ : std_logic;
signal \N__34659\ : std_logic;
signal \N__34656\ : std_logic;
signal \N__34655\ : std_logic;
signal \N__34654\ : std_logic;
signal \N__34651\ : std_logic;
signal \N__34646\ : std_logic;
signal \N__34641\ : std_logic;
signal \N__34640\ : std_logic;
signal \N__34639\ : std_logic;
signal \N__34636\ : std_logic;
signal \N__34633\ : std_logic;
signal \N__34630\ : std_logic;
signal \N__34629\ : std_logic;
signal \N__34626\ : std_logic;
signal \N__34621\ : std_logic;
signal \N__34618\ : std_logic;
signal \N__34615\ : std_logic;
signal \N__34612\ : std_logic;
signal \N__34609\ : std_logic;
signal \N__34604\ : std_logic;
signal \N__34599\ : std_logic;
signal \N__34598\ : std_logic;
signal \N__34597\ : std_logic;
signal \N__34594\ : std_logic;
signal \N__34589\ : std_logic;
signal \N__34584\ : std_logic;
signal \N__34581\ : std_logic;
signal \N__34578\ : std_logic;
signal \N__34575\ : std_logic;
signal \N__34572\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34566\ : std_logic;
signal \N__34563\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34557\ : std_logic;
signal \N__34556\ : std_logic;
signal \N__34555\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34540\ : std_logic;
signal \N__34537\ : std_logic;
signal \N__34532\ : std_logic;
signal \N__34529\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34521\ : std_logic;
signal \N__34518\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34512\ : std_logic;
signal \N__34511\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34505\ : std_logic;
signal \N__34502\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34494\ : std_logic;
signal \N__34491\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34485\ : std_logic;
signal \N__34482\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34476\ : std_logic;
signal \N__34473\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34467\ : std_logic;
signal \N__34464\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34458\ : std_logic;
signal \N__34457\ : std_logic;
signal \N__34456\ : std_logic;
signal \N__34455\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34450\ : std_logic;
signal \N__34449\ : std_logic;
signal \N__34442\ : std_logic;
signal \N__34433\ : std_logic;
signal \N__34428\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34422\ : std_logic;
signal \N__34421\ : std_logic;
signal \N__34420\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34414\ : std_logic;
signal \N__34411\ : std_logic;
signal \N__34404\ : std_logic;
signal \N__34403\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34397\ : std_logic;
signal \N__34392\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34386\ : std_logic;
signal \N__34383\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34376\ : std_logic;
signal \N__34375\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34369\ : std_logic;
signal \N__34366\ : std_logic;
signal \N__34359\ : std_logic;
signal \N__34358\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34351\ : std_logic;
signal \N__34348\ : std_logic;
signal \N__34343\ : std_logic;
signal \N__34340\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34334\ : std_logic;
signal \N__34333\ : std_logic;
signal \N__34332\ : std_logic;
signal \N__34331\ : std_logic;
signal \N__34330\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34314\ : std_logic;
signal \N__34313\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34307\ : std_logic;
signal \N__34302\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34296\ : std_logic;
signal \N__34295\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34289\ : std_logic;
signal \N__34286\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34280\ : std_logic;
signal \N__34277\ : std_logic;
signal \N__34276\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34269\ : std_logic;
signal \N__34266\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34260\ : std_logic;
signal \N__34257\ : std_logic;
signal \N__34248\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34244\ : std_logic;
signal \N__34241\ : std_logic;
signal \N__34240\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34234\ : std_logic;
signal \N__34231\ : std_logic;
signal \N__34224\ : std_logic;
signal \N__34221\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34217\ : std_logic;
signal \N__34216\ : std_logic;
signal \N__34213\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34207\ : std_logic;
signal \N__34204\ : std_logic;
signal \N__34197\ : std_logic;
signal \N__34194\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34190\ : std_logic;
signal \N__34189\ : std_logic;
signal \N__34186\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34180\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34170\ : std_logic;
signal \N__34169\ : std_logic;
signal \N__34168\ : std_logic;
signal \N__34167\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34163\ : std_logic;
signal \N__34154\ : std_logic;
signal \N__34149\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34143\ : std_logic;
signal \N__34140\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34132\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34126\ : std_logic;
signal \N__34125\ : std_logic;
signal \N__34122\ : std_logic;
signal \N__34117\ : std_logic;
signal \N__34116\ : std_logic;
signal \N__34113\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34107\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34099\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34091\ : std_logic;
signal \N__34086\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34080\ : std_logic;
signal \N__34077\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34071\ : std_logic;
signal \N__34068\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34062\ : std_logic;
signal \N__34059\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34053\ : std_logic;
signal \N__34050\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34046\ : std_logic;
signal \N__34043\ : std_logic;
signal \N__34040\ : std_logic;
signal \N__34037\ : std_logic;
signal \N__34034\ : std_logic;
signal \N__34031\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34017\ : std_logic;
signal \N__34014\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34008\ : std_logic;
signal \N__34005\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33994\ : std_logic;
signal \N__33991\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33980\ : std_logic;
signal \N__33977\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33971\ : std_logic;
signal \N__33968\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33959\ : std_logic;
signal \N__33956\ : std_logic;
signal \N__33951\ : std_logic;
signal \N__33950\ : std_logic;
signal \N__33949\ : std_logic;
signal \N__33948\ : std_logic;
signal \N__33947\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33938\ : std_logic;
signal \N__33937\ : std_logic;
signal \N__33936\ : std_logic;
signal \N__33935\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33926\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33922\ : std_logic;
signal \N__33921\ : std_logic;
signal \N__33920\ : std_logic;
signal \N__33919\ : std_logic;
signal \N__33918\ : std_logic;
signal \N__33917\ : std_logic;
signal \N__33916\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33886\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33846\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33825\ : std_logic;
signal \N__33822\ : std_logic;
signal \N__33821\ : std_logic;
signal \N__33818\ : std_logic;
signal \N__33815\ : std_logic;
signal \N__33812\ : std_logic;
signal \N__33807\ : std_logic;
signal \N__33804\ : std_logic;
signal \N__33801\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33783\ : std_logic;
signal \N__33780\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33776\ : std_logic;
signal \N__33775\ : std_logic;
signal \N__33772\ : std_logic;
signal \N__33769\ : std_logic;
signal \N__33766\ : std_logic;
signal \N__33761\ : std_logic;
signal \N__33758\ : std_logic;
signal \N__33755\ : std_logic;
signal \N__33752\ : std_logic;
signal \N__33747\ : std_logic;
signal \N__33744\ : std_logic;
signal \N__33741\ : std_logic;
signal \N__33738\ : std_logic;
signal \N__33737\ : std_logic;
signal \N__33734\ : std_logic;
signal \N__33731\ : std_logic;
signal \N__33730\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33704\ : std_logic;
signal \N__33703\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33683\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33674\ : std_logic;
signal \N__33673\ : std_logic;
signal \N__33670\ : std_logic;
signal \N__33665\ : std_logic;
signal \N__33662\ : std_logic;
signal \N__33659\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33648\ : std_logic;
signal \N__33645\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33639\ : std_logic;
signal \N__33636\ : std_logic;
signal \N__33635\ : std_logic;
signal \N__33630\ : std_logic;
signal \N__33627\ : std_logic;
signal \N__33624\ : std_logic;
signal \N__33621\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33612\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33597\ : std_logic;
signal \N__33594\ : std_logic;
signal \N__33591\ : std_logic;
signal \N__33588\ : std_logic;
signal \N__33585\ : std_logic;
signal \N__33582\ : std_logic;
signal \N__33579\ : std_logic;
signal \N__33576\ : std_logic;
signal \N__33573\ : std_logic;
signal \N__33570\ : std_logic;
signal \N__33567\ : std_logic;
signal \N__33564\ : std_logic;
signal \N__33561\ : std_logic;
signal \N__33558\ : std_logic;
signal \N__33557\ : std_logic;
signal \N__33556\ : std_logic;
signal \N__33553\ : std_logic;
signal \N__33550\ : std_logic;
signal \N__33547\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33537\ : std_logic;
signal \N__33534\ : std_logic;
signal \N__33531\ : std_logic;
signal \N__33528\ : std_logic;
signal \N__33525\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33515\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33501\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33486\ : std_logic;
signal \N__33483\ : std_logic;
signal \N__33480\ : std_logic;
signal \N__33479\ : std_logic;
signal \N__33476\ : std_logic;
signal \N__33473\ : std_logic;
signal \N__33470\ : std_logic;
signal \N__33465\ : std_logic;
signal \N__33462\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33450\ : std_logic;
signal \N__33447\ : std_logic;
signal \N__33444\ : std_logic;
signal \N__33441\ : std_logic;
signal \N__33438\ : std_logic;
signal \N__33435\ : std_logic;
signal \N__33432\ : std_logic;
signal \N__33431\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33425\ : std_logic;
signal \N__33422\ : std_logic;
signal \N__33419\ : std_logic;
signal \N__33416\ : std_logic;
signal \N__33413\ : std_logic;
signal \N__33408\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33399\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33393\ : std_logic;
signal \N__33390\ : std_logic;
signal \N__33387\ : std_logic;
signal \N__33384\ : std_logic;
signal \N__33381\ : std_logic;
signal \N__33378\ : std_logic;
signal \N__33375\ : std_logic;
signal \N__33372\ : std_logic;
signal \N__33369\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33362\ : std_logic;
signal \N__33359\ : std_logic;
signal \N__33356\ : std_logic;
signal \N__33353\ : std_logic;
signal \N__33350\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33342\ : std_logic;
signal \N__33339\ : std_logic;
signal \N__33336\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33327\ : std_logic;
signal \N__33324\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33318\ : std_logic;
signal \N__33315\ : std_logic;
signal \N__33312\ : std_logic;
signal \N__33309\ : std_logic;
signal \N__33306\ : std_logic;
signal \N__33303\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33279\ : std_logic;
signal \N__33276\ : std_logic;
signal \N__33273\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33258\ : std_logic;
signal \N__33255\ : std_logic;
signal \N__33252\ : std_logic;
signal \N__33249\ : std_logic;
signal \N__33246\ : std_logic;
signal \N__33243\ : std_logic;
signal \N__33240\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33228\ : std_logic;
signal \N__33225\ : std_logic;
signal \N__33222\ : std_logic;
signal \N__33219\ : std_logic;
signal \N__33216\ : std_logic;
signal \N__33213\ : std_logic;
signal \N__33210\ : std_logic;
signal \N__33207\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33198\ : std_logic;
signal \N__33195\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33186\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33174\ : std_logic;
signal \N__33171\ : std_logic;
signal \N__33168\ : std_logic;
signal \N__33165\ : std_logic;
signal \N__33162\ : std_logic;
signal \N__33159\ : std_logic;
signal \N__33156\ : std_logic;
signal \N__33153\ : std_logic;
signal \N__33150\ : std_logic;
signal \N__33147\ : std_logic;
signal \N__33144\ : std_logic;
signal \N__33141\ : std_logic;
signal \N__33138\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33132\ : std_logic;
signal \N__33129\ : std_logic;
signal \N__33126\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33120\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33102\ : std_logic;
signal \N__33099\ : std_logic;
signal \N__33096\ : std_logic;
signal \N__33093\ : std_logic;
signal \N__33090\ : std_logic;
signal \N__33087\ : std_logic;
signal \N__33084\ : std_logic;
signal \N__33081\ : std_logic;
signal \N__33078\ : std_logic;
signal \N__33075\ : std_logic;
signal \N__33072\ : std_logic;
signal \N__33069\ : std_logic;
signal \N__33066\ : std_logic;
signal \N__33063\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33057\ : std_logic;
signal \N__33054\ : std_logic;
signal \N__33051\ : std_logic;
signal \N__33048\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33036\ : std_logic;
signal \N__33033\ : std_logic;
signal \N__33030\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33021\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32997\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32993\ : std_logic;
signal \N__32992\ : std_logic;
signal \N__32989\ : std_logic;
signal \N__32986\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32982\ : std_logic;
signal \N__32977\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32970\ : std_logic;
signal \N__32967\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32952\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32950\ : std_logic;
signal \N__32949\ : std_logic;
signal \N__32946\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32919\ : std_logic;
signal \N__32916\ : std_logic;
signal \N__32913\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32900\ : std_logic;
signal \N__32899\ : std_logic;
signal \N__32896\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32883\ : std_logic;
signal \N__32878\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32872\ : std_logic;
signal \N__32865\ : std_logic;
signal \N__32862\ : std_logic;
signal \N__32859\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32856\ : std_logic;
signal \N__32855\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32838\ : std_logic;
signal \N__32835\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32826\ : std_logic;
signal \N__32825\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32814\ : std_logic;
signal \N__32811\ : std_logic;
signal \N__32806\ : std_logic;
signal \N__32799\ : std_logic;
signal \N__32796\ : std_logic;
signal \N__32793\ : std_logic;
signal \N__32790\ : std_logic;
signal \N__32787\ : std_logic;
signal \N__32784\ : std_logic;
signal \N__32783\ : std_logic;
signal \N__32782\ : std_logic;
signal \N__32777\ : std_logic;
signal \N__32774\ : std_logic;
signal \N__32771\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32764\ : std_logic;
signal \N__32761\ : std_logic;
signal \N__32758\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32750\ : std_logic;
signal \N__32745\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32743\ : std_logic;
signal \N__32740\ : std_logic;
signal \N__32733\ : std_logic;
signal \N__32730\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32724\ : std_logic;
signal \N__32721\ : std_logic;
signal \N__32718\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32712\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32706\ : std_logic;
signal \N__32703\ : std_logic;
signal \N__32702\ : std_logic;
signal \N__32699\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32697\ : std_logic;
signal \N__32696\ : std_logic;
signal \N__32693\ : std_logic;
signal \N__32688\ : std_logic;
signal \N__32685\ : std_logic;
signal \N__32682\ : std_logic;
signal \N__32673\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32671\ : std_logic;
signal \N__32668\ : std_logic;
signal \N__32667\ : std_logic;
signal \N__32666\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32658\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32646\ : std_logic;
signal \N__32643\ : std_logic;
signal \N__32640\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32636\ : std_logic;
signal \N__32635\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32633\ : std_logic;
signal \N__32632\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32621\ : std_logic;
signal \N__32618\ : std_logic;
signal \N__32613\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32602\ : std_logic;
signal \N__32599\ : std_logic;
signal \N__32596\ : std_logic;
signal \N__32593\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32591\ : std_logic;
signal \N__32588\ : std_logic;
signal \N__32585\ : std_logic;
signal \N__32582\ : std_logic;
signal \N__32577\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32567\ : std_logic;
signal \N__32566\ : std_logic;
signal \N__32561\ : std_logic;
signal \N__32558\ : std_logic;
signal \N__32557\ : std_logic;
signal \N__32552\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32541\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32539\ : std_logic;
signal \N__32538\ : std_logic;
signal \N__32529\ : std_logic;
signal \N__32526\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32517\ : std_logic;
signal \N__32516\ : std_logic;
signal \N__32513\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32506\ : std_logic;
signal \N__32503\ : std_logic;
signal \N__32500\ : std_logic;
signal \N__32497\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32490\ : std_logic;
signal \N__32489\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32485\ : std_logic;
signal \N__32482\ : std_logic;
signal \N__32479\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32473\ : std_logic;
signal \N__32470\ : std_logic;
signal \N__32465\ : std_logic;
signal \N__32462\ : std_logic;
signal \N__32451\ : std_logic;
signal \N__32448\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32433\ : std_logic;
signal \N__32430\ : std_logic;
signal \N__32427\ : std_logic;
signal \N__32424\ : std_logic;
signal \N__32421\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32412\ : std_logic;
signal \N__32409\ : std_logic;
signal \N__32406\ : std_logic;
signal \N__32403\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32397\ : std_logic;
signal \N__32394\ : std_logic;
signal \N__32391\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32385\ : std_logic;
signal \N__32382\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32376\ : std_logic;
signal \N__32373\ : std_logic;
signal \N__32370\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32363\ : std_logic;
signal \N__32362\ : std_logic;
signal \N__32361\ : std_logic;
signal \N__32360\ : std_logic;
signal \N__32357\ : std_logic;
signal \N__32350\ : std_logic;
signal \N__32347\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32337\ : std_logic;
signal \N__32336\ : std_logic;
signal \N__32331\ : std_logic;
signal \N__32328\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32313\ : std_logic;
signal \N__32312\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32306\ : std_logic;
signal \N__32303\ : std_logic;
signal \N__32298\ : std_logic;
signal \N__32297\ : std_logic;
signal \N__32294\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32280\ : std_logic;
signal \N__32277\ : std_logic;
signal \N__32276\ : std_logic;
signal \N__32273\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32271\ : std_logic;
signal \N__32268\ : std_logic;
signal \N__32265\ : std_logic;
signal \N__32260\ : std_logic;
signal \N__32257\ : std_logic;
signal \N__32250\ : std_logic;
signal \N__32247\ : std_logic;
signal \N__32244\ : std_logic;
signal \N__32241\ : std_logic;
signal \N__32238\ : std_logic;
signal \N__32235\ : std_logic;
signal \N__32232\ : std_logic;
signal \N__32229\ : std_logic;
signal \N__32226\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32222\ : std_logic;
signal \N__32219\ : std_logic;
signal \N__32216\ : std_logic;
signal \N__32213\ : std_logic;
signal \N__32208\ : std_logic;
signal \N__32207\ : std_logic;
signal \N__32204\ : std_logic;
signal \N__32201\ : std_logic;
signal \N__32198\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32188\ : std_logic;
signal \N__32185\ : std_logic;
signal \N__32182\ : std_logic;
signal \N__32177\ : std_logic;
signal \N__32172\ : std_logic;
signal \N__32171\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32167\ : std_logic;
signal \N__32164\ : std_logic;
signal \N__32161\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32149\ : std_logic;
signal \N__32142\ : std_logic;
signal \N__32139\ : std_logic;
signal \N__32136\ : std_logic;
signal \N__32133\ : std_logic;
signal \N__32130\ : std_logic;
signal \N__32127\ : std_logic;
signal \N__32124\ : std_logic;
signal \N__32123\ : std_logic;
signal \N__32120\ : std_logic;
signal \N__32117\ : std_logic;
signal \N__32114\ : std_logic;
signal \N__32111\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32105\ : std_logic;
signal \N__32102\ : std_logic;
signal \N__32097\ : std_logic;
signal \N__32094\ : std_logic;
signal \N__32091\ : std_logic;
signal \N__32088\ : std_logic;
signal \N__32085\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32072\ : std_logic;
signal \N__32067\ : std_logic;
signal \N__32064\ : std_logic;
signal \N__32061\ : std_logic;
signal \N__32058\ : std_logic;
signal \N__32057\ : std_logic;
signal \N__32052\ : std_logic;
signal \N__32049\ : std_logic;
signal \N__32046\ : std_logic;
signal \N__32043\ : std_logic;
signal \N__32040\ : std_logic;
signal \N__32039\ : std_logic;
signal \N__32036\ : std_logic;
signal \N__32031\ : std_logic;
signal \N__32028\ : std_logic;
signal \N__32025\ : std_logic;
signal \N__32022\ : std_logic;
signal \N__32019\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32013\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32007\ : std_logic;
signal \N__32004\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31981\ : std_logic;
signal \N__31978\ : std_logic;
signal \N__31975\ : std_logic;
signal \N__31972\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31962\ : std_logic;
signal \N__31959\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31953\ : std_logic;
signal \N__31950\ : std_logic;
signal \N__31947\ : std_logic;
signal \N__31944\ : std_logic;
signal \N__31941\ : std_logic;
signal \N__31938\ : std_logic;
signal \N__31935\ : std_logic;
signal \N__31932\ : std_logic;
signal \N__31929\ : std_logic;
signal \N__31926\ : std_logic;
signal \N__31923\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31914\ : std_logic;
signal \N__31911\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31899\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31890\ : std_logic;
signal \N__31887\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31881\ : std_logic;
signal \N__31878\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31863\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31854\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31842\ : std_logic;
signal \N__31839\ : std_logic;
signal \N__31836\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31815\ : std_logic;
signal \N__31812\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31803\ : std_logic;
signal \N__31800\ : std_logic;
signal \N__31797\ : std_logic;
signal \N__31794\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31785\ : std_logic;
signal \N__31782\ : std_logic;
signal \N__31779\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31773\ : std_logic;
signal \N__31770\ : std_logic;
signal \N__31767\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31761\ : std_logic;
signal \N__31758\ : std_logic;
signal \N__31755\ : std_logic;
signal \N__31752\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31746\ : std_logic;
signal \N__31743\ : std_logic;
signal \N__31740\ : std_logic;
signal \N__31737\ : std_logic;
signal \N__31734\ : std_logic;
signal \N__31731\ : std_logic;
signal \N__31728\ : std_logic;
signal \N__31725\ : std_logic;
signal \N__31722\ : std_logic;
signal \N__31719\ : std_logic;
signal \N__31716\ : std_logic;
signal \N__31713\ : std_logic;
signal \N__31710\ : std_logic;
signal \N__31707\ : std_logic;
signal \N__31704\ : std_logic;
signal \N__31701\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31689\ : std_logic;
signal \N__31686\ : std_logic;
signal \N__31683\ : std_logic;
signal \N__31680\ : std_logic;
signal \N__31677\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31671\ : std_logic;
signal \N__31668\ : std_logic;
signal \N__31665\ : std_logic;
signal \N__31662\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31650\ : std_logic;
signal \N__31647\ : std_logic;
signal \N__31644\ : std_logic;
signal \N__31641\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31623\ : std_logic;
signal \N__31620\ : std_logic;
signal \N__31617\ : std_logic;
signal \N__31614\ : std_logic;
signal \N__31611\ : std_logic;
signal \N__31608\ : std_logic;
signal \N__31605\ : std_logic;
signal \N__31602\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31590\ : std_logic;
signal \N__31589\ : std_logic;
signal \N__31586\ : std_logic;
signal \N__31583\ : std_logic;
signal \N__31580\ : std_logic;
signal \N__31575\ : std_logic;
signal \N__31572\ : std_logic;
signal \N__31569\ : std_logic;
signal \N__31566\ : std_logic;
signal \N__31563\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31557\ : std_logic;
signal \N__31554\ : std_logic;
signal \N__31551\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31545\ : std_logic;
signal \N__31542\ : std_logic;
signal \N__31539\ : std_logic;
signal \N__31536\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31530\ : std_logic;
signal \N__31527\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31518\ : std_logic;
signal \N__31515\ : std_logic;
signal \N__31512\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31503\ : std_logic;
signal \N__31500\ : std_logic;
signal \N__31497\ : std_logic;
signal \N__31494\ : std_logic;
signal \N__31491\ : std_logic;
signal \N__31488\ : std_logic;
signal \N__31487\ : std_logic;
signal \N__31482\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31477\ : std_logic;
signal \N__31474\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31468\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31458\ : std_logic;
signal \N__31457\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31451\ : std_logic;
signal \N__31448\ : std_logic;
signal \N__31445\ : std_logic;
signal \N__31442\ : std_logic;
signal \N__31439\ : std_logic;
signal \N__31436\ : std_logic;
signal \N__31433\ : std_logic;
signal \N__31430\ : std_logic;
signal \N__31427\ : std_logic;
signal \N__31418\ : std_logic;
signal \N__31413\ : std_logic;
signal \N__31410\ : std_logic;
signal \N__31407\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31395\ : std_logic;
signal \N__31392\ : std_logic;
signal \N__31389\ : std_logic;
signal \N__31386\ : std_logic;
signal \N__31385\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31383\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31372\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31340\ : std_logic;
signal \N__31337\ : std_logic;
signal \N__31336\ : std_logic;
signal \N__31333\ : std_logic;
signal \N__31330\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31317\ : std_logic;
signal \N__31314\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31308\ : std_logic;
signal \N__31305\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31301\ : std_logic;
signal \N__31298\ : std_logic;
signal \N__31293\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31282\ : std_logic;
signal \N__31281\ : std_logic;
signal \N__31280\ : std_logic;
signal \N__31275\ : std_logic;
signal \N__31268\ : std_logic;
signal \N__31263\ : std_logic;
signal \N__31262\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31260\ : std_logic;
signal \N__31259\ : std_logic;
signal \N__31258\ : std_logic;
signal \N__31257\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31255\ : std_logic;
signal \N__31248\ : std_logic;
signal \N__31241\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31227\ : std_logic;
signal \N__31226\ : std_logic;
signal \N__31225\ : std_logic;
signal \N__31222\ : std_logic;
signal \N__31219\ : std_logic;
signal \N__31218\ : std_logic;
signal \N__31215\ : std_logic;
signal \N__31208\ : std_logic;
signal \N__31203\ : std_logic;
signal \N__31200\ : std_logic;
signal \N__31197\ : std_logic;
signal \N__31194\ : std_logic;
signal \N__31191\ : std_logic;
signal \N__31188\ : std_logic;
signal \N__31185\ : std_logic;
signal \N__31184\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31172\ : std_logic;
signal \N__31171\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31163\ : std_logic;
signal \N__31162\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31160\ : std_logic;
signal \N__31157\ : std_logic;
signal \N__31154\ : std_logic;
signal \N__31147\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31139\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31128\ : std_logic;
signal \N__31125\ : std_logic;
signal \N__31124\ : std_logic;
signal \N__31123\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31119\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31113\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31101\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31092\ : std_logic;
signal \N__31091\ : std_logic;
signal \N__31090\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31078\ : std_logic;
signal \N__31071\ : std_logic;
signal \N__31068\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31044\ : std_logic;
signal \N__31041\ : std_logic;
signal \N__31038\ : std_logic;
signal \N__31035\ : std_logic;
signal \N__31032\ : std_logic;
signal \N__31029\ : std_logic;
signal \N__31028\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31026\ : std_logic;
signal \N__31023\ : std_logic;
signal \N__31020\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31014\ : std_logic;
signal \N__31005\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__30999\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30989\ : std_logic;
signal \N__30986\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30978\ : std_logic;
signal \N__30975\ : std_logic;
signal \N__30972\ : std_logic;
signal \N__30969\ : std_logic;
signal \N__30966\ : std_logic;
signal \N__30963\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30939\ : std_logic;
signal \N__30936\ : std_logic;
signal \N__30933\ : std_logic;
signal \N__30930\ : std_logic;
signal \N__30927\ : std_logic;
signal \N__30924\ : std_logic;
signal \N__30921\ : std_logic;
signal \N__30918\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30912\ : std_logic;
signal \N__30909\ : std_logic;
signal \N__30906\ : std_logic;
signal \N__30905\ : std_logic;
signal \N__30902\ : std_logic;
signal \N__30899\ : std_logic;
signal \N__30896\ : std_logic;
signal \N__30891\ : std_logic;
signal \N__30888\ : std_logic;
signal \N__30885\ : std_logic;
signal \N__30882\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30867\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30863\ : std_logic;
signal \N__30860\ : std_logic;
signal \N__30857\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30846\ : std_logic;
signal \N__30843\ : std_logic;
signal \N__30840\ : std_logic;
signal \N__30837\ : std_logic;
signal \N__30834\ : std_logic;
signal \N__30831\ : std_logic;
signal \N__30828\ : std_logic;
signal \N__30825\ : std_logic;
signal \N__30822\ : std_logic;
signal \N__30819\ : std_logic;
signal \N__30816\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30804\ : std_logic;
signal \N__30801\ : std_logic;
signal \N__30798\ : std_logic;
signal \N__30795\ : std_logic;
signal \N__30792\ : std_logic;
signal \N__30789\ : std_logic;
signal \N__30786\ : std_logic;
signal \N__30783\ : std_logic;
signal \N__30780\ : std_logic;
signal \N__30777\ : std_logic;
signal \N__30774\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30762\ : std_logic;
signal \N__30759\ : std_logic;
signal \N__30756\ : std_logic;
signal \N__30753\ : std_logic;
signal \N__30750\ : std_logic;
signal \N__30747\ : std_logic;
signal \N__30744\ : std_logic;
signal \N__30741\ : std_logic;
signal \N__30738\ : std_logic;
signal \N__30735\ : std_logic;
signal \N__30732\ : std_logic;
signal \N__30729\ : std_logic;
signal \N__30726\ : std_logic;
signal \N__30723\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30714\ : std_logic;
signal \N__30711\ : std_logic;
signal \N__30708\ : std_logic;
signal \N__30705\ : std_logic;
signal \N__30702\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30696\ : std_logic;
signal \N__30693\ : std_logic;
signal \N__30690\ : std_logic;
signal \N__30687\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30681\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30675\ : std_logic;
signal \N__30672\ : std_logic;
signal \N__30669\ : std_logic;
signal \N__30666\ : std_logic;
signal \N__30663\ : std_logic;
signal \N__30660\ : std_logic;
signal \N__30657\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30651\ : std_logic;
signal \N__30648\ : std_logic;
signal \N__30645\ : std_logic;
signal \N__30642\ : std_logic;
signal \N__30639\ : std_logic;
signal \N__30636\ : std_logic;
signal \N__30633\ : std_logic;
signal \N__30630\ : std_logic;
signal \N__30627\ : std_logic;
signal \N__30624\ : std_logic;
signal \N__30621\ : std_logic;
signal \N__30618\ : std_logic;
signal \N__30615\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30609\ : std_logic;
signal \N__30608\ : std_logic;
signal \N__30603\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30595\ : std_logic;
signal \N__30592\ : std_logic;
signal \N__30589\ : std_logic;
signal \N__30584\ : std_logic;
signal \N__30581\ : std_logic;
signal \N__30576\ : std_logic;
signal \N__30573\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30567\ : std_logic;
signal \N__30564\ : std_logic;
signal \N__30561\ : std_logic;
signal \N__30558\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30554\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30542\ : std_logic;
signal \N__30537\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30531\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30525\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30519\ : std_logic;
signal \N__30516\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30514\ : std_logic;
signal \N__30513\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30507\ : std_logic;
signal \N__30504\ : std_logic;
signal \N__30501\ : std_logic;
signal \N__30498\ : std_logic;
signal \N__30495\ : std_logic;
signal \N__30492\ : std_logic;
signal \N__30489\ : std_logic;
signal \N__30484\ : std_logic;
signal \N__30477\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30474\ : std_logic;
signal \N__30473\ : std_logic;
signal \N__30472\ : std_logic;
signal \N__30471\ : std_logic;
signal \N__30464\ : std_logic;
signal \N__30463\ : std_logic;
signal \N__30462\ : std_logic;
signal \N__30461\ : std_logic;
signal \N__30460\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30458\ : std_logic;
signal \N__30455\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30449\ : std_logic;
signal \N__30446\ : std_logic;
signal \N__30443\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30421\ : std_logic;
signal \N__30418\ : std_logic;
signal \N__30413\ : std_logic;
signal \N__30410\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30402\ : std_logic;
signal \N__30397\ : std_logic;
signal \N__30394\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30379\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30363\ : std_logic;
signal \N__30360\ : std_logic;
signal \N__30357\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30351\ : std_logic;
signal \N__30350\ : std_logic;
signal \N__30349\ : std_logic;
signal \N__30346\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30336\ : std_logic;
signal \N__30335\ : std_logic;
signal \N__30332\ : std_logic;
signal \N__30329\ : std_logic;
signal \N__30324\ : std_logic;
signal \N__30323\ : std_logic;
signal \N__30320\ : std_logic;
signal \N__30317\ : std_logic;
signal \N__30312\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30300\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30293\ : std_logic;
signal \N__30288\ : std_logic;
signal \N__30285\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30281\ : std_logic;
signal \N__30278\ : std_logic;
signal \N__30273\ : std_logic;
signal \N__30270\ : std_logic;
signal \N__30267\ : std_logic;
signal \N__30264\ : std_logic;
signal \N__30261\ : std_logic;
signal \N__30260\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30256\ : std_logic;
signal \N__30251\ : std_logic;
signal \N__30246\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30242\ : std_logic;
signal \N__30239\ : std_logic;
signal \N__30238\ : std_logic;
signal \N__30235\ : std_logic;
signal \N__30232\ : std_logic;
signal \N__30229\ : std_logic;
signal \N__30226\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30216\ : std_logic;
signal \N__30213\ : std_logic;
signal \N__30210\ : std_logic;
signal \N__30207\ : std_logic;
signal \N__30204\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30202\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30189\ : std_logic;
signal \N__30186\ : std_logic;
signal \N__30183\ : std_logic;
signal \N__30180\ : std_logic;
signal \N__30177\ : std_logic;
signal \N__30174\ : std_logic;
signal \N__30171\ : std_logic;
signal \N__30168\ : std_logic;
signal \N__30165\ : std_logic;
signal \N__30162\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30156\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30141\ : std_logic;
signal \N__30138\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30122\ : std_logic;
signal \N__30121\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30112\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30106\ : std_logic;
signal \N__30099\ : std_logic;
signal \N__30096\ : std_logic;
signal \N__30093\ : std_logic;
signal \N__30090\ : std_logic;
signal \N__30087\ : std_logic;
signal \N__30084\ : std_logic;
signal \N__30083\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30081\ : std_logic;
signal \N__30078\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30071\ : std_logic;
signal \N__30068\ : std_logic;
signal \N__30063\ : std_logic;
signal \N__30054\ : std_logic;
signal \N__30053\ : std_logic;
signal \N__30052\ : std_logic;
signal \N__30049\ : std_logic;
signal \N__30046\ : std_logic;
signal \N__30041\ : std_logic;
signal \N__30036\ : std_logic;
signal \N__30035\ : std_logic;
signal \N__30034\ : std_logic;
signal \N__30033\ : std_logic;
signal \N__30030\ : std_logic;
signal \N__30027\ : std_logic;
signal \N__30026\ : std_logic;
signal \N__30023\ : std_logic;
signal \N__30020\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30012\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29996\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29988\ : std_logic;
signal \N__29987\ : std_logic;
signal \N__29986\ : std_logic;
signal \N__29983\ : std_logic;
signal \N__29976\ : std_logic;
signal \N__29973\ : std_logic;
signal \N__29970\ : std_logic;
signal \N__29969\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29962\ : std_logic;
signal \N__29959\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29957\ : std_logic;
signal \N__29952\ : std_logic;
signal \N__29951\ : std_logic;
signal \N__29950\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29942\ : std_logic;
signal \N__29941\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29932\ : std_logic;
signal \N__29929\ : std_logic;
signal \N__29924\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29920\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29910\ : std_logic;
signal \N__29905\ : std_logic;
signal \N__29900\ : std_logic;
signal \N__29895\ : std_logic;
signal \N__29892\ : std_logic;
signal \N__29889\ : std_logic;
signal \N__29888\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29877\ : std_logic;
signal \N__29874\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29862\ : std_logic;
signal \N__29859\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29855\ : std_logic;
signal \N__29852\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29841\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29820\ : std_logic;
signal \N__29817\ : std_logic;
signal \N__29814\ : std_logic;
signal \N__29811\ : std_logic;
signal \N__29808\ : std_logic;
signal \N__29805\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29790\ : std_logic;
signal \N__29787\ : std_logic;
signal \N__29784\ : std_logic;
signal \N__29781\ : std_logic;
signal \N__29778\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29769\ : std_logic;
signal \N__29766\ : std_logic;
signal \N__29763\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29757\ : std_logic;
signal \N__29754\ : std_logic;
signal \N__29751\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29742\ : std_logic;
signal \N__29739\ : std_logic;
signal \N__29736\ : std_logic;
signal \N__29733\ : std_logic;
signal \N__29730\ : std_logic;
signal \N__29727\ : std_logic;
signal \N__29724\ : std_logic;
signal \N__29721\ : std_logic;
signal \N__29718\ : std_logic;
signal \N__29715\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29709\ : std_logic;
signal \N__29706\ : std_logic;
signal \N__29703\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29697\ : std_logic;
signal \N__29694\ : std_logic;
signal \N__29691\ : std_logic;
signal \N__29690\ : std_logic;
signal \N__29689\ : std_logic;
signal \N__29686\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29670\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29664\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29658\ : std_logic;
signal \N__29655\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29646\ : std_logic;
signal \N__29643\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29637\ : std_logic;
signal \N__29634\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29625\ : std_logic;
signal \N__29622\ : std_logic;
signal \N__29619\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29601\ : std_logic;
signal \N__29598\ : std_logic;
signal \N__29595\ : std_logic;
signal \N__29592\ : std_logic;
signal \N__29589\ : std_logic;
signal \N__29586\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29577\ : std_logic;
signal \N__29574\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29565\ : std_logic;
signal \N__29562\ : std_logic;
signal \N__29559\ : std_logic;
signal \N__29556\ : std_logic;
signal \N__29553\ : std_logic;
signal \N__29550\ : std_logic;
signal \N__29547\ : std_logic;
signal \N__29544\ : std_logic;
signal \N__29541\ : std_logic;
signal \N__29538\ : std_logic;
signal \N__29535\ : std_logic;
signal \N__29532\ : std_logic;
signal \N__29529\ : std_logic;
signal \N__29526\ : std_logic;
signal \N__29523\ : std_logic;
signal \N__29520\ : std_logic;
signal \N__29517\ : std_logic;
signal \N__29514\ : std_logic;
signal \N__29511\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29505\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29487\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29481\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29463\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29451\ : std_logic;
signal \N__29448\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29436\ : std_logic;
signal \N__29433\ : std_logic;
signal \N__29430\ : std_logic;
signal \N__29427\ : std_logic;
signal \N__29424\ : std_logic;
signal \N__29421\ : std_logic;
signal \N__29418\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29412\ : std_logic;
signal \N__29409\ : std_logic;
signal \N__29406\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29399\ : std_logic;
signal \N__29394\ : std_logic;
signal \N__29393\ : std_logic;
signal \N__29392\ : std_logic;
signal \N__29391\ : std_logic;
signal \N__29390\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29374\ : std_logic;
signal \N__29367\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29365\ : std_logic;
signal \N__29364\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29353\ : std_logic;
signal \N__29350\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29340\ : std_logic;
signal \N__29337\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29325\ : std_logic;
signal \N__29322\ : std_logic;
signal \N__29319\ : std_logic;
signal \N__29316\ : std_logic;
signal \N__29313\ : std_logic;
signal \N__29310\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29301\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29283\ : std_logic;
signal \N__29280\ : std_logic;
signal \N__29277\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29271\ : std_logic;
signal \N__29268\ : std_logic;
signal \N__29265\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29259\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29247\ : std_logic;
signal \N__29244\ : std_logic;
signal \N__29241\ : std_logic;
signal \N__29238\ : std_logic;
signal \N__29235\ : std_logic;
signal \N__29234\ : std_logic;
signal \N__29229\ : std_logic;
signal \N__29226\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29223\ : std_logic;
signal \N__29222\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29220\ : std_logic;
signal \N__29219\ : std_logic;
signal \N__29216\ : std_logic;
signal \N__29209\ : std_logic;
signal \N__29204\ : std_logic;
signal \N__29199\ : std_logic;
signal \N__29190\ : std_logic;
signal \N__29189\ : std_logic;
signal \N__29186\ : std_logic;
signal \N__29183\ : std_logic;
signal \N__29178\ : std_logic;
signal \N__29177\ : std_logic;
signal \N__29172\ : std_logic;
signal \N__29169\ : std_logic;
signal \N__29168\ : std_logic;
signal \N__29167\ : std_logic;
signal \N__29166\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29148\ : std_logic;
signal \N__29147\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29135\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29126\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29118\ : std_logic;
signal \N__29117\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29106\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29100\ : std_logic;
signal \N__29099\ : std_logic;
signal \N__29096\ : std_logic;
signal \N__29095\ : std_logic;
signal \N__29092\ : std_logic;
signal \N__29089\ : std_logic;
signal \N__29086\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29066\ : std_logic;
signal \N__29061\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29057\ : std_logic;
signal \N__29054\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29048\ : std_logic;
signal \N__29045\ : std_logic;
signal \N__29042\ : std_logic;
signal \N__29041\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29037\ : std_logic;
signal \N__29034\ : std_logic;
signal \N__29033\ : std_logic;
signal \N__29030\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29024\ : std_logic;
signal \N__29021\ : std_logic;
signal \N__29016\ : std_logic;
signal \N__29007\ : std_logic;
signal \N__29006\ : std_logic;
signal \N__29003\ : std_logic;
signal \N__29000\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28995\ : std_logic;
signal \N__28992\ : std_logic;
signal \N__28989\ : std_logic;
signal \N__28986\ : std_logic;
signal \N__28983\ : std_logic;
signal \N__28980\ : std_logic;
signal \N__28977\ : std_logic;
signal \N__28974\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28958\ : std_logic;
signal \N__28957\ : std_logic;
signal \N__28956\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28946\ : std_logic;
signal \N__28941\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28935\ : std_logic;
signal \N__28932\ : std_logic;
signal \N__28929\ : std_logic;
signal \N__28926\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28920\ : std_logic;
signal \N__28917\ : std_logic;
signal \N__28914\ : std_logic;
signal \N__28911\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28908\ : std_logic;
signal \N__28905\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28897\ : std_logic;
signal \N__28890\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28886\ : std_logic;
signal \N__28883\ : std_logic;
signal \N__28880\ : std_logic;
signal \N__28875\ : std_logic;
signal \N__28874\ : std_logic;
signal \N__28871\ : std_logic;
signal \N__28868\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28853\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28849\ : std_logic;
signal \N__28848\ : std_logic;
signal \N__28847\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28841\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28812\ : std_logic;
signal \N__28809\ : std_logic;
signal \N__28806\ : std_logic;
signal \N__28803\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28796\ : std_logic;
signal \N__28793\ : std_logic;
signal \N__28790\ : std_logic;
signal \N__28787\ : std_logic;
signal \N__28782\ : std_logic;
signal \N__28779\ : std_logic;
signal \N__28776\ : std_logic;
signal \N__28773\ : std_logic;
signal \N__28770\ : std_logic;
signal \N__28767\ : std_logic;
signal \N__28764\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28755\ : std_logic;
signal \N__28752\ : std_logic;
signal \N__28749\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28740\ : std_logic;
signal \N__28737\ : std_logic;
signal \N__28734\ : std_logic;
signal \N__28731\ : std_logic;
signal \N__28728\ : std_logic;
signal \N__28725\ : std_logic;
signal \N__28722\ : std_logic;
signal \N__28719\ : std_logic;
signal \N__28716\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28710\ : std_logic;
signal \N__28707\ : std_logic;
signal \N__28704\ : std_logic;
signal \N__28701\ : std_logic;
signal \N__28698\ : std_logic;
signal \N__28695\ : std_logic;
signal \N__28692\ : std_logic;
signal \N__28689\ : std_logic;
signal \N__28686\ : std_logic;
signal \N__28683\ : std_logic;
signal \N__28680\ : std_logic;
signal \N__28677\ : std_logic;
signal \N__28674\ : std_logic;
signal \N__28671\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28662\ : std_logic;
signal \N__28659\ : std_logic;
signal \N__28656\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28638\ : std_logic;
signal \N__28635\ : std_logic;
signal \N__28632\ : std_logic;
signal \N__28629\ : std_logic;
signal \N__28626\ : std_logic;
signal \N__28623\ : std_logic;
signal \N__28620\ : std_logic;
signal \N__28617\ : std_logic;
signal \N__28614\ : std_logic;
signal \N__28611\ : std_logic;
signal \N__28608\ : std_logic;
signal \N__28605\ : std_logic;
signal \N__28602\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28596\ : std_logic;
signal \N__28593\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28584\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28577\ : std_logic;
signal \N__28574\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28562\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28550\ : std_logic;
signal \N__28547\ : std_logic;
signal \N__28542\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28536\ : std_logic;
signal \N__28533\ : std_logic;
signal \N__28530\ : std_logic;
signal \N__28527\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28509\ : std_logic;
signal \N__28506\ : std_logic;
signal \N__28503\ : std_logic;
signal \N__28500\ : std_logic;
signal \N__28497\ : std_logic;
signal \N__28494\ : std_logic;
signal \N__28491\ : std_logic;
signal \N__28488\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28479\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28467\ : std_logic;
signal \N__28464\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28455\ : std_logic;
signal \N__28452\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28434\ : std_logic;
signal \N__28431\ : std_logic;
signal \N__28428\ : std_logic;
signal \N__28425\ : std_logic;
signal \N__28422\ : std_logic;
signal \N__28419\ : std_logic;
signal \N__28416\ : std_logic;
signal \N__28413\ : std_logic;
signal \N__28410\ : std_logic;
signal \N__28407\ : std_logic;
signal \N__28404\ : std_logic;
signal \N__28401\ : std_logic;
signal \N__28398\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28392\ : std_logic;
signal \N__28389\ : std_logic;
signal \N__28386\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28380\ : std_logic;
signal \N__28377\ : std_logic;
signal \N__28374\ : std_logic;
signal \N__28371\ : std_logic;
signal \N__28368\ : std_logic;
signal \N__28365\ : std_logic;
signal \N__28362\ : std_logic;
signal \N__28359\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28353\ : std_logic;
signal \N__28350\ : std_logic;
signal \N__28347\ : std_logic;
signal \N__28344\ : std_logic;
signal \N__28341\ : std_logic;
signal \N__28338\ : std_logic;
signal \N__28335\ : std_logic;
signal \N__28332\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28326\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28321\ : std_logic;
signal \N__28314\ : std_logic;
signal \N__28311\ : std_logic;
signal \N__28308\ : std_logic;
signal \N__28305\ : std_logic;
signal \N__28302\ : std_logic;
signal \N__28299\ : std_logic;
signal \N__28296\ : std_logic;
signal \N__28293\ : std_logic;
signal \N__28290\ : std_logic;
signal \N__28287\ : std_logic;
signal \N__28284\ : std_logic;
signal \N__28281\ : std_logic;
signal \N__28278\ : std_logic;
signal \N__28275\ : std_logic;
signal \N__28272\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28266\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28242\ : std_logic;
signal \N__28239\ : std_logic;
signal \N__28236\ : std_logic;
signal \N__28233\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28227\ : std_logic;
signal \N__28224\ : std_logic;
signal \N__28221\ : std_logic;
signal \N__28218\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28203\ : std_logic;
signal \N__28200\ : std_logic;
signal \N__28197\ : std_logic;
signal \N__28194\ : std_logic;
signal \N__28191\ : std_logic;
signal \N__28188\ : std_logic;
signal \N__28185\ : std_logic;
signal \N__28182\ : std_logic;
signal \N__28181\ : std_logic;
signal \N__28178\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28168\ : std_logic;
signal \N__28165\ : std_logic;
signal \N__28162\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28146\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28134\ : std_logic;
signal \N__28131\ : std_logic;
signal \N__28128\ : std_logic;
signal \N__28125\ : std_logic;
signal \N__28122\ : std_logic;
signal \N__28119\ : std_logic;
signal \N__28116\ : std_logic;
signal \N__28113\ : std_logic;
signal \N__28110\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28104\ : std_logic;
signal \N__28101\ : std_logic;
signal \N__28098\ : std_logic;
signal \N__28095\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28089\ : std_logic;
signal \N__28086\ : std_logic;
signal \N__28083\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28074\ : std_logic;
signal \N__28071\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28065\ : std_logic;
signal \N__28062\ : std_logic;
signal \N__28059\ : std_logic;
signal \N__28056\ : std_logic;
signal \N__28053\ : std_logic;
signal \N__28050\ : std_logic;
signal \N__28047\ : std_logic;
signal \N__28044\ : std_logic;
signal \N__28041\ : std_logic;
signal \N__28038\ : std_logic;
signal \N__28035\ : std_logic;
signal \N__28032\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28023\ : std_logic;
signal \N__28020\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28014\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27999\ : std_logic;
signal \N__27996\ : std_logic;
signal \N__27993\ : std_logic;
signal \N__27990\ : std_logic;
signal \N__27987\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27978\ : std_logic;
signal \N__27977\ : std_logic;
signal \N__27974\ : std_logic;
signal \N__27971\ : std_logic;
signal \N__27966\ : std_logic;
signal \N__27965\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27954\ : std_logic;
signal \N__27951\ : std_logic;
signal \N__27948\ : std_logic;
signal \N__27945\ : std_logic;
signal \N__27942\ : std_logic;
signal \N__27939\ : std_logic;
signal \N__27936\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27930\ : std_logic;
signal \N__27927\ : std_logic;
signal \N__27924\ : std_logic;
signal \N__27921\ : std_logic;
signal \N__27918\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27911\ : std_logic;
signal \N__27908\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27900\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27894\ : std_logic;
signal \N__27891\ : std_logic;
signal \N__27888\ : std_logic;
signal \N__27885\ : std_logic;
signal \N__27884\ : std_logic;
signal \N__27881\ : std_logic;
signal \N__27878\ : std_logic;
signal \N__27873\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27858\ : std_logic;
signal \N__27855\ : std_logic;
signal \N__27854\ : std_logic;
signal \N__27851\ : std_logic;
signal \N__27848\ : std_logic;
signal \N__27845\ : std_logic;
signal \N__27840\ : std_logic;
signal \N__27837\ : std_logic;
signal \N__27834\ : std_logic;
signal \N__27831\ : std_logic;
signal \N__27828\ : std_logic;
signal \N__27827\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27823\ : std_logic;
signal \N__27822\ : std_logic;
signal \N__27821\ : std_logic;
signal \N__27818\ : std_logic;
signal \N__27817\ : std_logic;
signal \N__27814\ : std_logic;
signal \N__27803\ : std_logic;
signal \N__27798\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27792\ : std_logic;
signal \N__27789\ : std_logic;
signal \N__27788\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27786\ : std_logic;
signal \N__27785\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27783\ : std_logic;
signal \N__27782\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27780\ : std_logic;
signal \N__27779\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27777\ : std_logic;
signal \N__27776\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27774\ : std_logic;
signal \N__27773\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27771\ : std_logic;
signal \N__27770\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27768\ : std_logic;
signal \N__27765\ : std_logic;
signal \N__27762\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27728\ : std_logic;
signal \N__27719\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27707\ : std_logic;
signal \N__27704\ : std_logic;
signal \N__27701\ : std_logic;
signal \N__27698\ : std_logic;
signal \N__27695\ : std_logic;
signal \N__27690\ : std_logic;
signal \N__27687\ : std_logic;
signal \N__27684\ : std_logic;
signal \N__27681\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27669\ : std_logic;
signal \N__27666\ : std_logic;
signal \N__27665\ : std_logic;
signal \N__27662\ : std_logic;
signal \N__27659\ : std_logic;
signal \N__27654\ : std_logic;
signal \N__27653\ : std_logic;
signal \N__27650\ : std_logic;
signal \N__27647\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27638\ : std_logic;
signal \N__27635\ : std_logic;
signal \N__27632\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27626\ : std_logic;
signal \N__27623\ : std_logic;
signal \N__27620\ : std_logic;
signal \N__27615\ : std_logic;
signal \N__27612\ : std_logic;
signal \N__27611\ : std_logic;
signal \N__27608\ : std_logic;
signal \N__27605\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27599\ : std_logic;
signal \N__27598\ : std_logic;
signal \N__27597\ : std_logic;
signal \N__27596\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27584\ : std_logic;
signal \N__27579\ : std_logic;
signal \N__27578\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27519\ : std_logic;
signal \N__27516\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27510\ : std_logic;
signal \N__27507\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27501\ : std_logic;
signal \N__27498\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27492\ : std_logic;
signal \N__27489\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27483\ : std_logic;
signal \N__27480\ : std_logic;
signal \N__27477\ : std_logic;
signal \N__27474\ : std_logic;
signal \N__27471\ : std_logic;
signal \N__27468\ : std_logic;
signal \N__27465\ : std_logic;
signal \N__27462\ : std_logic;
signal \N__27459\ : std_logic;
signal \N__27456\ : std_logic;
signal \N__27453\ : std_logic;
signal \N__27450\ : std_logic;
signal \N__27447\ : std_logic;
signal \N__27444\ : std_logic;
signal \N__27441\ : std_logic;
signal \N__27438\ : std_logic;
signal \N__27435\ : std_logic;
signal \N__27432\ : std_logic;
signal \N__27429\ : std_logic;
signal \N__27426\ : std_logic;
signal \N__27423\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27417\ : std_logic;
signal \N__27414\ : std_logic;
signal \N__27411\ : std_logic;
signal \N__27408\ : std_logic;
signal \N__27405\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27396\ : std_logic;
signal \N__27393\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27384\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27378\ : std_logic;
signal \N__27375\ : std_logic;
signal \N__27372\ : std_logic;
signal \N__27369\ : std_logic;
signal \N__27366\ : std_logic;
signal \N__27363\ : std_logic;
signal \N__27360\ : std_logic;
signal \N__27357\ : std_logic;
signal \N__27354\ : std_logic;
signal \N__27351\ : std_logic;
signal \N__27348\ : std_logic;
signal \N__27345\ : std_logic;
signal \N__27342\ : std_logic;
signal \N__27339\ : std_logic;
signal \N__27336\ : std_logic;
signal \N__27333\ : std_logic;
signal \N__27330\ : std_logic;
signal \N__27327\ : std_logic;
signal \N__27324\ : std_logic;
signal \N__27321\ : std_logic;
signal \N__27318\ : std_logic;
signal \N__27315\ : std_logic;
signal \N__27312\ : std_logic;
signal \N__27309\ : std_logic;
signal \N__27306\ : std_logic;
signal \N__27303\ : std_logic;
signal \N__27300\ : std_logic;
signal \N__27297\ : std_logic;
signal \N__27294\ : std_logic;
signal \N__27291\ : std_logic;
signal \N__27288\ : std_logic;
signal \N__27285\ : std_logic;
signal \N__27282\ : std_logic;
signal \N__27279\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27264\ : std_logic;
signal \N__27261\ : std_logic;
signal \N__27258\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27252\ : std_logic;
signal \N__27249\ : std_logic;
signal \N__27246\ : std_logic;
signal \N__27243\ : std_logic;
signal \N__27240\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27232\ : std_logic;
signal \N__27229\ : std_logic;
signal \N__27226\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27210\ : std_logic;
signal \N__27209\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27207\ : std_logic;
signal \N__27204\ : std_logic;
signal \N__27199\ : std_logic;
signal \N__27196\ : std_logic;
signal \N__27195\ : std_logic;
signal \N__27194\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27183\ : std_logic;
signal \N__27182\ : std_logic;
signal \N__27177\ : std_logic;
signal \N__27174\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27161\ : std_logic;
signal \N__27150\ : std_logic;
signal \N__27149\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27147\ : std_logic;
signal \N__27146\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27144\ : std_logic;
signal \N__27143\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27141\ : std_logic;
signal \N__27140\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27136\ : std_logic;
signal \N__27135\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27133\ : std_logic;
signal \N__27132\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27125\ : std_logic;
signal \N__27114\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27107\ : std_logic;
signal \N__27098\ : std_logic;
signal \N__27083\ : std_logic;
signal \N__27080\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27068\ : std_logic;
signal \N__27065\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27047\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27035\ : std_logic;
signal \N__27032\ : std_logic;
signal \N__27027\ : std_logic;
signal \N__27024\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27012\ : std_logic;
signal \N__27009\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26999\ : std_logic;
signal \N__26998\ : std_logic;
signal \N__26997\ : std_logic;
signal \N__26996\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26994\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26990\ : std_logic;
signal \N__26983\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26976\ : std_logic;
signal \N__26973\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26958\ : std_logic;
signal \N__26955\ : std_logic;
signal \N__26948\ : std_logic;
signal \N__26937\ : std_logic;
signal \N__26934\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26932\ : std_logic;
signal \N__26931\ : std_logic;
signal \N__26928\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26923\ : std_logic;
signal \N__26920\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26911\ : std_logic;
signal \N__26906\ : std_logic;
signal \N__26895\ : std_logic;
signal \N__26894\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26889\ : std_logic;
signal \N__26888\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26868\ : std_logic;
signal \N__26865\ : std_logic;
signal \N__26862\ : std_logic;
signal \N__26859\ : std_logic;
signal \N__26856\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26841\ : std_logic;
signal \N__26838\ : std_logic;
signal \N__26835\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26820\ : std_logic;
signal \N__26817\ : std_logic;
signal \N__26814\ : std_logic;
signal \N__26811\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26805\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26781\ : std_logic;
signal \N__26778\ : std_logic;
signal \N__26775\ : std_logic;
signal \N__26772\ : std_logic;
signal \N__26769\ : std_logic;
signal \N__26766\ : std_logic;
signal \N__26763\ : std_logic;
signal \N__26760\ : std_logic;
signal \N__26757\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26733\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26724\ : std_logic;
signal \N__26721\ : std_logic;
signal \N__26718\ : std_logic;
signal \N__26715\ : std_logic;
signal \N__26712\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26700\ : std_logic;
signal \N__26697\ : std_logic;
signal \N__26694\ : std_logic;
signal \N__26691\ : std_logic;
signal \N__26688\ : std_logic;
signal \N__26685\ : std_logic;
signal \N__26682\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26672\ : std_logic;
signal \N__26669\ : std_logic;
signal \N__26666\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26655\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26647\ : std_logic;
signal \N__26644\ : std_logic;
signal \N__26637\ : std_logic;
signal \N__26636\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26613\ : std_logic;
signal \N__26610\ : std_logic;
signal \N__26607\ : std_logic;
signal \N__26604\ : std_logic;
signal \N__26601\ : std_logic;
signal \N__26598\ : std_logic;
signal \N__26595\ : std_logic;
signal \N__26592\ : std_logic;
signal \N__26589\ : std_logic;
signal \N__26586\ : std_logic;
signal \N__26583\ : std_logic;
signal \N__26580\ : std_logic;
signal \N__26577\ : std_logic;
signal \N__26574\ : std_logic;
signal \N__26571\ : std_logic;
signal \N__26568\ : std_logic;
signal \N__26565\ : std_logic;
signal \N__26562\ : std_logic;
signal \N__26559\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26552\ : std_logic;
signal \N__26549\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26545\ : std_logic;
signal \N__26542\ : std_logic;
signal \N__26539\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26530\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26524\ : std_logic;
signal \N__26519\ : std_logic;
signal \N__26514\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26510\ : std_logic;
signal \N__26509\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26502\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26496\ : std_logic;
signal \N__26493\ : std_logic;
signal \N__26490\ : std_logic;
signal \N__26487\ : std_logic;
signal \N__26482\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26472\ : std_logic;
signal \N__26469\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26465\ : std_logic;
signal \N__26464\ : std_logic;
signal \N__26461\ : std_logic;
signal \N__26458\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26451\ : std_logic;
signal \N__26448\ : std_logic;
signal \N__26445\ : std_logic;
signal \N__26442\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26424\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26413\ : std_logic;
signal \N__26412\ : std_logic;
signal \N__26409\ : std_logic;
signal \N__26404\ : std_logic;
signal \N__26401\ : std_logic;
signal \N__26398\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26388\ : std_logic;
signal \N__26385\ : std_logic;
signal \N__26384\ : std_logic;
signal \N__26381\ : std_logic;
signal \N__26380\ : std_logic;
signal \N__26377\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26367\ : std_logic;
signal \N__26364\ : std_logic;
signal \N__26361\ : std_logic;
signal \N__26358\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26352\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26339\ : std_logic;
signal \N__26338\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26336\ : std_logic;
signal \N__26335\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26333\ : std_logic;
signal \N__26332\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26330\ : std_logic;
signal \N__26329\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26327\ : std_logic;
signal \N__26326\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26324\ : std_logic;
signal \N__26321\ : std_logic;
signal \N__26320\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26316\ : std_logic;
signal \N__26313\ : std_logic;
signal \N__26312\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26302\ : std_logic;
signal \N__26297\ : std_logic;
signal \N__26296\ : std_logic;
signal \N__26293\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26288\ : std_logic;
signal \N__26285\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26276\ : std_logic;
signal \N__26273\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26271\ : std_logic;
signal \N__26268\ : std_logic;
signal \N__26265\ : std_logic;
signal \N__26264\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26258\ : std_logic;
signal \N__26249\ : std_logic;
signal \N__26246\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26230\ : std_logic;
signal \N__26213\ : std_logic;
signal \N__26202\ : std_logic;
signal \N__26187\ : std_logic;
signal \N__26186\ : std_logic;
signal \N__26183\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26170\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26157\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26147\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26139\ : std_logic;
signal \N__26136\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26121\ : std_logic;
signal \N__26118\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26108\ : std_logic;
signal \N__26105\ : std_logic;
signal \N__26100\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26096\ : std_logic;
signal \N__26093\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26082\ : std_logic;
signal \N__26079\ : std_logic;
signal \N__26078\ : std_logic;
signal \N__26075\ : std_logic;
signal \N__26072\ : std_logic;
signal \N__26069\ : std_logic;
signal \N__26064\ : std_logic;
signal \N__26061\ : std_logic;
signal \N__26058\ : std_logic;
signal \N__26057\ : std_logic;
signal \N__26054\ : std_logic;
signal \N__26051\ : std_logic;
signal \N__26048\ : std_logic;
signal \N__26043\ : std_logic;
signal \N__26040\ : std_logic;
signal \N__26039\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26037\ : std_logic;
signal \N__26036\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26024\ : std_logic;
signal \N__26019\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26013\ : std_logic;
signal \N__26010\ : std_logic;
signal \N__26009\ : std_logic;
signal \N__26006\ : std_logic;
signal \N__26003\ : std_logic;
signal \N__26000\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25991\ : std_logic;
signal \N__25990\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25971\ : std_logic;
signal \N__25968\ : std_logic;
signal \N__25965\ : std_logic;
signal \N__25962\ : std_logic;
signal \N__25959\ : std_logic;
signal \N__25958\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25938\ : std_logic;
signal \N__25935\ : std_logic;
signal \N__25932\ : std_logic;
signal \N__25929\ : std_logic;
signal \N__25926\ : std_logic;
signal \N__25925\ : std_logic;
signal \N__25922\ : std_logic;
signal \N__25919\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25915\ : std_logic;
signal \N__25912\ : std_logic;
signal \N__25909\ : std_logic;
signal \N__25906\ : std_logic;
signal \N__25899\ : std_logic;
signal \N__25896\ : std_logic;
signal \N__25893\ : std_logic;
signal \N__25890\ : std_logic;
signal \N__25887\ : std_logic;
signal \N__25884\ : std_logic;
signal \N__25883\ : std_logic;
signal \N__25880\ : std_logic;
signal \N__25877\ : std_logic;
signal \N__25874\ : std_logic;
signal \N__25869\ : std_logic;
signal \N__25866\ : std_logic;
signal \N__25863\ : std_logic;
signal \N__25860\ : std_logic;
signal \N__25857\ : std_logic;
signal \N__25854\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25845\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25841\ : std_logic;
signal \N__25840\ : std_logic;
signal \N__25839\ : std_logic;
signal \N__25838\ : std_logic;
signal \N__25835\ : std_logic;
signal \N__25832\ : std_logic;
signal \N__25829\ : std_logic;
signal \N__25824\ : std_logic;
signal \N__25821\ : std_logic;
signal \N__25812\ : std_logic;
signal \N__25809\ : std_logic;
signal \N__25808\ : std_logic;
signal \N__25805\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25802\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25789\ : std_logic;
signal \N__25782\ : std_logic;
signal \N__25781\ : std_logic;
signal \N__25780\ : std_logic;
signal \N__25779\ : std_logic;
signal \N__25778\ : std_logic;
signal \N__25775\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25763\ : std_logic;
signal \N__25760\ : std_logic;
signal \N__25755\ : std_logic;
signal \N__25752\ : std_logic;
signal \N__25751\ : std_logic;
signal \N__25748\ : std_logic;
signal \N__25747\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25745\ : std_logic;
signal \N__25744\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25742\ : std_logic;
signal \N__25741\ : std_logic;
signal \N__25740\ : std_logic;
signal \N__25737\ : std_logic;
signal \N__25736\ : std_logic;
signal \N__25733\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25711\ : std_logic;
signal \N__25704\ : std_logic;
signal \N__25701\ : std_logic;
signal \N__25698\ : std_logic;
signal \N__25697\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25695\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25686\ : std_logic;
signal \N__25683\ : std_logic;
signal \N__25682\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25673\ : std_logic;
signal \N__25670\ : std_logic;
signal \N__25665\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25653\ : std_logic;
signal \N__25650\ : std_logic;
signal \N__25647\ : std_logic;
signal \N__25644\ : std_logic;
signal \N__25641\ : std_logic;
signal \N__25638\ : std_logic;
signal \N__25635\ : std_logic;
signal \N__25632\ : std_logic;
signal \N__25629\ : std_logic;
signal \N__25628\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25626\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25617\ : std_logic;
signal \N__25616\ : std_logic;
signal \N__25613\ : std_logic;
signal \N__25608\ : std_logic;
signal \N__25605\ : std_logic;
signal \N__25602\ : std_logic;
signal \N__25595\ : std_logic;
signal \N__25590\ : std_logic;
signal \N__25587\ : std_logic;
signal \N__25584\ : std_logic;
signal \N__25583\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25578\ : std_logic;
signal \N__25577\ : std_logic;
signal \N__25574\ : std_logic;
signal \N__25569\ : std_logic;
signal \N__25566\ : std_logic;
signal \N__25563\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25557\ : std_logic;
signal \N__25554\ : std_logic;
signal \N__25545\ : std_logic;
signal \N__25542\ : std_logic;
signal \N__25539\ : std_logic;
signal \N__25536\ : std_logic;
signal \N__25535\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25530\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25524\ : std_logic;
signal \N__25523\ : std_logic;
signal \N__25520\ : std_logic;
signal \N__25517\ : std_logic;
signal \N__25514\ : std_logic;
signal \N__25509\ : std_logic;
signal \N__25506\ : std_logic;
signal \N__25503\ : std_logic;
signal \N__25496\ : std_logic;
signal \N__25491\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25487\ : std_logic;
signal \N__25484\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25477\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25460\ : std_logic;
signal \N__25459\ : std_logic;
signal \N__25458\ : std_logic;
signal \N__25453\ : std_logic;
signal \N__25448\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25441\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25437\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25422\ : std_logic;
signal \N__25419\ : std_logic;
signal \N__25416\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25404\ : std_logic;
signal \N__25401\ : std_logic;
signal \N__25398\ : std_logic;
signal \N__25395\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25385\ : std_logic;
signal \N__25382\ : std_logic;
signal \N__25379\ : std_logic;
signal \N__25376\ : std_logic;
signal \N__25373\ : std_logic;
signal \N__25370\ : std_logic;
signal \N__25367\ : std_logic;
signal \N__25364\ : std_logic;
signal \N__25361\ : std_logic;
signal \N__25358\ : std_logic;
signal \N__25355\ : std_logic;
signal \N__25352\ : std_logic;
signal \N__25349\ : std_logic;
signal \N__25346\ : std_logic;
signal \N__25343\ : std_logic;
signal \N__25340\ : std_logic;
signal \N__25337\ : std_logic;
signal \N__25334\ : std_logic;
signal \N__25331\ : std_logic;
signal \N__25328\ : std_logic;
signal \N__25325\ : std_logic;
signal \N__25322\ : std_logic;
signal \N__25319\ : std_logic;
signal \N__25316\ : std_logic;
signal \N__25313\ : std_logic;
signal \N__25310\ : std_logic;
signal \N__25307\ : std_logic;
signal \N__25304\ : std_logic;
signal \N__25301\ : std_logic;
signal \N__25298\ : std_logic;
signal \N__25295\ : std_logic;
signal \N__25292\ : std_logic;
signal \N__25289\ : std_logic;
signal \N__25284\ : std_logic;
signal \N__25283\ : std_logic;
signal \N__25280\ : std_logic;
signal \N__25277\ : std_logic;
signal \N__25274\ : std_logic;
signal \N__25271\ : std_logic;
signal \N__25268\ : std_logic;
signal \N__25265\ : std_logic;
signal \N__25262\ : std_logic;
signal \N__25259\ : std_logic;
signal \N__25256\ : std_logic;
signal \N__25253\ : std_logic;
signal \N__25250\ : std_logic;
signal \N__25247\ : std_logic;
signal \N__25244\ : std_logic;
signal \N__25241\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25232\ : std_logic;
signal \N__25229\ : std_logic;
signal \N__25226\ : std_logic;
signal \N__25223\ : std_logic;
signal \N__25220\ : std_logic;
signal \N__25217\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25208\ : std_logic;
signal \N__25205\ : std_logic;
signal \N__25202\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25196\ : std_logic;
signal \N__25193\ : std_logic;
signal \N__25190\ : std_logic;
signal \N__25187\ : std_logic;
signal \N__25182\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25175\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25169\ : std_logic;
signal \N__25166\ : std_logic;
signal \N__25163\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25157\ : std_logic;
signal \N__25154\ : std_logic;
signal \N__25151\ : std_logic;
signal \N__25148\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25142\ : std_logic;
signal \N__25139\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25130\ : std_logic;
signal \N__25127\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25121\ : std_logic;
signal \N__25118\ : std_logic;
signal \N__25115\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25097\ : std_logic;
signal \N__25094\ : std_logic;
signal \N__25091\ : std_logic;
signal \N__25088\ : std_logic;
signal \N__25085\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25077\ : std_logic;
signal \N__25076\ : std_logic;
signal \N__25075\ : std_logic;
signal \N__25074\ : std_logic;
signal \N__25071\ : std_logic;
signal \N__25064\ : std_logic;
signal \N__25059\ : std_logic;
signal \N__25056\ : std_logic;
signal \N__25053\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25044\ : std_logic;
signal \N__25041\ : std_logic;
signal \N__25038\ : std_logic;
signal \N__25035\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25023\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25017\ : std_logic;
signal \N__25014\ : std_logic;
signal \N__25011\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__24998\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24974\ : std_logic;
signal \N__24971\ : std_logic;
signal \N__24968\ : std_logic;
signal \N__24965\ : std_logic;
signal \N__24962\ : std_logic;
signal \N__24959\ : std_logic;
signal \N__24956\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24950\ : std_logic;
signal \N__24947\ : std_logic;
signal \N__24944\ : std_logic;
signal \N__24941\ : std_logic;
signal \N__24938\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24932\ : std_logic;
signal \N__24929\ : std_logic;
signal \N__24926\ : std_logic;
signal \N__24923\ : std_logic;
signal \N__24920\ : std_logic;
signal \N__24917\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24911\ : std_logic;
signal \N__24908\ : std_logic;
signal \N__24905\ : std_logic;
signal \N__24902\ : std_logic;
signal \N__24899\ : std_logic;
signal \N__24896\ : std_logic;
signal \N__24891\ : std_logic;
signal \N__24888\ : std_logic;
signal \N__24887\ : std_logic;
signal \N__24884\ : std_logic;
signal \N__24881\ : std_logic;
signal \N__24876\ : std_logic;
signal \N__24873\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24858\ : std_logic;
signal \N__24855\ : std_logic;
signal \N__24852\ : std_logic;
signal \N__24849\ : std_logic;
signal \N__24846\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24840\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24836\ : std_logic;
signal \N__24833\ : std_logic;
signal \N__24830\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24822\ : std_logic;
signal \N__24819\ : std_logic;
signal \N__24818\ : std_logic;
signal \N__24815\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24804\ : std_logic;
signal \N__24803\ : std_logic;
signal \N__24800\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24782\ : std_logic;
signal \N__24779\ : std_logic;
signal \N__24776\ : std_logic;
signal \N__24773\ : std_logic;
signal \N__24770\ : std_logic;
signal \N__24767\ : std_logic;
signal \N__24764\ : std_logic;
signal \N__24761\ : std_logic;
signal \N__24758\ : std_logic;
signal \N__24755\ : std_logic;
signal \N__24752\ : std_logic;
signal \N__24749\ : std_logic;
signal \N__24746\ : std_logic;
signal \N__24743\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24737\ : std_logic;
signal \N__24734\ : std_logic;
signal \N__24731\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24722\ : std_logic;
signal \N__24719\ : std_logic;
signal \N__24716\ : std_logic;
signal \N__24713\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24702\ : std_logic;
signal \N__24699\ : std_logic;
signal \N__24698\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24679\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24671\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24665\ : std_logic;
signal \N__24662\ : std_logic;
signal \N__24661\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24657\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24651\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24639\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24629\ : std_logic;
signal \N__24624\ : std_logic;
signal \N__24621\ : std_logic;
signal \N__24620\ : std_logic;
signal \N__24619\ : std_logic;
signal \N__24616\ : std_logic;
signal \N__24613\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24605\ : std_logic;
signal \N__24602\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24596\ : std_logic;
signal \N__24593\ : std_logic;
signal \N__24588\ : std_logic;
signal \N__24585\ : std_logic;
signal \N__24584\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24564\ : std_logic;
signal \N__24557\ : std_logic;
signal \N__24554\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24548\ : std_logic;
signal \N__24545\ : std_logic;
signal \N__24542\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24533\ : std_logic;
signal \N__24532\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24523\ : std_logic;
signal \N__24520\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24513\ : std_logic;
signal \N__24510\ : std_logic;
signal \N__24505\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24491\ : std_logic;
signal \N__24488\ : std_logic;
signal \N__24485\ : std_logic;
signal \N__24484\ : std_logic;
signal \N__24483\ : std_logic;
signal \N__24478\ : std_logic;
signal \N__24475\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24467\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24459\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24453\ : std_logic;
signal \N__24452\ : std_logic;
signal \N__24449\ : std_logic;
signal \N__24446\ : std_logic;
signal \N__24445\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24434\ : std_logic;
signal \N__24431\ : std_logic;
signal \N__24430\ : std_logic;
signal \N__24425\ : std_logic;
signal \N__24422\ : std_logic;
signal \N__24417\ : std_logic;
signal \N__24414\ : std_logic;
signal \N__24411\ : std_logic;
signal \N__24408\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24392\ : std_logic;
signal \N__24391\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24387\ : std_logic;
signal \N__24384\ : std_logic;
signal \N__24381\ : std_logic;
signal \N__24378\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24372\ : std_logic;
signal \N__24369\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24359\ : std_logic;
signal \N__24354\ : std_logic;
signal \N__24353\ : std_logic;
signal \N__24350\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24345\ : std_logic;
signal \N__24342\ : std_logic;
signal \N__24339\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24328\ : std_logic;
signal \N__24323\ : std_logic;
signal \N__24318\ : std_logic;
signal \N__24317\ : std_logic;
signal \N__24314\ : std_logic;
signal \N__24311\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24304\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24293\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24287\ : std_logic;
signal \N__24284\ : std_logic;
signal \N__24279\ : std_logic;
signal \N__24276\ : std_logic;
signal \N__24275\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24262\ : std_logic;
signal \N__24259\ : std_logic;
signal \N__24256\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24248\ : std_logic;
signal \N__24245\ : std_logic;
signal \N__24240\ : std_logic;
signal \N__24239\ : std_logic;
signal \N__24236\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24232\ : std_logic;
signal \N__24231\ : std_logic;
signal \N__24228\ : std_logic;
signal \N__24225\ : std_logic;
signal \N__24222\ : std_logic;
signal \N__24219\ : std_logic;
signal \N__24216\ : std_logic;
signal \N__24213\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24203\ : std_logic;
signal \N__24198\ : std_logic;
signal \N__24197\ : std_logic;
signal \N__24194\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24189\ : std_logic;
signal \N__24186\ : std_logic;
signal \N__24183\ : std_logic;
signal \N__24180\ : std_logic;
signal \N__24177\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24167\ : std_logic;
signal \N__24164\ : std_logic;
signal \N__24159\ : std_logic;
signal \N__24158\ : std_logic;
signal \N__24155\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24150\ : std_logic;
signal \N__24147\ : std_logic;
signal \N__24144\ : std_logic;
signal \N__24141\ : std_logic;
signal \N__24138\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24128\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24120\ : std_logic;
signal \N__24119\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24117\ : std_logic;
signal \N__24114\ : std_logic;
signal \N__24111\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24105\ : std_logic;
signal \N__24102\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24083\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24077\ : std_logic;
signal \N__24074\ : std_logic;
signal \N__24073\ : std_logic;
signal \N__24070\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24066\ : std_logic;
signal \N__24063\ : std_logic;
signal \N__24060\ : std_logic;
signal \N__24057\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24047\ : std_logic;
signal \N__24042\ : std_logic;
signal \N__24041\ : std_logic;
signal \N__24038\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24033\ : std_logic;
signal \N__24030\ : std_logic;
signal \N__24027\ : std_logic;
signal \N__24024\ : std_logic;
signal \N__24021\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24011\ : std_logic;
signal \N__24006\ : std_logic;
signal \N__24005\ : std_logic;
signal \N__24002\ : std_logic;
signal \N__23999\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23988\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23979\ : std_logic;
signal \N__23976\ : std_logic;
signal \N__23967\ : std_logic;
signal \N__23964\ : std_logic;
signal \N__23963\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23961\ : std_logic;
signal \N__23958\ : std_logic;
signal \N__23955\ : std_logic;
signal \N__23952\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23946\ : std_logic;
signal \N__23943\ : std_logic;
signal \N__23940\ : std_logic;
signal \N__23937\ : std_logic;
signal \N__23934\ : std_logic;
signal \N__23927\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23921\ : std_logic;
signal \N__23920\ : std_logic;
signal \N__23917\ : std_logic;
signal \N__23914\ : std_logic;
signal \N__23913\ : std_logic;
signal \N__23910\ : std_logic;
signal \N__23907\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23888\ : std_logic;
signal \N__23883\ : std_logic;
signal \N__23882\ : std_logic;
signal \N__23879\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23861\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23855\ : std_logic;
signal \N__23852\ : std_logic;
signal \N__23847\ : std_logic;
signal \N__23844\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23840\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23836\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23830\ : std_logic;
signal \N__23827\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23819\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23815\ : std_logic;
signal \N__23812\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23799\ : std_logic;
signal \N__23798\ : std_logic;
signal \N__23795\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23790\ : std_logic;
signal \N__23787\ : std_logic;
signal \N__23784\ : std_logic;
signal \N__23781\ : std_logic;
signal \N__23778\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23768\ : std_logic;
signal \N__23763\ : std_logic;
signal \N__23760\ : std_logic;
signal \N__23757\ : std_logic;
signal \N__23754\ : std_logic;
signal \N__23751\ : std_logic;
signal \N__23748\ : std_logic;
signal \N__23745\ : std_logic;
signal \N__23742\ : std_logic;
signal \N__23739\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23726\ : std_logic;
signal \N__23721\ : std_logic;
signal \N__23720\ : std_logic;
signal \N__23717\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23698\ : std_logic;
signal \N__23693\ : std_logic;
signal \N__23690\ : std_logic;
signal \N__23685\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23681\ : std_logic;
signal \N__23678\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23674\ : std_logic;
signal \N__23671\ : std_logic;
signal \N__23668\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23660\ : std_logic;
signal \N__23659\ : std_logic;
signal \N__23654\ : std_logic;
signal \N__23651\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23640\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23628\ : std_logic;
signal \N__23625\ : std_logic;
signal \N__23622\ : std_logic;
signal \N__23621\ : std_logic;
signal \N__23618\ : std_logic;
signal \N__23615\ : std_logic;
signal \N__23610\ : std_logic;
signal \N__23607\ : std_logic;
signal \N__23606\ : std_logic;
signal \N__23603\ : std_logic;
signal \N__23600\ : std_logic;
signal \N__23597\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23591\ : std_logic;
signal \N__23588\ : std_logic;
signal \N__23587\ : std_logic;
signal \N__23582\ : std_logic;
signal \N__23579\ : std_logic;
signal \N__23574\ : std_logic;
signal \N__23573\ : std_logic;
signal \N__23568\ : std_logic;
signal \N__23565\ : std_logic;
signal \N__23564\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23547\ : std_logic;
signal \N__23546\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23529\ : std_logic;
signal \N__23528\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23507\ : std_logic;
signal \N__23506\ : std_logic;
signal \N__23503\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23497\ : std_logic;
signal \N__23490\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23486\ : std_logic;
signal \N__23485\ : std_logic;
signal \N__23480\ : std_logic;
signal \N__23477\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23471\ : std_logic;
signal \N__23468\ : std_logic;
signal \N__23463\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23454\ : std_logic;
signal \N__23451\ : std_logic;
signal \N__23450\ : std_logic;
signal \N__23449\ : std_logic;
signal \N__23448\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23446\ : std_logic;
signal \N__23443\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23441\ : std_logic;
signal \N__23438\ : std_logic;
signal \N__23433\ : std_logic;
signal \N__23428\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23406\ : std_logic;
signal \N__23405\ : std_logic;
signal \N__23404\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23402\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23390\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23383\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23367\ : std_logic;
signal \N__23366\ : std_logic;
signal \N__23363\ : std_logic;
signal \N__23360\ : std_logic;
signal \N__23357\ : std_logic;
signal \N__23354\ : std_logic;
signal \N__23349\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23347\ : std_logic;
signal \N__23344\ : std_logic;
signal \N__23341\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23331\ : std_logic;
signal \N__23328\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23316\ : std_logic;
signal \N__23313\ : std_logic;
signal \N__23310\ : std_logic;
signal \N__23309\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23301\ : std_logic;
signal \N__23298\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23288\ : std_logic;
signal \N__23285\ : std_logic;
signal \N__23282\ : std_logic;
signal \N__23279\ : std_logic;
signal \N__23276\ : std_logic;
signal \N__23273\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23262\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23247\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23235\ : std_logic;
signal \N__23232\ : std_logic;
signal \N__23229\ : std_logic;
signal \N__23226\ : std_logic;
signal \N__23223\ : std_logic;
signal \N__23220\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23214\ : std_logic;
signal \N__23211\ : std_logic;
signal \N__23208\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23196\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23184\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23169\ : std_logic;
signal \N__23166\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23154\ : std_logic;
signal \N__23151\ : std_logic;
signal \N__23148\ : std_logic;
signal \N__23145\ : std_logic;
signal \N__23142\ : std_logic;
signal \N__23139\ : std_logic;
signal \N__23136\ : std_logic;
signal \N__23133\ : std_logic;
signal \N__23130\ : std_logic;
signal \N__23127\ : std_logic;
signal \N__23124\ : std_logic;
signal \N__23121\ : std_logic;
signal \N__23118\ : std_logic;
signal \N__23115\ : std_logic;
signal \N__23112\ : std_logic;
signal \N__23109\ : std_logic;
signal \N__23106\ : std_logic;
signal \N__23103\ : std_logic;
signal \N__23100\ : std_logic;
signal \N__23097\ : std_logic;
signal \N__23094\ : std_logic;
signal \N__23091\ : std_logic;
signal \N__23088\ : std_logic;
signal \N__23087\ : std_logic;
signal \N__23084\ : std_logic;
signal \N__23081\ : std_logic;
signal \N__23078\ : std_logic;
signal \N__23075\ : std_logic;
signal \N__23070\ : std_logic;
signal \N__23067\ : std_logic;
signal \N__23064\ : std_logic;
signal \N__23061\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23055\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23043\ : std_logic;
signal \N__23040\ : std_logic;
signal \N__23037\ : std_logic;
signal \N__23034\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23022\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23009\ : std_logic;
signal \N__23004\ : std_logic;
signal \N__23001\ : std_logic;
signal \N__22998\ : std_logic;
signal \N__22995\ : std_logic;
signal \N__22992\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22986\ : std_logic;
signal \N__22985\ : std_logic;
signal \N__22978\ : std_logic;
signal \N__22973\ : std_logic;
signal \N__22968\ : std_logic;
signal \N__22965\ : std_logic;
signal \N__22962\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22958\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22954\ : std_logic;
signal \N__22951\ : std_logic;
signal \N__22948\ : std_logic;
signal \N__22941\ : std_logic;
signal \N__22938\ : std_logic;
signal \N__22935\ : std_logic;
signal \N__22932\ : std_logic;
signal \N__22929\ : std_logic;
signal \N__22926\ : std_logic;
signal \N__22923\ : std_logic;
signal \N__22922\ : std_logic;
signal \N__22919\ : std_logic;
signal \N__22916\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22908\ : std_logic;
signal \N__22905\ : std_logic;
signal \N__22902\ : std_logic;
signal \N__22899\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22887\ : std_logic;
signal \N__22884\ : std_logic;
signal \N__22883\ : std_logic;
signal \N__22882\ : std_logic;
signal \N__22879\ : std_logic;
signal \N__22876\ : std_logic;
signal \N__22873\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22860\ : std_logic;
signal \N__22859\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22856\ : std_logic;
signal \N__22855\ : std_logic;
signal \N__22852\ : std_logic;
signal \N__22847\ : std_logic;
signal \N__22840\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22830\ : std_logic;
signal \N__22827\ : std_logic;
signal \N__22826\ : std_logic;
signal \N__22825\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22805\ : std_logic;
signal \N__22804\ : std_logic;
signal \N__22801\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22788\ : std_logic;
signal \N__22787\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22767\ : std_logic;
signal \N__22764\ : std_logic;
signal \N__22763\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22755\ : std_logic;
signal \N__22752\ : std_logic;
signal \N__22751\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22745\ : std_logic;
signal \N__22744\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22734\ : std_logic;
signal \N__22731\ : std_logic;
signal \N__22724\ : std_logic;
signal \N__22713\ : std_logic;
signal \N__22712\ : std_logic;
signal \N__22707\ : std_logic;
signal \N__22706\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22704\ : std_logic;
signal \N__22703\ : std_logic;
signal \N__22700\ : std_logic;
signal \N__22697\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22683\ : std_logic;
signal \N__22682\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22673\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22665\ : std_logic;
signal \N__22662\ : std_logic;
signal \N__22659\ : std_logic;
signal \N__22658\ : std_logic;
signal \N__22653\ : std_logic;
signal \N__22650\ : std_logic;
signal \N__22649\ : std_logic;
signal \N__22646\ : std_logic;
signal \N__22643\ : std_logic;
signal \N__22638\ : std_logic;
signal \N__22637\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22626\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22614\ : std_logic;
signal \N__22611\ : std_logic;
signal \N__22608\ : std_logic;
signal \N__22605\ : std_logic;
signal \N__22602\ : std_logic;
signal \N__22599\ : std_logic;
signal \N__22596\ : std_logic;
signal \N__22593\ : std_logic;
signal \N__22590\ : std_logic;
signal \N__22587\ : std_logic;
signal \N__22584\ : std_logic;
signal \N__22581\ : std_logic;
signal \N__22578\ : std_logic;
signal \N__22575\ : std_logic;
signal \N__22572\ : std_logic;
signal \N__22569\ : std_logic;
signal \N__22566\ : std_logic;
signal \N__22563\ : std_logic;
signal \N__22560\ : std_logic;
signal \N__22557\ : std_logic;
signal \N__22554\ : std_logic;
signal \N__22551\ : std_logic;
signal \N__22548\ : std_logic;
signal \N__22545\ : std_logic;
signal \N__22542\ : std_logic;
signal \N__22539\ : std_logic;
signal \N__22536\ : std_logic;
signal \N__22533\ : std_logic;
signal \N__22530\ : std_logic;
signal \N__22527\ : std_logic;
signal \N__22524\ : std_logic;
signal \N__22521\ : std_logic;
signal \N__22518\ : std_logic;
signal \N__22517\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22500\ : std_logic;
signal \N__22499\ : std_logic;
signal \N__22496\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22488\ : std_logic;
signal \N__22487\ : std_logic;
signal \N__22482\ : std_logic;
signal \N__22479\ : std_logic;
signal \N__22476\ : std_logic;
signal \N__22475\ : std_logic;
signal \N__22474\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22455\ : std_logic;
signal \N__22452\ : std_logic;
signal \N__22449\ : std_logic;
signal \N__22446\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22437\ : std_logic;
signal \N__22434\ : std_logic;
signal \N__22433\ : std_logic;
signal \N__22430\ : std_logic;
signal \N__22427\ : std_logic;
signal \N__22424\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22416\ : std_logic;
signal \N__22415\ : std_logic;
signal \N__22414\ : std_logic;
signal \N__22413\ : std_logic;
signal \N__22412\ : std_logic;
signal \N__22405\ : std_logic;
signal \N__22400\ : std_logic;
signal \N__22395\ : std_logic;
signal \N__22392\ : std_logic;
signal \N__22389\ : std_logic;
signal \N__22386\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22374\ : std_logic;
signal \N__22371\ : std_logic;
signal \N__22368\ : std_logic;
signal \N__22365\ : std_logic;
signal \N__22362\ : std_logic;
signal \N__22359\ : std_logic;
signal \N__22356\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22350\ : std_logic;
signal \N__22347\ : std_logic;
signal \N__22344\ : std_logic;
signal \N__22341\ : std_logic;
signal \N__22338\ : std_logic;
signal \N__22335\ : std_logic;
signal \N__22332\ : std_logic;
signal \N__22329\ : std_logic;
signal \N__22326\ : std_logic;
signal clock_ibuf_gb_io_gb_input : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal mcu_sclk_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net\ : std_logic;
signal \bfn_5_16_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_17_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_375\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_i\ : std_logic;
signal \N_1821_0\ : std_logic;
signal sdin1_c : std_logic;
signal sdin0_c : std_logic;
signal mcu_data_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93Z0Z_0_cascade_\ : std_logic;
signal sclk1_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32Z0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.un2_count_bits_1_0_a2_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_8\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\ : std_logic;
signal \bfn_6_18_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4\ : std_logic;
signal \bfn_6_19_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_333\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_376\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.dout_read\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_237_cascade_\ : std_logic;
signal \N_85_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_3\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_370_i\ : std_logic;
signal \N_1820_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_u_i_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.sclk_u_i_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_7 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_7 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_7_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_7\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_7_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_7\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1Z0Z_23_cascade_\ : std_logic;
signal \N_29\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_read\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01Z0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_reti_0_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_8\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_369_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.csb_u_i_a2_0_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_331_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.m7_0_a2_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_459_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_8 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_466_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_448_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1826_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_5 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_5\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_6 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_6\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_7 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_7\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1827_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_7 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_863\ : std_logic;
signal s1_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_iZ0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_596_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_597\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_oZ0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1615_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.csb_u_i_a2_0_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0\ : std_logic;
signal \N_1822_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.csb_u_i_a2_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0\ : std_logic;
signal \bfn_9_19_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_a2_1_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_22\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_op\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0\ : std_logic;
signal \bfn_9_22_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_391_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_455_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_454_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_453_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_463_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_1 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_1 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_1_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_1 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_1_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_1_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_5_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_5\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_5 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_5 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_5_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_6\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_21\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_22\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.dout_op\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_12\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_15\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_10\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_391\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_1\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_10 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_3_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_3 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_3 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_3_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_31 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_31 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_31_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_31\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_31_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_31\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_27 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_28 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_29 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_30 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_31 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_31\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_3 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_4 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_4\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_4_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_4\ : std_logic;
signal \bfn_11_15_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m7_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996_cascade_\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0\ : std_logic;
signal \bfn_11_19_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_3\ : std_logic;
signal sync_50hz_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_410_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_68_0_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_8 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_8 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_8_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_8_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_8\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_14 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_14 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_14_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_14 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_14_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_14_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_14\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_22 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_30 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_30 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_30_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_30\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_30_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_30\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_30\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_30\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_30\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_31 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_31\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_31\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_4\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_4 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_26 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_26 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_26 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_0_26\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_1_26_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_26 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_21 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_29 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_3 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_907\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_30 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_621\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_31 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_610\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_1 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_316\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_5 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_885\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_6 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_874\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_4 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_4 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_4\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_30 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_4 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_8 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_0 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_11 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_12 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_13 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_14 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_786\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_15 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_20 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15Z0Z_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_19\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_i_a2_1_1_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9\ : std_logic;
signal \bfn_12_20_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.en_ch_cnt_0_a2_0_a2_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1867_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un40_0_a2_4_a2_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16\ : std_logic;
signal sda_o : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_22_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_22\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_22 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_22 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_22\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_22\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_22\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_28 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_28 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_28_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_28\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_28_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_28\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_28\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_15 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_15 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_15_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_15 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_775\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_15_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_15_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_15\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_23 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_17 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_17 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_17_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_17 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_17_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_17_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_17\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_25 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_4_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_4_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_4 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRLZ0Z7_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_6_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_6\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_6 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_6 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_841\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_9_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_6_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3QZ0Z5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_5\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1615\ : std_logic;
signal \N_1614_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_28 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_643\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_5\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_4 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_896\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_291_reti_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_276i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_retZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_4_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_2_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_0_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_o3_i_a2_1_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_5\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ns_i_a2_1_1_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_2\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_2_cascade_\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_10\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_68_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_410_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_state_7\ : std_logic;
signal \bfn_13_23_0_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetterZ0\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_Control_StartUp_inst.rst_neg_i\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_22\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_2 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_13 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_13 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_13_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_13 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_797\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_13_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_13_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_18 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_18 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_18_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_18_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_18\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_18\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_15\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_13_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3QZ0Z5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_4\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_4\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_9\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_22 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3Z0Z_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1959_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0_cascade_\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_Control_StartUp_inst.N_8_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.en_count_bits_0_i_a2_0_a2_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_277_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_18\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967i_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_276_reti\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_8_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_2_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1945\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1844\ : std_logic;
signal \N_528_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.n_state41\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_state_19\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_275_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_275_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_2_cascade_\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_59\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_2\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_2 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_2 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_2_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_2_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_2\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_10 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_10 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_10_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_10 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_830\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_10_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_10_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_10\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_18 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_18\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_11 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_11 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_11_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_11 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_819\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_11_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_11_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_19 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_20 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_20 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_20_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_20 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_283\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_20_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_20_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_6\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_6 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_6_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRLZ0Z7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_7\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_6\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_6 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_5 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_5 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRLZ0Z7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_5\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_5 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_14 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_242_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_5 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_16 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_18 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1911\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_8 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1920\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m20_0_a2_4_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_11_0_i_0_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1394_cascade_\ : std_logic;
signal s_sda_i_g : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1392\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1381_0_cascade_\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_state_i_2_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.end_conf_a\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1817_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_0_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1873_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1874_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_2_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1950\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1949_cascade_\ : std_logic;
signal stop_fpga2_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.end_conf_b\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_112\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_4\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_111\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_119\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_120\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_36\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_118\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_37\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_38\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_33\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_34\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_35\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_76\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_17 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_753\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_19 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_2 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_918\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_22 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_698\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_23 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_2\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_25 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_27 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_19 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_19 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_731\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_19\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_19_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_19\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_19\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_19\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_0 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_0 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_0_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_21 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_1\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_18 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_18\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_20 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_20\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_15_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_14\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_14_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGHZ0Z5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_14_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_14\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_14 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_23_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDDZ0Z7_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_6 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_6\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_3 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_4 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_6 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_0Z0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_30\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1654_cascade_\ : std_logic;
signal \N_12_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_7 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0_cascade_\ : std_logic;
signal \N_12_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_0_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_1786_2\ : std_logic;
signal \N_979\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_id_prdata_1_4_u_i_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2_cascade_\ : std_logic;
signal \N_1838_0_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1379_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1400_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1374_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1399_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1395_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_0_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1409_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1372_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1880\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1848_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1884_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392_reti\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0_a2_6_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_li_0_1\ : std_logic;
signal \c_state_ret_12_RNIDMPS1_0\ : std_logic;
signal \c_state_ret_12_RNIDMPS1_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.clr_sys_reg\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_1 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_349\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_7\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_31\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_32\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_113\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_114\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_110\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_39\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_77\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_78\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_40\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_67\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_68\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_115\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_116\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_117\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa\ : std_logic;
signal rst_n_c_i : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_12 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_12 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_12_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_12 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_808\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_12_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_12\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_12_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_12\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_11 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_11\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_12 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_12\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_13 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_13\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_14 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_14\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_15 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_15\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_16 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_17 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_17\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_2 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_2\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_24 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_24\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_19 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_19\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_25 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_27 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_27\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_28 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_28\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_28\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_29 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_29\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_3 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_3 : std_logic;
signal serial_out_testing_c : std_logic;
signal rst_n_c : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1965\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_522_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.start_conf_b\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_20 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_20_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DDZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_22\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_conf\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1831_0\ : std_logic;
signal \N_1614\ : std_logic;
signal \N_1841_0_cascade_\ : std_logic;
signal \N_1613_cascade_\ : std_logic;
signal \N_1860_0\ : std_logic;
signal \N_202_0\ : std_logic;
signal \N_1859_0\ : std_logic;
signal \N_1861_0\ : std_logic;
signal \N_1613\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_604\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.s_command_4\ : std_logic;
signal \I2C_top_level_inst1.s_command_5\ : std_logic;
signal \I2C_top_level_inst1.s_command_6\ : std_logic;
signal \N_1803\ : std_logic;
signal \N_1803_cascade_\ : std_logic;
signal \I2C_top_level_inst1.s_command_7\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6Z0Z_26\ : std_logic;
signal \I2C_top_level_inst1.N_327_i\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_113_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4\ : std_logic;
signal \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_3_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_5_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_2_1\ : std_logic;
signal \I2C_top_level_inst1.N_4_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.N_259\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1848_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7Z0Z_26\ : std_logic;
signal \I2C_top_level_inst1.s_sda_o_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.s_sda_o_txZ0\ : std_logic;
signal \I2C_top_level_inst1.s_sda_o_qZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.start_conf_a\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1855_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1855_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1857_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1857_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_384\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1854_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1840_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_383\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8Z0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_state_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1862\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.N_1816_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_state_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_reti_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_6\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_11\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_48\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_51\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_10\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_55\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_121\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_14\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_12\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_13\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_8\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_9\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_15\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_79\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_16\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_17\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_18\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_107\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_69\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_106\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_47\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_94\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_104\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_105\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_46\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_91\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_92\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_93\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_95\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_96\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_97\ : std_logic;
signal enable_config_c : std_logic;
signal elec_config_out_c : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_24\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_24_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_24\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_24 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_24 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_24_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_24\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_23 : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_10 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_10\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_24 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_676\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_23\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_687\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_23\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_23_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_23\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_23 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_23 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_23_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_23\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_20\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_21 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_21 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_21_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_21 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1320\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1896\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_21_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_21\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_21\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_21_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_30\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_13 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_31\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_14 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_22_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_22\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_22 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_22_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDDZ0Z7\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_22 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_22\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_20 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_30\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_22 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_8_0_m2_ns_1_cascade_\ : std_logic;
signal \N_1842_0\ : std_logic;
signal \N_1842_0_cascade_\ : std_logic;
signal \N_1841_0\ : std_logic;
signal \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C_net\ : std_logic;
signal \bfn_18_18_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_CO\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_addr_RNI3UAS1_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.c_addr_RNI50BS1_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93STZ0Z1\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rstZ0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNOZ0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_3_cascade_\ : std_logic;
signal \N_1975\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNOZ0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0\ : std_logic;
signal \bfn_18_20_0_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.paddr_fsm_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_2 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_3 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_4 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_5 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_6 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_7\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_8 : std_logic;
signal \bfn_18_21_0_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_9 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_10 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_11 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_12 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_13 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_14 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_14\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_paddr_fsm_15 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_86\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_54\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_s_data_system_o_0 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_52\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_53\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_87\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_88\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_49\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_50\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_89\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_90\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_85\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_1\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_101\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_66\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_102\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_103\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_84\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_41\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_100\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_42\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_43\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_44\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_45\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_70\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_71\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_74\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_75\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_98\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_99\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_72\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_73\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_83\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_82\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_80\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_81\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_29 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_29 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_29_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_29\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_29\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_29_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_632\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_29\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_29\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_7 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_8_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_6\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_7\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_24\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_28\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_1Z0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_27\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_7\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_7 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_8\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_8 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_8 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_8 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_8_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8DZ0Z7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14_cascade_\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_8 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_20\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_20 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_12 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_0_12_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_2_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_0_i_12_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_13\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_13 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_13\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_5 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_6 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_7 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_8 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_12\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_12 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_12 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_12\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_11_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFHZ0Z5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_1\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_2\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_3\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_4\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_5\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_6\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_7\ : std_logic;
signal \I2C_top_level_inst1.s_load_addr1\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_3\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_4\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_4\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_5\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_5\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_6\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_6\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_7\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_7\ : std_logic;
signal \N_396\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_4_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNOZ0Z_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.s_no_restart\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_304_0\ : std_logic;
signal \I2C_top_level_inst1.s_ack\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_6\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_5\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_2\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_3\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_4\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_21\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_27\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_22\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_23\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_108\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_109\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_19\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_20\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_24\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_124\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_125\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_122\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_123\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_25\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_26\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_27 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_27 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_27_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_27\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_27\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_27_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_654\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_27\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_27\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_16 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_16 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_16_cascade_\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_16 : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_16 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_764\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_16_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_16\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_16\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_16_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_16\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_24 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_24\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_22 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_4 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_5 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_6 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_15_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_14\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_15\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_4 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_20 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_20 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_12 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_22 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_14 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_15 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_16 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_11 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_11 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_11_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_13\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_13 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_23\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_10 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_10 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_2 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_2 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_11 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_11\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_11 : std_logic;
signal \bfn_20_17_0_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_CO\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_4\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_7\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7\ : std_logic;
signal \bfn_20_18_0_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_12\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_15\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_103_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_291_cascade_\ : std_logic;
signal \I2C_top_level_inst1.s_load_addr0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_6_0_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1378\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_1676_cascade_\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21\ : std_logic;
signal \c_state_RNIEVJ7_22_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_77_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_300_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_FSM_inst.N_1425_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_64\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_65\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_128\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_126\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_127\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_28\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_29\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_30\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_62\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_63\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_58\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_59\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_60\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_61\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_56\ : std_logic;
signal \serializer_mod_inst.shift_regZ0Z_57\ : std_logic;
signal \serializer_mod_inst.un22_next_state_1_cascade_\ : std_logic;
signal \serializer_mod_inst.un22_next_state\ : std_logic;
signal \serializer_mod_inst.current_stateZ0Z_1\ : std_logic;
signal \serializer_mod_inst.current_stateZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_0 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_940\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_25\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_3Z0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_16\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_7 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_7\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_17_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_16\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_17 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_11\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_21_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LHZ0Z5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_21 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_21 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_21_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDDZ0Z7\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_21 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_21 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_21\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_11 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_12 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_21 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_30\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_13 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_31\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_15 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_13 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_31\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_15 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_24\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_17 : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_10\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_9 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i_cascade_\ : std_logic;
signal \s_paddr_I2C_5\ : std_logic;
signal \s_paddr_I2C_4\ : std_logic;
signal \s_paddr_I2C_6\ : std_logic;
signal \s_paddr_I2C_7\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_5\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_2_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_1_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0_cascade_\ : std_logic;
signal \s_paddr_I2C_2\ : std_logic;
signal \s_paddr_I2C_1\ : std_logic;
signal \s_paddr_I2C_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_7_3_i_a2_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0\ : std_logic;
signal \I2C_top_level_inst1.s_addr1_o_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_8_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_CO\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1651\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1652\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_0_4_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_0_1_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_279_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_0_1_7_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_268_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_10_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_18_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1605_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_0\ : std_logic;
signal \I2C_top_level_inst1.s_command_0\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_1\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_2\ : std_logic;
signal \I2C_top_level_inst1.s_data_ireg_3\ : std_logic;
signal scl_c_g : std_logic;
signal \I2C_top_level_inst1.s_load_command\ : std_logic;
signal \serializer_mod_inst.un1_counter_srlto6_3\ : std_logic;
signal \serializer_mod_inst.un1_counter_srlto6_4_cascade_\ : std_logic;
signal \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\ : std_logic;
signal \serializer_mod_inst.un22_next_state_5\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_0\ : std_logic;
signal \bfn_21_27_0_\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_1\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_0\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_2\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_1\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_3\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_2\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_4\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_3\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_5\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_4\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_6\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_5\ : std_logic;
signal \serializer_mod_inst.next_state32_i\ : std_logic;
signal \serializer_mod_inst.counter_sr_cry_6\ : std_logic;
signal \serializer_mod_inst.counter_srZ0Z_7\ : std_logic;
signal \serializer_mod_inst.counter_sre_0_i\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_15 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_24\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_2Z0Z_26\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_27\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_28\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_29\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_7 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_19 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_19 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_0 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_0 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_18 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_18_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9DZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_19\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_18 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_27\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_28\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_29\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_23 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_23 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_23_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.dout_conf\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALHZ0Z5\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_21\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_22\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_23 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_23 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_23\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_9 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_10 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_10 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_10 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_10_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_10\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_9 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_8\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_9\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_2 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_3 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_3 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_3 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_3\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_2 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_2\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_6_0_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_607\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_15_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_1_15\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_322\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_267\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_394\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_267_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_1_1_i_m2_1_9_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_101\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_1_2_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_372_cascade_\ : std_logic;
signal \N_409\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_a3_1_0_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_412_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_1_14\ : std_logic;
signal \N_410\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_1_0_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_24_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_11_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_11_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_2_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_86_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_95_0\ : std_logic;
signal \I2C_top_level_inst1.s_stop\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_844_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1754_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_1\ : std_logic;
signal scl_c : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0\ : std_logic;
signal \I2C_top_level_inst1.s_command_1\ : std_logic;
signal \I2C_top_level_inst1.s_command_2\ : std_logic;
signal \I2C_top_level_inst1.s_command_3\ : std_logic;
signal \I2C_top_level_inst1.s_load_wdata\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.s_start\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.s_r_w\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_27\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_29\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_23 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_19\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_19 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_19 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_19\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_18 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_18 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_18 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_18_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_18\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_25 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_25 : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_25_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_25_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_665\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_25\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_16 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_17 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_17 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_17_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_17\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_16 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGHZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_15\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_16\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_31\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_14 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_15 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_24\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_16 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_28\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_17 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_2 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RLZ0Z7_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_2\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkstopmask_1 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_clkctrovf_1 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_3_26\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_4093_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_26\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_g\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0\ : std_logic;
signal \s_paddr_I2C_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_230_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_0_sqmuxa\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_2_sqmuxa\ : std_logic;
signal \s_paddr_I2C_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_230\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_4\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_365_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_4_0_a2_2_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_676_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_address\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1606_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1565_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_5_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_6_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_7_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_11_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_23_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_288\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_288_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_23\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_115\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_904\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un30_i_a2_9_a2_4_a2_0_1_2_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_291\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_0_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_232_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_2_1_cascade_\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_20\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_4_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_232\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_1_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_2_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_231\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_212\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_211\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1653_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_122_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_208\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_239\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_239_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_294\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_1_0_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_0_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1776\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_209\ : std_logic;
signal s_sda_i : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_16\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_15\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_15\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_16\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_17\ : std_logic;
signal \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_19 : std_logic;
signal \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_29\ : std_logic;
signal \N_1592_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_9\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_10\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_10\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_11\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_11\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_12\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_14\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_14\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_13\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_12\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_13\ : std_logic;
signal \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_0 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_0 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_interrupts_1 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_config_1 : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_1 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_1\ : std_logic;
signal cemf_module_64ch_ctrl_inst1_data_coarseovf_0 : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2QZ0Z5_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0_cascade_\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_0\ : std_logic;
signal \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net\ : std_logic;
signal \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_18\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_17\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_18\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_19\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_20\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_19\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_20\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_21\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_21\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_22\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_22\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_23\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_23\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_24\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_24\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_25\ : std_logic;
signal \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_25\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_26\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_26\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_27\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_27\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_28\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_28\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_29\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_29\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_30\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_30\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_31\ : std_logic;
signal \I2C_top_level_inst1.s_sda_o_reg\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_0\ : std_logic;
signal \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_1\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_2\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_3\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_3\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_4\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_4\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_5\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_5\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_6\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_6\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_7\ : std_logic;
signal \I2C_top_level_inst1.s_enable_desp_tx\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_7\ : std_logic;
signal \I2C_top_level_inst1_s_data_oreg_8\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_8\ : std_logic;
signal \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\ : std_logic;
signal \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0\ : std_logic;
signal rst_n_c_i_g : std_logic;
signal \c_state_RNIEVJ7_22\ : std_logic;
signal \I2C_top_level_inst1.s_load_rdata2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o3_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1802\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1609_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0\ : std_logic;
signal \I2C_top_level_inst1.s_addr0_o_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_691\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_295_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_277\ : std_logic;
signal \N_552_i\ : std_logic;
signal \N_1838_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_295\ : std_logic;
signal \N_73_i_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1_s_burst\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_19\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_274_cascade_\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_276\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_245\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1669_cascade_\ : std_logic;
signal clock_c_g : std_logic;
signal \I2C_top_level_inst1.c_state4_0_i_g\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_2_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_0_2_cascade_\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0\ : std_logic;
signal \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666_2\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal next_sequence_wire : std_logic;
signal stop_fpga2_wire : std_logic;
signal stop1_wire : std_logic;
signal s0_wire : std_logic;
signal mcu_data_wire : std_logic;
signal start1_wire : std_logic;
signal rst_n_wire : std_logic;
signal scl_wire : std_logic;
signal dout0_wire : std_logic;
signal stop0_wire : std_logic;
signal s2_wire : std_logic;
signal mcu_sclk_wire : std_logic;
signal frame_sync_wire : std_logic;
signal sdin0_wire : std_logic;
signal sdin1_wire : std_logic;
signal dout1_wire : std_logic;
signal csb1_wire : std_logic;
signal sclk1_wire : std_logic;
signal sclk0_wire : std_logic;
signal s1_wire : std_logic;
signal enable_config_wire : std_logic;
signal sync_50hz_wire : std_logic;
signal serial_out_testing_wire : std_logic;
signal start0_wire : std_logic;
signal s3_wire : std_logic;
signal elec_config_out_wire : std_logic;
signal csb0_wire : std_logic;
signal clock_wire : std_logic;
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_WDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_WADDR_wire\ : std_logic_vector(10 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_MASK_wire\ : std_logic_vector(15 downto 0);
signal \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_WDATA_wire\ : std_logic_vector(15 downto 0);

begin
    next_sequence <= next_sequence_wire;
    stop_fpga2 <= stop_fpga2_wire;
    stop1 <= stop1_wire;
    s0 <= s0_wire;
    mcu_data <= mcu_data_wire;
    start1 <= start1_wire;
    rst_n_wire <= rst_n;
    scl_wire <= scl;
    dout0 <= dout0_wire;
    stop0 <= stop0_wire;
    s2 <= s2_wire;
    mcu_sclk <= mcu_sclk_wire;
    frame_sync <= frame_sync_wire;
    sdin0_wire <= sdin0;
    sdin1_wire <= sdin1;
    dout1 <= dout1_wire;
    csb1 <= csb1_wire;
    sclk1 <= sclk1_wire;
    sclk0 <= sclk0_wire;
    s1 <= s1_wire;
    enable_config <= enable_config_wire;
    sync_50hz_wire <= sync_50hz;
    serial_out_testing <= serial_out_testing_wire;
    start0 <= start0_wire;
    s3 <= s3_wire;
    elec_config_out <= elec_config_out_wire;
    csb0 <= csb0_wire;
    clock_wire <= clock;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_15 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_14 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_13 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_12 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_11 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_10 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_9 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_8 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_7 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_6 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_5 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_4 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_3 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_2 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_1 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_0 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24740\&\N__24935\&\N__25112\&\N__25316\&\N__36044\&\N__25214\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24731\&\N__24932\&\N__25109\&\N__25313\&\N__36041\&\N__25211\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_WDATA_wire\ <= \N__23921\&\N__23963\&\N__24005\&\N__24042\&\N__24483\&\N__24697\&\N__24275\&\N__26186\&\N__33976\&\N__26384\&\N__24353\&\N__24392\&\N__23798\&\N__24619\&\N__23684\&\N__23721\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_31 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_30 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_29 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_28 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_27 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_26 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_25 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_24 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_23 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_22 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_21 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_20 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_19 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_18 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_17 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_16 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24728\&\N__24923\&\N__25100\&\N__25304\&\N__36032\&\N__25202\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24719\&\N__24920\&\N__25097\&\N__25301\&\N__36029\&\N__25199\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_WDATA_wire\ <= \N__26553\&\N__24666\&\N__24077\&\N__24445\&\N__24533\&\N__24158\&\N__24240\&\N__24584\&\N__24198\&\N__24317\&\N__24119\&\N__23841\&\N__26424\&\N__26469\&\N__26514\&\N__23883\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_31 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_30 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_29 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_28 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_27 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_26 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_25 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_24 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_23 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_22 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_21 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_20 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_19 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_18 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_17 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_16 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24800\&\N__24995\&\N__25172\&\N__25376\&\N__36104\&\N__25274\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24791\&\N__24992\&\N__25169\&\N__25373\&\N__36101\&\N__25271\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_WDATA_wire\ <= \N__26552\&\N__24665\&\N__24078\&\N__24459\&\N__24534\&\N__24159\&\N__24239\&\N__24588\&\N__24197\&\N__24318\&\N__24120\&\N__23840\&\N__26419\&\N__26464\&\N__26509\&\N__23882\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_15 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_14 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_13 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_12 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_11 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_10 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_9 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_8 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_7 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_6 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_5 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_4 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_3 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_2 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_1 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_0 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24807\&\N__25005\&\N__25182\&\N__25386\&\N__36114\&\N__25284\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24803\&\N__25004\&\N__25181\&\N__25385\&\N__36113\&\N__25283\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_WDATA_wire\ <= \N__23922\&\N__23964\&\N__24006\&\N__24041\&\N__24495\&\N__24702\&\N__24279\&\N__26187\&\N__34005\&\N__26385\&\N__24354\&\N__24393\&\N__23799\&\N__24624\&\N__23685\&\N__23720\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_31 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_30 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_29 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_28 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_27 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_26 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_25 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_24 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_23 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_22 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_21 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_20 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_19 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_18 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_17 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_16 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24752\&\N__24947\&\N__25124\&\N__25328\&\N__36056\&\N__25226\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24743\&\N__24944\&\N__25121\&\N__25325\&\N__36053\&\N__25223\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_WDATA_wire\ <= \N__26548\&\N__24661\&\N__24069\&\N__24430\&\N__24513\&\N__24150\&\N__24235\&\N__24564\&\N__24193\&\N__24310\&\N__24117\&\N__23836\&\N__26420\&\N__26465\&\N__26510\&\N__23878\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_15 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_14 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_13 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_12 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_11 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_10 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_9 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_8 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_7 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_6 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_5 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_4 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_3 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_2 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_1 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_0 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24788\&\N__24983\&\N__25160\&\N__25364\&\N__36092\&\N__25262\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24779\&\N__24980\&\N__25157\&\N__25361\&\N__36089\&\N__25259\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_WDATA_wire\ <= \N__23920\&\N__23961\&\N__23998\&\N__24033\&\N__24491\&\N__24698\&\N__24274\&\N__26182\&\N__34001\&\N__26380\&\N__24349\&\N__24387\&\N__23794\&\N__24620\&\N__23659\&\N__23698\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_15 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_14 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_13 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_12 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_11 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_10 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_9 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_8 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_7 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_6 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_5 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_4 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_3 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_2 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_1 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_0 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24764\&\N__24959\&\N__25136\&\N__25340\&\N__36068\&\N__25238\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24755\&\N__24956\&\N__25133\&\N__25337\&\N__36065\&\N__25235\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_WDATA_wire\ <= \N__23913\&\N__23962\&\N__23991\&\N__24037\&\N__24484\&\N__24679\&\N__24255\&\N__26169\&\N__33994\&\N__26376\&\N__24345\&\N__24391\&\N__23790\&\N__24601\&\N__23677\&\N__23716\;
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_31 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(15);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_30 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(14);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_29 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(13);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_28 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(12);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_27 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(11);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_26 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(10);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_25 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(9);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_24 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(8);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_23 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(7);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_22 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(6);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_21 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(5);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_20 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(4);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_19 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(3);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_18 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(2);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_17 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(1);
    cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_16 <= \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\(0);
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24776\&\N__24971\&\N__25148\&\N__25352\&\N__36080\&\N__25250\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_WADDR_wire\ <= '0'&'0'&'0'&'0'&'0'&\N__24767\&\N__24968\&\N__25145\&\N__25349\&\N__36077\&\N__25247\;
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_MASK_wire\ <= '0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0'&'0';
    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_WDATA_wire\ <= \N__26538\&\N__24657\&\N__24073\&\N__24452\&\N__24532\&\N__24154\&\N__24231\&\N__24583\&\N__24189\&\N__24292\&\N__24118\&\N__23818\&\N__26412\&\N__26457\&\N__26502\&\N__23860\;

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65640\,
            RE => \N__39325\,
            WCLKE => \N__24887\,
            WCLK => \N__65641\,
            WE => \N__39314\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65665\,
            RE => \N__39296\,
            WCLKE => \N__24891\,
            WCLK => \N__65666\,
            WE => \N__39305\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65524\,
            RE => \N__39401\,
            WCLKE => \N__23739\,
            WCLK => \N__65525\,
            WE => \N__39396\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65515\,
            RE => \N__39402\,
            WCLKE => \N__23732\,
            WCLK => \N__65516\,
            WE => \N__39400\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65614\,
            RE => \N__39336\,
            WCLKE => \N__24549\,
            WCLK => \N__65615\,
            WE => \N__39350\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65544\,
            RE => \N__39392\,
            WCLKE => \N__26637\,
            WCLK => \N__65545\,
            WE => \N__39381\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.mem_mem_0_0_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65594\,
            RE => \N__39362\,
            WCLKE => \N__24548\,
            WCLK => \N__65593\,
            WE => \N__39373\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical\ : SB_RAM40_4K
    generic map (
            WRITE_MODE => 0,
            READ_MODE => 0,
            INIT_0 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_8 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_9 => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_A => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_B => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_C => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_D => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_E => x"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_F => x"0000000000000000000000000000000000000000000000000000000000000000"
        )
    port map (
            RDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RDATA_wire\,
            RADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_RADDR_wire\,
            WADDR => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_WADDR_wire\,
            MASK => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_MASK_wire\,
            WDATA => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.mem_mem_0_1_physical_WDATA_wire\,
            RCLKE => 'H',
            RCLK => \N__65569\,
            RE => \N__39382\,
            WCLKE => \N__26636\,
            WCLK => \N__65570\,
            WE => \N__39374\
        );

    \next_sequence_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67138\,
            DIN => \N__67137\,
            DOUT => \N__67136\,
            PACKAGEPIN => next_sequence_wire
        );

    \next_sequence_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67138\,
            PADOUT => \N__67137\,
            PADIN => \N__67136\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__31524\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \stop_fpga2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67129\,
            DIN => \N__67128\,
            DOUT => \N__67127\,
            PACKAGEPIN => stop_fpga2_wire
        );

    \stop_fpga2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67129\,
            PADOUT => \N__67128\,
            PADIN => \N__67127\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__33015\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \stop1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67120\,
            DIN => \N__67119\,
            DOUT => \N__67118\,
            PACKAGEPIN => stop1_wire
        );

    \stop1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67120\,
            PADOUT => \N__67119\,
            PADIN => \N__67118\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67111\,
            DIN => \N__67110\,
            DOUT => \N__67109\,
            PACKAGEPIN => s0_wire
        );

    \s0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67111\,
            PADOUT => \N__67110\,
            PADIN => \N__67109\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \mcu_data_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67102\,
            DIN => \N__67101\,
            DOUT => \N__67100\,
            PACKAGEPIN => mcu_data_wire
        );

    \mcu_data_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67102\,
            PADOUT => \N__67101\,
            PADIN => \N__67100\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22536\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67093\,
            DIN => \N__67092\,
            DOUT => \N__67091\,
            PACKAGEPIN => start1_wire
        );

    \start1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67093\,
            PADOUT => \N__67092\,
            PADIN => \N__67091\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \rst_n_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67084\,
            DIN => \N__67083\,
            DOUT => \N__67082\,
            PACKAGEPIN => rst_n_wire
        );

    \rst_n_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__67084\,
            PADOUT => \N__67083\,
            PADIN => \N__67082\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => rst_n_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \scl_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67075\,
            DIN => \N__67074\,
            DOUT => \N__67073\,
            PACKAGEPIN => scl_wire
        );

    \scl_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__67075\,
            PADOUT => \N__67074\,
            PADIN => \N__67073\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => scl_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67066\,
            DIN => \N__67065\,
            DOUT => \N__67064\,
            PACKAGEPIN => dout0_wire
        );

    \dout0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67066\,
            PADOUT => \N__67065\,
            PADIN => \N__67064\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23139\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \stop0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67057\,
            DIN => \N__67056\,
            DOUT => \N__67055\,
            PACKAGEPIN => stop0_wire
        );

    \stop0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67057\,
            PADOUT => \N__67056\,
            PADIN => \N__67055\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s2_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67048\,
            DIN => \N__67047\,
            DOUT => \N__67046\,
            PACKAGEPIN => s2_wire
        );

    \s2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67048\,
            PADOUT => \N__67047\,
            PADIN => \N__67046\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24840\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \mcu_sclk_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67039\,
            DIN => \N__67038\,
            DOUT => \N__67037\,
            PACKAGEPIN => mcu_sclk_wire
        );

    \mcu_sclk_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67039\,
            PADOUT => \N__67038\,
            PADIN => \N__67037\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22359\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \frame_sync_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67030\,
            DIN => \N__67029\,
            DOUT => \N__67028\,
            PACKAGEPIN => frame_sync_wire
        );

    \frame_sync_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67030\,
            PADOUT => \N__67029\,
            PADIN => \N__67028\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sdin0_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67021\,
            DIN => \N__67020\,
            DOUT => \N__67019\,
            PACKAGEPIN => sdin0_wire
        );

    \sdin0_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__67021\,
            PADOUT => \N__67020\,
            PADIN => \N__67019\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sdin0_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sdin1_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67012\,
            DIN => \N__67011\,
            DOUT => \N__67010\,
            PACKAGEPIN => sdin1_wire
        );

    \sdin1_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__67012\,
            PADOUT => \N__67011\,
            PADIN => \N__67010\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sdin1_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \dout1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__67003\,
            DIN => \N__67002\,
            DOUT => \N__67001\,
            PACKAGEPIN => dout1_wire
        );

    \dout1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__67003\,
            PADOUT => \N__67002\,
            PADIN => \N__67001\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23265\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \csb1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66994\,
            DIN => \N__66993\,
            DOUT => \N__66992\,
            PACKAGEPIN => csb1_wire
        );

    \csb1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66994\,
            PADOUT => \N__66993\,
            PADIN => \N__66992\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__25653\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sclk1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66985\,
            DIN => \N__66984\,
            DOUT => \N__66983\,
            PACKAGEPIN => sclk1_wire
        );

    \sclk1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66985\,
            PADOUT => \N__66984\,
            PADIN => \N__66983\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22899\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sclk0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66976\,
            DIN => \N__66975\,
            DOUT => \N__66974\,
            PACKAGEPIN => sclk0_wire
        );

    \sclk0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66976\,
            PADOUT => \N__66975\,
            PADIN => \N__66974\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__22593\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s1_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66967\,
            DIN => \N__66966\,
            DOUT => \N__66965\,
            PACKAGEPIN => s1_wire
        );

    \s1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66967\,
            PADOUT => \N__66966\,
            PADIN => \N__66965\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__24836\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \enable_config_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66958\,
            DIN => \N__66957\,
            DOUT => \N__66956\,
            PACKAGEPIN => enable_config_wire
        );

    \enable_config_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66958\,
            PADOUT => \N__66957\,
            PADIN => \N__66956\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37449\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \sync_50hz_ibuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66949\,
            DIN => \N__66948\,
            DOUT => \N__66947\,
            PACKAGEPIN => sync_50hz_wire
        );

    \sync_50hz_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__66949\,
            PADOUT => \N__66948\,
            PADIN => \N__66947\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => sync_50hz_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \serial_out_testing_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66940\,
            DIN => \N__66939\,
            DOUT => \N__66938\,
            PACKAGEPIN => serial_out_testing_wire
        );

    \serial_out_testing_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66940\,
            PADOUT => \N__66939\,
            PADIN => \N__66938\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__35508\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \start0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66931\,
            DIN => \N__66930\,
            DOUT => \N__66929\,
            PACKAGEPIN => start0_wire
        );

    \start0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66931\,
            PADOUT => \N__66930\,
            PADIN => \N__66929\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \s3_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66922\,
            DIN => \N__66921\,
            DOUT => \N__66920\,
            PACKAGEPIN => s3_wire
        );

    \s3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66922\,
            PADOUT => \N__66921\,
            PADIN => \N__66920\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \elec_config_out_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66913\,
            DIN => \N__66912\,
            DOUT => \N__66911\,
            PACKAGEPIN => elec_config_out_wire
        );

    \elec_config_out_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66913\,
            PADOUT => \N__66912\,
            PADIN => \N__66911\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__37437\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \csb0_obuf_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66904\,
            DIN => \N__66903\,
            DOUT => \N__66902\,
            PACKAGEPIN => csb0_wire
        );

    \csb0_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__66904\,
            PADOUT => \N__66903\,
            PADIN => \N__66902\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__23064\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \IO_PIN_INST_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66895\,
            DIN => \N__66894\,
            DOUT => \N__66893\,
            PACKAGEPIN => sda
        );

    \IO_PIN_INST_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "101001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__66895\,
            PADOUT => \N__66894\,
            PADIN => \N__66893\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => \N__29340\,
            DIN0 => s_sda_i,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clock_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__66886\,
            DIN => \N__66885\,
            DOUT => \N__66884\,
            PACKAGEPIN => clock_wire
        );

    \clock_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__66886\,
            PADOUT => \N__66885\,
            PADIN => \N__66884\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clock_ibuf_gb_io_gb_input,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__16711\ : InMux
    port map (
            O => \N__66867\,
            I => \N__66863\
        );

    \I__16710\ : InMux
    port map (
            O => \N__66866\,
            I => \N__66860\
        );

    \I__16709\ : LocalMux
    port map (
            O => \N__66863\,
            I => \N__66857\
        );

    \I__16708\ : LocalMux
    port map (
            O => \N__66860\,
            I => \N__66854\
        );

    \I__16707\ : Span4Mux_h
    port map (
            O => \N__66857\,
            I => \N__66847\
        );

    \I__16706\ : Span4Mux_v
    port map (
            O => \N__66854\,
            I => \N__66844\
        );

    \I__16705\ : InMux
    port map (
            O => \N__66853\,
            I => \N__66839\
        );

    \I__16704\ : InMux
    port map (
            O => \N__66852\,
            I => \N__66839\
        );

    \I__16703\ : InMux
    port map (
            O => \N__66851\,
            I => \N__66834\
        );

    \I__16702\ : InMux
    port map (
            O => \N__66850\,
            I => \N__66834\
        );

    \I__16701\ : Odrv4
    port map (
            O => \N__66847\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0\
        );

    \I__16700\ : Odrv4
    port map (
            O => \N__66844\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0\
        );

    \I__16699\ : LocalMux
    port map (
            O => \N__66839\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0\
        );

    \I__16698\ : LocalMux
    port map (
            O => \N__66834\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0\
        );

    \I__16697\ : CascadeMux
    port map (
            O => \N__66825\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0_cascade_\
        );

    \I__16696\ : CascadeMux
    port map (
            O => \N__66822\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_0_2_cascade_\
        );

    \I__16695\ : CascadeMux
    port map (
            O => \N__66819\,
            I => \N__66816\
        );

    \I__16694\ : InMux
    port map (
            O => \N__66816\,
            I => \N__66806\
        );

    \I__16693\ : InMux
    port map (
            O => \N__66815\,
            I => \N__66806\
        );

    \I__16692\ : InMux
    port map (
            O => \N__66814\,
            I => \N__66806\
        );

    \I__16691\ : CascadeMux
    port map (
            O => \N__66813\,
            I => \N__66803\
        );

    \I__16690\ : LocalMux
    port map (
            O => \N__66806\,
            I => \N__66800\
        );

    \I__16689\ : InMux
    port map (
            O => \N__66803\,
            I => \N__66795\
        );

    \I__16688\ : Span4Mux_v
    port map (
            O => \N__66800\,
            I => \N__66791\
        );

    \I__16687\ : InMux
    port map (
            O => \N__66799\,
            I => \N__66784\
        );

    \I__16686\ : InMux
    port map (
            O => \N__66798\,
            I => \N__66781\
        );

    \I__16685\ : LocalMux
    port map (
            O => \N__66795\,
            I => \N__66776\
        );

    \I__16684\ : InMux
    port map (
            O => \N__66794\,
            I => \N__66773\
        );

    \I__16683\ : Span4Mux_v
    port map (
            O => \N__66791\,
            I => \N__66770\
        );

    \I__16682\ : InMux
    port map (
            O => \N__66790\,
            I => \N__66764\
        );

    \I__16681\ : InMux
    port map (
            O => \N__66789\,
            I => \N__66764\
        );

    \I__16680\ : InMux
    port map (
            O => \N__66788\,
            I => \N__66759\
        );

    \I__16679\ : InMux
    port map (
            O => \N__66787\,
            I => \N__66759\
        );

    \I__16678\ : LocalMux
    port map (
            O => \N__66784\,
            I => \N__66756\
        );

    \I__16677\ : LocalMux
    port map (
            O => \N__66781\,
            I => \N__66752\
        );

    \I__16676\ : InMux
    port map (
            O => \N__66780\,
            I => \N__66747\
        );

    \I__16675\ : InMux
    port map (
            O => \N__66779\,
            I => \N__66747\
        );

    \I__16674\ : Span4Mux_v
    port map (
            O => \N__66776\,
            I => \N__66744\
        );

    \I__16673\ : LocalMux
    port map (
            O => \N__66773\,
            I => \N__66739\
        );

    \I__16672\ : Span4Mux_h
    port map (
            O => \N__66770\,
            I => \N__66739\
        );

    \I__16671\ : InMux
    port map (
            O => \N__66769\,
            I => \N__66736\
        );

    \I__16670\ : LocalMux
    port map (
            O => \N__66764\,
            I => \N__66731\
        );

    \I__16669\ : LocalMux
    port map (
            O => \N__66759\,
            I => \N__66731\
        );

    \I__16668\ : Span4Mux_h
    port map (
            O => \N__66756\,
            I => \N__66728\
        );

    \I__16667\ : InMux
    port map (
            O => \N__66755\,
            I => \N__66725\
        );

    \I__16666\ : Span4Mux_h
    port map (
            O => \N__66752\,
            I => \N__66720\
        );

    \I__16665\ : LocalMux
    port map (
            O => \N__66747\,
            I => \N__66720\
        );

    \I__16664\ : Span4Mux_h
    port map (
            O => \N__66744\,
            I => \N__66715\
        );

    \I__16663\ : Span4Mux_h
    port map (
            O => \N__66739\,
            I => \N__66715\
        );

    \I__16662\ : LocalMux
    port map (
            O => \N__66736\,
            I => \N__66708\
        );

    \I__16661\ : Span4Mux_v
    port map (
            O => \N__66731\,
            I => \N__66708\
        );

    \I__16660\ : Span4Mux_v
    port map (
            O => \N__66728\,
            I => \N__66708\
        );

    \I__16659\ : LocalMux
    port map (
            O => \N__66725\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8\
        );

    \I__16658\ : Odrv4
    port map (
            O => \N__66720\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8\
        );

    \I__16657\ : Odrv4
    port map (
            O => \N__66715\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8\
        );

    \I__16656\ : Odrv4
    port map (
            O => \N__66708\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8\
        );

    \I__16655\ : InMux
    port map (
            O => \N__66699\,
            I => \N__66696\
        );

    \I__16654\ : LocalMux
    port map (
            O => \N__66696\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_2\
        );

    \I__16653\ : CascadeMux
    port map (
            O => \N__66693\,
            I => \N__66688\
        );

    \I__16652\ : InMux
    port map (
            O => \N__66692\,
            I => \N__66684\
        );

    \I__16651\ : InMux
    port map (
            O => \N__66691\,
            I => \N__66681\
        );

    \I__16650\ : InMux
    port map (
            O => \N__66688\,
            I => \N__66677\
        );

    \I__16649\ : InMux
    port map (
            O => \N__66687\,
            I => \N__66670\
        );

    \I__16648\ : LocalMux
    port map (
            O => \N__66684\,
            I => \N__66665\
        );

    \I__16647\ : LocalMux
    port map (
            O => \N__66681\,
            I => \N__66665\
        );

    \I__16646\ : InMux
    port map (
            O => \N__66680\,
            I => \N__66662\
        );

    \I__16645\ : LocalMux
    port map (
            O => \N__66677\,
            I => \N__66659\
        );

    \I__16644\ : CascadeMux
    port map (
            O => \N__66676\,
            I => \N__66655\
        );

    \I__16643\ : InMux
    port map (
            O => \N__66675\,
            I => \N__66650\
        );

    \I__16642\ : InMux
    port map (
            O => \N__66674\,
            I => \N__66645\
        );

    \I__16641\ : InMux
    port map (
            O => \N__66673\,
            I => \N__66645\
        );

    \I__16640\ : LocalMux
    port map (
            O => \N__66670\,
            I => \N__66640\
        );

    \I__16639\ : Span4Mux_v
    port map (
            O => \N__66665\,
            I => \N__66640\
        );

    \I__16638\ : LocalMux
    port map (
            O => \N__66662\,
            I => \N__66637\
        );

    \I__16637\ : Span4Mux_h
    port map (
            O => \N__66659\,
            I => \N__66634\
        );

    \I__16636\ : InMux
    port map (
            O => \N__66658\,
            I => \N__66627\
        );

    \I__16635\ : InMux
    port map (
            O => \N__66655\,
            I => \N__66627\
        );

    \I__16634\ : InMux
    port map (
            O => \N__66654\,
            I => \N__66627\
        );

    \I__16633\ : InMux
    port map (
            O => \N__66653\,
            I => \N__66624\
        );

    \I__16632\ : LocalMux
    port map (
            O => \N__66650\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16631\ : LocalMux
    port map (
            O => \N__66645\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16630\ : Odrv4
    port map (
            O => \N__66640\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16629\ : Odrv12
    port map (
            O => \N__66637\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16628\ : Odrv4
    port map (
            O => \N__66634\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16627\ : LocalMux
    port map (
            O => \N__66627\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16626\ : LocalMux
    port map (
            O => \N__66624\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\
        );

    \I__16625\ : CascadeMux
    port map (
            O => \N__66609\,
            I => \N__66604\
        );

    \I__16624\ : InMux
    port map (
            O => \N__66608\,
            I => \N__66599\
        );

    \I__16623\ : InMux
    port map (
            O => \N__66607\,
            I => \N__66594\
        );

    \I__16622\ : InMux
    port map (
            O => \N__66604\,
            I => \N__66594\
        );

    \I__16621\ : InMux
    port map (
            O => \N__66603\,
            I => \N__66590\
        );

    \I__16620\ : InMux
    port map (
            O => \N__66602\,
            I => \N__66587\
        );

    \I__16619\ : LocalMux
    port map (
            O => \N__66599\,
            I => \N__66582\
        );

    \I__16618\ : LocalMux
    port map (
            O => \N__66594\,
            I => \N__66582\
        );

    \I__16617\ : InMux
    port map (
            O => \N__66593\,
            I => \N__66579\
        );

    \I__16616\ : LocalMux
    port map (
            O => \N__66590\,
            I => \N__66574\
        );

    \I__16615\ : LocalMux
    port map (
            O => \N__66587\,
            I => \N__66574\
        );

    \I__16614\ : Span4Mux_h
    port map (
            O => \N__66582\,
            I => \N__66571\
        );

    \I__16613\ : LocalMux
    port map (
            O => \N__66579\,
            I => \N__66568\
        );

    \I__16612\ : Odrv4
    port map (
            O => \N__66574\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0\
        );

    \I__16611\ : Odrv4
    port map (
            O => \N__66571\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0\
        );

    \I__16610\ : Odrv12
    port map (
            O => \N__66568\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0\
        );

    \I__16609\ : InMux
    port map (
            O => \N__66561\,
            I => \N__66556\
        );

    \I__16608\ : InMux
    port map (
            O => \N__66560\,
            I => \N__66545\
        );

    \I__16607\ : InMux
    port map (
            O => \N__66559\,
            I => \N__66542\
        );

    \I__16606\ : LocalMux
    port map (
            O => \N__66556\,
            I => \N__66539\
        );

    \I__16605\ : InMux
    port map (
            O => \N__66555\,
            I => \N__66536\
        );

    \I__16604\ : InMux
    port map (
            O => \N__66554\,
            I => \N__66533\
        );

    \I__16603\ : InMux
    port map (
            O => \N__66553\,
            I => \N__66522\
        );

    \I__16602\ : InMux
    port map (
            O => \N__66552\,
            I => \N__66522\
        );

    \I__16601\ : InMux
    port map (
            O => \N__66551\,
            I => \N__66522\
        );

    \I__16600\ : InMux
    port map (
            O => \N__66550\,
            I => \N__66522\
        );

    \I__16599\ : InMux
    port map (
            O => \N__66549\,
            I => \N__66522\
        );

    \I__16598\ : InMux
    port map (
            O => \N__66548\,
            I => \N__66519\
        );

    \I__16597\ : LocalMux
    port map (
            O => \N__66545\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16596\ : LocalMux
    port map (
            O => \N__66542\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16595\ : Odrv4
    port map (
            O => \N__66539\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16594\ : LocalMux
    port map (
            O => \N__66536\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16593\ : LocalMux
    port map (
            O => \N__66533\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16592\ : LocalMux
    port map (
            O => \N__66522\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16591\ : LocalMux
    port map (
            O => \N__66519\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\
        );

    \I__16590\ : InMux
    port map (
            O => \N__66504\,
            I => \N__66499\
        );

    \I__16589\ : InMux
    port map (
            O => \N__66503\,
            I => \N__66489\
        );

    \I__16588\ : InMux
    port map (
            O => \N__66502\,
            I => \N__66486\
        );

    \I__16587\ : LocalMux
    port map (
            O => \N__66499\,
            I => \N__66483\
        );

    \I__16586\ : InMux
    port map (
            O => \N__66498\,
            I => \N__66478\
        );

    \I__16585\ : InMux
    port map (
            O => \N__66497\,
            I => \N__66478\
        );

    \I__16584\ : InMux
    port map (
            O => \N__66496\,
            I => \N__66471\
        );

    \I__16583\ : InMux
    port map (
            O => \N__66495\,
            I => \N__66471\
        );

    \I__16582\ : InMux
    port map (
            O => \N__66494\,
            I => \N__66471\
        );

    \I__16581\ : InMux
    port map (
            O => \N__66493\,
            I => \N__66466\
        );

    \I__16580\ : InMux
    port map (
            O => \N__66492\,
            I => \N__66466\
        );

    \I__16579\ : LocalMux
    port map (
            O => \N__66489\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\
        );

    \I__16578\ : LocalMux
    port map (
            O => \N__66486\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\
        );

    \I__16577\ : Odrv4
    port map (
            O => \N__66483\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\
        );

    \I__16576\ : LocalMux
    port map (
            O => \N__66478\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\
        );

    \I__16575\ : LocalMux
    port map (
            O => \N__66471\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\
        );

    \I__16574\ : LocalMux
    port map (
            O => \N__66466\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\
        );

    \I__16573\ : InMux
    port map (
            O => \N__66453\,
            I => \N__66450\
        );

    \I__16572\ : LocalMux
    port map (
            O => \N__66450\,
            I => \N__66446\
        );

    \I__16571\ : CascadeMux
    port map (
            O => \N__66449\,
            I => \N__66443\
        );

    \I__16570\ : Span4Mux_v
    port map (
            O => \N__66446\,
            I => \N__66440\
        );

    \I__16569\ : InMux
    port map (
            O => \N__66443\,
            I => \N__66437\
        );

    \I__16568\ : Span4Mux_v
    port map (
            O => \N__66440\,
            I => \N__66432\
        );

    \I__16567\ : LocalMux
    port map (
            O => \N__66437\,
            I => \N__66432\
        );

    \I__16566\ : Span4Mux_v
    port map (
            O => \N__66432\,
            I => \N__66428\
        );

    \I__16565\ : InMux
    port map (
            O => \N__66431\,
            I => \N__66425\
        );

    \I__16564\ : Odrv4
    port map (
            O => \N__66428\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0\
        );

    \I__16563\ : LocalMux
    port map (
            O => \N__66425\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0\
        );

    \I__16562\ : InMux
    port map (
            O => \N__66420\,
            I => \N__66416\
        );

    \I__16561\ : CascadeMux
    port map (
            O => \N__66419\,
            I => \N__66413\
        );

    \I__16560\ : LocalMux
    port map (
            O => \N__66416\,
            I => \N__66407\
        );

    \I__16559\ : InMux
    port map (
            O => \N__66413\,
            I => \N__66402\
        );

    \I__16558\ : InMux
    port map (
            O => \N__66412\,
            I => \N__66402\
        );

    \I__16557\ : InMux
    port map (
            O => \N__66411\,
            I => \N__66397\
        );

    \I__16556\ : InMux
    port map (
            O => \N__66410\,
            I => \N__66397\
        );

    \I__16555\ : Span4Mux_v
    port map (
            O => \N__66407\,
            I => \N__66394\
        );

    \I__16554\ : LocalMux
    port map (
            O => \N__66402\,
            I => \N__66389\
        );

    \I__16553\ : LocalMux
    port map (
            O => \N__66397\,
            I => \N__66389\
        );

    \I__16552\ : Odrv4
    port map (
            O => \N__66394\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0\
        );

    \I__16551\ : Odrv4
    port map (
            O => \N__66389\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0\
        );

    \I__16550\ : InMux
    port map (
            O => \N__66384\,
            I => \N__66379\
        );

    \I__16549\ : InMux
    port map (
            O => \N__66383\,
            I => \N__66370\
        );

    \I__16548\ : InMux
    port map (
            O => \N__66382\,
            I => \N__66370\
        );

    \I__16547\ : LocalMux
    port map (
            O => \N__66379\,
            I => \N__66367\
        );

    \I__16546\ : InMux
    port map (
            O => \N__66378\,
            I => \N__66364\
        );

    \I__16545\ : InMux
    port map (
            O => \N__66377\,
            I => \N__66361\
        );

    \I__16544\ : InMux
    port map (
            O => \N__66376\,
            I => \N__66356\
        );

    \I__16543\ : InMux
    port map (
            O => \N__66375\,
            I => \N__66356\
        );

    \I__16542\ : LocalMux
    port map (
            O => \N__66370\,
            I => \N__66353\
        );

    \I__16541\ : Span4Mux_h
    port map (
            O => \N__66367\,
            I => \N__66346\
        );

    \I__16540\ : LocalMux
    port map (
            O => \N__66364\,
            I => \N__66346\
        );

    \I__16539\ : LocalMux
    port map (
            O => \N__66361\,
            I => \N__66346\
        );

    \I__16538\ : LocalMux
    port map (
            O => \N__66356\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0\
        );

    \I__16537\ : Odrv12
    port map (
            O => \N__66353\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0\
        );

    \I__16536\ : Odrv4
    port map (
            O => \N__66346\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0\
        );

    \I__16535\ : InMux
    port map (
            O => \N__66339\,
            I => \N__66336\
        );

    \I__16534\ : LocalMux
    port map (
            O => \N__66336\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666_2\
        );

    \I__16533\ : CascadeMux
    port map (
            O => \N__66333\,
            I => \N__66330\
        );

    \I__16532\ : InMux
    port map (
            O => \N__66330\,
            I => \N__66321\
        );

    \I__16531\ : InMux
    port map (
            O => \N__66329\,
            I => \N__66312\
        );

    \I__16530\ : InMux
    port map (
            O => \N__66328\,
            I => \N__66312\
        );

    \I__16529\ : InMux
    port map (
            O => \N__66327\,
            I => \N__66312\
        );

    \I__16528\ : InMux
    port map (
            O => \N__66326\,
            I => \N__66312\
        );

    \I__16527\ : InMux
    port map (
            O => \N__66325\,
            I => \N__66309\
        );

    \I__16526\ : InMux
    port map (
            O => \N__66324\,
            I => \N__66306\
        );

    \I__16525\ : LocalMux
    port map (
            O => \N__66321\,
            I => \N__66303\
        );

    \I__16524\ : LocalMux
    port map (
            O => \N__66312\,
            I => \N__66300\
        );

    \I__16523\ : LocalMux
    port map (
            O => \N__66309\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17\
        );

    \I__16522\ : LocalMux
    port map (
            O => \N__66306\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17\
        );

    \I__16521\ : Odrv12
    port map (
            O => \N__66303\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17\
        );

    \I__16520\ : Odrv4
    port map (
            O => \N__66300\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17\
        );

    \I__16519\ : InMux
    port map (
            O => \N__66291\,
            I => \N__66287\
        );

    \I__16518\ : InMux
    port map (
            O => \N__66290\,
            I => \N__66284\
        );

    \I__16517\ : LocalMux
    port map (
            O => \N__66287\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_295\
        );

    \I__16516\ : LocalMux
    port map (
            O => \N__66284\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_295\
        );

    \I__16515\ : CascadeMux
    port map (
            O => \N__66279\,
            I => \N_73_i_0_cascade_\
        );

    \I__16514\ : InMux
    port map (
            O => \N__66276\,
            I => \N__66268\
        );

    \I__16513\ : InMux
    port map (
            O => \N__66275\,
            I => \N__66268\
        );

    \I__16512\ : InMux
    port map (
            O => \N__66274\,
            I => \N__66265\
        );

    \I__16511\ : InMux
    port map (
            O => \N__66273\,
            I => \N__66261\
        );

    \I__16510\ : LocalMux
    port map (
            O => \N__66268\,
            I => \N__66256\
        );

    \I__16509\ : LocalMux
    port map (
            O => \N__66265\,
            I => \N__66256\
        );

    \I__16508\ : InMux
    port map (
            O => \N__66264\,
            I => \N__66252\
        );

    \I__16507\ : LocalMux
    port map (
            O => \N__66261\,
            I => \N__66248\
        );

    \I__16506\ : Span4Mux_v
    port map (
            O => \N__66256\,
            I => \N__66245\
        );

    \I__16505\ : InMux
    port map (
            O => \N__66255\,
            I => \N__66240\
        );

    \I__16504\ : LocalMux
    port map (
            O => \N__66252\,
            I => \N__66237\
        );

    \I__16503\ : InMux
    port map (
            O => \N__66251\,
            I => \N__66234\
        );

    \I__16502\ : Span4Mux_v
    port map (
            O => \N__66248\,
            I => \N__66229\
        );

    \I__16501\ : Span4Mux_h
    port map (
            O => \N__66245\,
            I => \N__66229\
        );

    \I__16500\ : InMux
    port map (
            O => \N__66244\,
            I => \N__66226\
        );

    \I__16499\ : InMux
    port map (
            O => \N__66243\,
            I => \N__66223\
        );

    \I__16498\ : LocalMux
    port map (
            O => \N__66240\,
            I => \N__66220\
        );

    \I__16497\ : Span4Mux_h
    port map (
            O => \N__66237\,
            I => \N__66215\
        );

    \I__16496\ : LocalMux
    port map (
            O => \N__66234\,
            I => \N__66215\
        );

    \I__16495\ : Span4Mux_h
    port map (
            O => \N__66229\,
            I => \N__66210\
        );

    \I__16494\ : LocalMux
    port map (
            O => \N__66226\,
            I => \N__66210\
        );

    \I__16493\ : LocalMux
    port map (
            O => \N__66223\,
            I => \I2C_top_level_inst1_s_burst\
        );

    \I__16492\ : Odrv12
    port map (
            O => \N__66220\,
            I => \I2C_top_level_inst1_s_burst\
        );

    \I__16491\ : Odrv4
    port map (
            O => \N__66215\,
            I => \I2C_top_level_inst1_s_burst\
        );

    \I__16490\ : Odrv4
    port map (
            O => \N__66210\,
            I => \I2C_top_level_inst1_s_burst\
        );

    \I__16489\ : InMux
    port map (
            O => \N__66201\,
            I => \N__66198\
        );

    \I__16488\ : LocalMux
    port map (
            O => \N__66198\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_19\
        );

    \I__16487\ : CascadeMux
    port map (
            O => \N__66195\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_274_cascade_\
        );

    \I__16486\ : CascadeMux
    port map (
            O => \N__66192\,
            I => \N__66188\
        );

    \I__16485\ : InMux
    port map (
            O => \N__66191\,
            I => \N__66175\
        );

    \I__16484\ : InMux
    port map (
            O => \N__66188\,
            I => \N__66175\
        );

    \I__16483\ : InMux
    port map (
            O => \N__66187\,
            I => \N__66175\
        );

    \I__16482\ : InMux
    port map (
            O => \N__66186\,
            I => \N__66175\
        );

    \I__16481\ : InMux
    port map (
            O => \N__66185\,
            I => \N__66169\
        );

    \I__16480\ : InMux
    port map (
            O => \N__66184\,
            I => \N__66169\
        );

    \I__16479\ : LocalMux
    port map (
            O => \N__66175\,
            I => \N__66160\
        );

    \I__16478\ : InMux
    port map (
            O => \N__66174\,
            I => \N__66157\
        );

    \I__16477\ : LocalMux
    port map (
            O => \N__66169\,
            I => \N__66151\
        );

    \I__16476\ : InMux
    port map (
            O => \N__66168\,
            I => \N__66143\
        );

    \I__16475\ : InMux
    port map (
            O => \N__66167\,
            I => \N__66143\
        );

    \I__16474\ : InMux
    port map (
            O => \N__66166\,
            I => \N__66143\
        );

    \I__16473\ : InMux
    port map (
            O => \N__66165\,
            I => \N__66138\
        );

    \I__16472\ : InMux
    port map (
            O => \N__66164\,
            I => \N__66138\
        );

    \I__16471\ : InMux
    port map (
            O => \N__66163\,
            I => \N__66135\
        );

    \I__16470\ : Span4Mux_h
    port map (
            O => \N__66160\,
            I => \N__66130\
        );

    \I__16469\ : LocalMux
    port map (
            O => \N__66157\,
            I => \N__66130\
        );

    \I__16468\ : CascadeMux
    port map (
            O => \N__66156\,
            I => \N__66126\
        );

    \I__16467\ : CascadeMux
    port map (
            O => \N__66155\,
            I => \N__66122\
        );

    \I__16466\ : CascadeMux
    port map (
            O => \N__66154\,
            I => \N__66119\
        );

    \I__16465\ : Span4Mux_v
    port map (
            O => \N__66151\,
            I => \N__66115\
        );

    \I__16464\ : InMux
    port map (
            O => \N__66150\,
            I => \N__66112\
        );

    \I__16463\ : LocalMux
    port map (
            O => \N__66143\,
            I => \N__66106\
        );

    \I__16462\ : LocalMux
    port map (
            O => \N__66138\,
            I => \N__66102\
        );

    \I__16461\ : LocalMux
    port map (
            O => \N__66135\,
            I => \N__66099\
        );

    \I__16460\ : Span4Mux_h
    port map (
            O => \N__66130\,
            I => \N__66096\
        );

    \I__16459\ : InMux
    port map (
            O => \N__66129\,
            I => \N__66086\
        );

    \I__16458\ : InMux
    port map (
            O => \N__66126\,
            I => \N__66086\
        );

    \I__16457\ : InMux
    port map (
            O => \N__66125\,
            I => \N__66086\
        );

    \I__16456\ : InMux
    port map (
            O => \N__66122\,
            I => \N__66079\
        );

    \I__16455\ : InMux
    port map (
            O => \N__66119\,
            I => \N__66079\
        );

    \I__16454\ : InMux
    port map (
            O => \N__66118\,
            I => \N__66079\
        );

    \I__16453\ : Span4Mux_v
    port map (
            O => \N__66115\,
            I => \N__66074\
        );

    \I__16452\ : LocalMux
    port map (
            O => \N__66112\,
            I => \N__66074\
        );

    \I__16451\ : InMux
    port map (
            O => \N__66111\,
            I => \N__66067\
        );

    \I__16450\ : InMux
    port map (
            O => \N__66110\,
            I => \N__66067\
        );

    \I__16449\ : InMux
    port map (
            O => \N__66109\,
            I => \N__66067\
        );

    \I__16448\ : Span4Mux_v
    port map (
            O => \N__66106\,
            I => \N__66064\
        );

    \I__16447\ : InMux
    port map (
            O => \N__66105\,
            I => \N__66061\
        );

    \I__16446\ : Span4Mux_h
    port map (
            O => \N__66102\,
            I => \N__66054\
        );

    \I__16445\ : Span4Mux_h
    port map (
            O => \N__66099\,
            I => \N__66054\
        );

    \I__16444\ : Span4Mux_v
    port map (
            O => \N__66096\,
            I => \N__66054\
        );

    \I__16443\ : InMux
    port map (
            O => \N__66095\,
            I => \N__66051\
        );

    \I__16442\ : InMux
    port map (
            O => \N__66094\,
            I => \N__66046\
        );

    \I__16441\ : InMux
    port map (
            O => \N__66093\,
            I => \N__66046\
        );

    \I__16440\ : LocalMux
    port map (
            O => \N__66086\,
            I => \N__66041\
        );

    \I__16439\ : LocalMux
    port map (
            O => \N__66079\,
            I => \N__66041\
        );

    \I__16438\ : Span4Mux_h
    port map (
            O => \N__66074\,
            I => \N__66038\
        );

    \I__16437\ : LocalMux
    port map (
            O => \N__66067\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16436\ : Odrv4
    port map (
            O => \N__66064\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16435\ : LocalMux
    port map (
            O => \N__66061\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16434\ : Odrv4
    port map (
            O => \N__66054\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16433\ : LocalMux
    port map (
            O => \N__66051\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16432\ : LocalMux
    port map (
            O => \N__66046\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16431\ : Odrv4
    port map (
            O => \N__66041\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16430\ : Odrv4
    port map (
            O => \N__66038\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\
        );

    \I__16429\ : InMux
    port map (
            O => \N__66021\,
            I => \N__66012\
        );

    \I__16428\ : InMux
    port map (
            O => \N__66020\,
            I => \N__66012\
        );

    \I__16427\ : InMux
    port map (
            O => \N__66019\,
            I => \N__66009\
        );

    \I__16426\ : InMux
    port map (
            O => \N__66018\,
            I => \N__66006\
        );

    \I__16425\ : InMux
    port map (
            O => \N__66017\,
            I => \N__66003\
        );

    \I__16424\ : LocalMux
    port map (
            O => \N__66012\,
            I => \N__65998\
        );

    \I__16423\ : LocalMux
    port map (
            O => \N__66009\,
            I => \N__65998\
        );

    \I__16422\ : LocalMux
    port map (
            O => \N__66006\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19\
        );

    \I__16421\ : LocalMux
    port map (
            O => \N__66003\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19\
        );

    \I__16420\ : Odrv4
    port map (
            O => \N__65998\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19\
        );

    \I__16419\ : InMux
    port map (
            O => \N__65991\,
            I => \N__65988\
        );

    \I__16418\ : LocalMux
    port map (
            O => \N__65988\,
            I => \N__65982\
        );

    \I__16417\ : CascadeMux
    port map (
            O => \N__65987\,
            I => \N__65979\
        );

    \I__16416\ : CascadeMux
    port map (
            O => \N__65986\,
            I => \N__65975\
        );

    \I__16415\ : InMux
    port map (
            O => \N__65985\,
            I => \N__65971\
        );

    \I__16414\ : Span4Mux_v
    port map (
            O => \N__65982\,
            I => \N__65968\
        );

    \I__16413\ : InMux
    port map (
            O => \N__65979\,
            I => \N__65965\
        );

    \I__16412\ : InMux
    port map (
            O => \N__65978\,
            I => \N__65962\
        );

    \I__16411\ : InMux
    port map (
            O => \N__65975\,
            I => \N__65957\
        );

    \I__16410\ : InMux
    port map (
            O => \N__65974\,
            I => \N__65957\
        );

    \I__16409\ : LocalMux
    port map (
            O => \N__65971\,
            I => \N__65946\
        );

    \I__16408\ : Sp12to4
    port map (
            O => \N__65968\,
            I => \N__65946\
        );

    \I__16407\ : LocalMux
    port map (
            O => \N__65965\,
            I => \N__65946\
        );

    \I__16406\ : LocalMux
    port map (
            O => \N__65962\,
            I => \N__65946\
        );

    \I__16405\ : LocalMux
    port map (
            O => \N__65957\,
            I => \N__65946\
        );

    \I__16404\ : Span12Mux_h
    port map (
            O => \N__65946\,
            I => \N__65942\
        );

    \I__16403\ : InMux
    port map (
            O => \N__65945\,
            I => \N__65939\
        );

    \I__16402\ : Odrv12
    port map (
            O => \N__65942\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6\
        );

    \I__16401\ : LocalMux
    port map (
            O => \N__65939\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6\
        );

    \I__16400\ : InMux
    port map (
            O => \N__65934\,
            I => \N__65927\
        );

    \I__16399\ : InMux
    port map (
            O => \N__65933\,
            I => \N__65927\
        );

    \I__16398\ : CascadeMux
    port map (
            O => \N__65932\,
            I => \N__65923\
        );

    \I__16397\ : LocalMux
    port map (
            O => \N__65927\,
            I => \N__65920\
        );

    \I__16396\ : InMux
    port map (
            O => \N__65926\,
            I => \N__65915\
        );

    \I__16395\ : InMux
    port map (
            O => \N__65923\,
            I => \N__65915\
        );

    \I__16394\ : Span4Mux_h
    port map (
            O => \N__65920\,
            I => \N__65909\
        );

    \I__16393\ : LocalMux
    port map (
            O => \N__65915\,
            I => \N__65909\
        );

    \I__16392\ : InMux
    port map (
            O => \N__65914\,
            I => \N__65906\
        );

    \I__16391\ : Span4Mux_h
    port map (
            O => \N__65909\,
            I => \N__65903\
        );

    \I__16390\ : LocalMux
    port map (
            O => \N__65906\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2\
        );

    \I__16389\ : Odrv4
    port map (
            O => \N__65903\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2\
        );

    \I__16388\ : CascadeMux
    port map (
            O => \N__65898\,
            I => \N__65894\
        );

    \I__16387\ : InMux
    port map (
            O => \N__65897\,
            I => \N__65889\
        );

    \I__16386\ : InMux
    port map (
            O => \N__65894\,
            I => \N__65884\
        );

    \I__16385\ : InMux
    port map (
            O => \N__65893\,
            I => \N__65884\
        );

    \I__16384\ : InMux
    port map (
            O => \N__65892\,
            I => \N__65881\
        );

    \I__16383\ : LocalMux
    port map (
            O => \N__65889\,
            I => \N__65878\
        );

    \I__16382\ : LocalMux
    port map (
            O => \N__65884\,
            I => \N__65873\
        );

    \I__16381\ : LocalMux
    port map (
            O => \N__65881\,
            I => \N__65873\
        );

    \I__16380\ : Span4Mux_v
    port map (
            O => \N__65878\,
            I => \N__65866\
        );

    \I__16379\ : Span4Mux_v
    port map (
            O => \N__65873\,
            I => \N__65866\
        );

    \I__16378\ : InMux
    port map (
            O => \N__65872\,
            I => \N__65861\
        );

    \I__16377\ : InMux
    port map (
            O => \N__65871\,
            I => \N__65861\
        );

    \I__16376\ : Odrv4
    port map (
            O => \N__65866\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2\
        );

    \I__16375\ : LocalMux
    port map (
            O => \N__65861\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2\
        );

    \I__16374\ : InMux
    port map (
            O => \N__65856\,
            I => \N__65853\
        );

    \I__16373\ : LocalMux
    port map (
            O => \N__65853\,
            I => \N__65849\
        );

    \I__16372\ : InMux
    port map (
            O => \N__65852\,
            I => \N__65845\
        );

    \I__16371\ : Span4Mux_v
    port map (
            O => \N__65849\,
            I => \N__65842\
        );

    \I__16370\ : InMux
    port map (
            O => \N__65848\,
            I => \N__65839\
        );

    \I__16369\ : LocalMux
    port map (
            O => \N__65845\,
            I => \N__65836\
        );

    \I__16368\ : Odrv4
    port map (
            O => \N__65842\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2\
        );

    \I__16367\ : LocalMux
    port map (
            O => \N__65839\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2\
        );

    \I__16366\ : Odrv4
    port map (
            O => \N__65836\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2\
        );

    \I__16365\ : InMux
    port map (
            O => \N__65829\,
            I => \N__65826\
        );

    \I__16364\ : LocalMux
    port map (
            O => \N__65826\,
            I => \N__65823\
        );

    \I__16363\ : Odrv4
    port map (
            O => \N__65823\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_276\
        );

    \I__16362\ : InMux
    port map (
            O => \N__65820\,
            I => \N__65816\
        );

    \I__16361\ : InMux
    port map (
            O => \N__65819\,
            I => \N__65813\
        );

    \I__16360\ : LocalMux
    port map (
            O => \N__65816\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1\
        );

    \I__16359\ : LocalMux
    port map (
            O => \N__65813\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1\
        );

    \I__16358\ : CascadeMux
    port map (
            O => \N__65808\,
            I => \N__65804\
        );

    \I__16357\ : CascadeMux
    port map (
            O => \N__65807\,
            I => \N__65801\
        );

    \I__16356\ : InMux
    port map (
            O => \N__65804\,
            I => \N__65797\
        );

    \I__16355\ : InMux
    port map (
            O => \N__65801\,
            I => \N__65792\
        );

    \I__16354\ : InMux
    port map (
            O => \N__65800\,
            I => \N__65792\
        );

    \I__16353\ : LocalMux
    port map (
            O => \N__65797\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_245\
        );

    \I__16352\ : LocalMux
    port map (
            O => \N__65792\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_245\
        );

    \I__16351\ : InMux
    port map (
            O => \N__65787\,
            I => \N__65784\
        );

    \I__16350\ : LocalMux
    port map (
            O => \N__65784\,
            I => \N__65780\
        );

    \I__16349\ : InMux
    port map (
            O => \N__65783\,
            I => \N__65777\
        );

    \I__16348\ : Odrv4
    port map (
            O => \N__65780\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0\
        );

    \I__16347\ : LocalMux
    port map (
            O => \N__65777\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0\
        );

    \I__16346\ : CascadeMux
    port map (
            O => \N__65772\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1669_cascade_\
        );

    \I__16345\ : InMux
    port map (
            O => \N__65769\,
            I => \N__65764\
        );

    \I__16344\ : InMux
    port map (
            O => \N__65768\,
            I => \N__65761\
        );

    \I__16343\ : InMux
    port map (
            O => \N__65767\,
            I => \N__65758\
        );

    \I__16342\ : LocalMux
    port map (
            O => \N__65764\,
            I => \N__65755\
        );

    \I__16341\ : LocalMux
    port map (
            O => \N__65761\,
            I => \N__65710\
        );

    \I__16340\ : LocalMux
    port map (
            O => \N__65758\,
            I => \N__65707\
        );

    \I__16339\ : Glb2LocalMux
    port map (
            O => \N__65755\,
            I => \N__65034\
        );

    \I__16338\ : ClkMux
    port map (
            O => \N__65754\,
            I => \N__65034\
        );

    \I__16337\ : ClkMux
    port map (
            O => \N__65753\,
            I => \N__65034\
        );

    \I__16336\ : ClkMux
    port map (
            O => \N__65752\,
            I => \N__65034\
        );

    \I__16335\ : ClkMux
    port map (
            O => \N__65751\,
            I => \N__65034\
        );

    \I__16334\ : ClkMux
    port map (
            O => \N__65750\,
            I => \N__65034\
        );

    \I__16333\ : ClkMux
    port map (
            O => \N__65749\,
            I => \N__65034\
        );

    \I__16332\ : ClkMux
    port map (
            O => \N__65748\,
            I => \N__65034\
        );

    \I__16331\ : ClkMux
    port map (
            O => \N__65747\,
            I => \N__65034\
        );

    \I__16330\ : ClkMux
    port map (
            O => \N__65746\,
            I => \N__65034\
        );

    \I__16329\ : ClkMux
    port map (
            O => \N__65745\,
            I => \N__65034\
        );

    \I__16328\ : ClkMux
    port map (
            O => \N__65744\,
            I => \N__65034\
        );

    \I__16327\ : ClkMux
    port map (
            O => \N__65743\,
            I => \N__65034\
        );

    \I__16326\ : ClkMux
    port map (
            O => \N__65742\,
            I => \N__65034\
        );

    \I__16325\ : ClkMux
    port map (
            O => \N__65741\,
            I => \N__65034\
        );

    \I__16324\ : ClkMux
    port map (
            O => \N__65740\,
            I => \N__65034\
        );

    \I__16323\ : ClkMux
    port map (
            O => \N__65739\,
            I => \N__65034\
        );

    \I__16322\ : ClkMux
    port map (
            O => \N__65738\,
            I => \N__65034\
        );

    \I__16321\ : ClkMux
    port map (
            O => \N__65737\,
            I => \N__65034\
        );

    \I__16320\ : ClkMux
    port map (
            O => \N__65736\,
            I => \N__65034\
        );

    \I__16319\ : ClkMux
    port map (
            O => \N__65735\,
            I => \N__65034\
        );

    \I__16318\ : ClkMux
    port map (
            O => \N__65734\,
            I => \N__65034\
        );

    \I__16317\ : ClkMux
    port map (
            O => \N__65733\,
            I => \N__65034\
        );

    \I__16316\ : ClkMux
    port map (
            O => \N__65732\,
            I => \N__65034\
        );

    \I__16315\ : ClkMux
    port map (
            O => \N__65731\,
            I => \N__65034\
        );

    \I__16314\ : ClkMux
    port map (
            O => \N__65730\,
            I => \N__65034\
        );

    \I__16313\ : ClkMux
    port map (
            O => \N__65729\,
            I => \N__65034\
        );

    \I__16312\ : ClkMux
    port map (
            O => \N__65728\,
            I => \N__65034\
        );

    \I__16311\ : ClkMux
    port map (
            O => \N__65727\,
            I => \N__65034\
        );

    \I__16310\ : ClkMux
    port map (
            O => \N__65726\,
            I => \N__65034\
        );

    \I__16309\ : ClkMux
    port map (
            O => \N__65725\,
            I => \N__65034\
        );

    \I__16308\ : ClkMux
    port map (
            O => \N__65724\,
            I => \N__65034\
        );

    \I__16307\ : ClkMux
    port map (
            O => \N__65723\,
            I => \N__65034\
        );

    \I__16306\ : ClkMux
    port map (
            O => \N__65722\,
            I => \N__65034\
        );

    \I__16305\ : ClkMux
    port map (
            O => \N__65721\,
            I => \N__65034\
        );

    \I__16304\ : ClkMux
    port map (
            O => \N__65720\,
            I => \N__65034\
        );

    \I__16303\ : ClkMux
    port map (
            O => \N__65719\,
            I => \N__65034\
        );

    \I__16302\ : ClkMux
    port map (
            O => \N__65718\,
            I => \N__65034\
        );

    \I__16301\ : ClkMux
    port map (
            O => \N__65717\,
            I => \N__65034\
        );

    \I__16300\ : ClkMux
    port map (
            O => \N__65716\,
            I => \N__65034\
        );

    \I__16299\ : ClkMux
    port map (
            O => \N__65715\,
            I => \N__65034\
        );

    \I__16298\ : ClkMux
    port map (
            O => \N__65714\,
            I => \N__65034\
        );

    \I__16297\ : ClkMux
    port map (
            O => \N__65713\,
            I => \N__65034\
        );

    \I__16296\ : Glb2LocalMux
    port map (
            O => \N__65710\,
            I => \N__65034\
        );

    \I__16295\ : Glb2LocalMux
    port map (
            O => \N__65707\,
            I => \N__65034\
        );

    \I__16294\ : ClkMux
    port map (
            O => \N__65706\,
            I => \N__65034\
        );

    \I__16293\ : ClkMux
    port map (
            O => \N__65705\,
            I => \N__65034\
        );

    \I__16292\ : ClkMux
    port map (
            O => \N__65704\,
            I => \N__65034\
        );

    \I__16291\ : ClkMux
    port map (
            O => \N__65703\,
            I => \N__65034\
        );

    \I__16290\ : ClkMux
    port map (
            O => \N__65702\,
            I => \N__65034\
        );

    \I__16289\ : ClkMux
    port map (
            O => \N__65701\,
            I => \N__65034\
        );

    \I__16288\ : ClkMux
    port map (
            O => \N__65700\,
            I => \N__65034\
        );

    \I__16287\ : ClkMux
    port map (
            O => \N__65699\,
            I => \N__65034\
        );

    \I__16286\ : ClkMux
    port map (
            O => \N__65698\,
            I => \N__65034\
        );

    \I__16285\ : ClkMux
    port map (
            O => \N__65697\,
            I => \N__65034\
        );

    \I__16284\ : ClkMux
    port map (
            O => \N__65696\,
            I => \N__65034\
        );

    \I__16283\ : ClkMux
    port map (
            O => \N__65695\,
            I => \N__65034\
        );

    \I__16282\ : ClkMux
    port map (
            O => \N__65694\,
            I => \N__65034\
        );

    \I__16281\ : ClkMux
    port map (
            O => \N__65693\,
            I => \N__65034\
        );

    \I__16280\ : ClkMux
    port map (
            O => \N__65692\,
            I => \N__65034\
        );

    \I__16279\ : ClkMux
    port map (
            O => \N__65691\,
            I => \N__65034\
        );

    \I__16278\ : ClkMux
    port map (
            O => \N__65690\,
            I => \N__65034\
        );

    \I__16277\ : ClkMux
    port map (
            O => \N__65689\,
            I => \N__65034\
        );

    \I__16276\ : ClkMux
    port map (
            O => \N__65688\,
            I => \N__65034\
        );

    \I__16275\ : ClkMux
    port map (
            O => \N__65687\,
            I => \N__65034\
        );

    \I__16274\ : ClkMux
    port map (
            O => \N__65686\,
            I => \N__65034\
        );

    \I__16273\ : ClkMux
    port map (
            O => \N__65685\,
            I => \N__65034\
        );

    \I__16272\ : ClkMux
    port map (
            O => \N__65684\,
            I => \N__65034\
        );

    \I__16271\ : ClkMux
    port map (
            O => \N__65683\,
            I => \N__65034\
        );

    \I__16270\ : ClkMux
    port map (
            O => \N__65682\,
            I => \N__65034\
        );

    \I__16269\ : ClkMux
    port map (
            O => \N__65681\,
            I => \N__65034\
        );

    \I__16268\ : ClkMux
    port map (
            O => \N__65680\,
            I => \N__65034\
        );

    \I__16267\ : ClkMux
    port map (
            O => \N__65679\,
            I => \N__65034\
        );

    \I__16266\ : ClkMux
    port map (
            O => \N__65678\,
            I => \N__65034\
        );

    \I__16265\ : ClkMux
    port map (
            O => \N__65677\,
            I => \N__65034\
        );

    \I__16264\ : ClkMux
    port map (
            O => \N__65676\,
            I => \N__65034\
        );

    \I__16263\ : ClkMux
    port map (
            O => \N__65675\,
            I => \N__65034\
        );

    \I__16262\ : ClkMux
    port map (
            O => \N__65674\,
            I => \N__65034\
        );

    \I__16261\ : ClkMux
    port map (
            O => \N__65673\,
            I => \N__65034\
        );

    \I__16260\ : ClkMux
    port map (
            O => \N__65672\,
            I => \N__65034\
        );

    \I__16259\ : ClkMux
    port map (
            O => \N__65671\,
            I => \N__65034\
        );

    \I__16258\ : ClkMux
    port map (
            O => \N__65670\,
            I => \N__65034\
        );

    \I__16257\ : ClkMux
    port map (
            O => \N__65669\,
            I => \N__65034\
        );

    \I__16256\ : ClkMux
    port map (
            O => \N__65668\,
            I => \N__65034\
        );

    \I__16255\ : ClkMux
    port map (
            O => \N__65667\,
            I => \N__65034\
        );

    \I__16254\ : ClkMux
    port map (
            O => \N__65666\,
            I => \N__65034\
        );

    \I__16253\ : ClkMux
    port map (
            O => \N__65665\,
            I => \N__65034\
        );

    \I__16252\ : ClkMux
    port map (
            O => \N__65664\,
            I => \N__65034\
        );

    \I__16251\ : ClkMux
    port map (
            O => \N__65663\,
            I => \N__65034\
        );

    \I__16250\ : ClkMux
    port map (
            O => \N__65662\,
            I => \N__65034\
        );

    \I__16249\ : ClkMux
    port map (
            O => \N__65661\,
            I => \N__65034\
        );

    \I__16248\ : ClkMux
    port map (
            O => \N__65660\,
            I => \N__65034\
        );

    \I__16247\ : ClkMux
    port map (
            O => \N__65659\,
            I => \N__65034\
        );

    \I__16246\ : ClkMux
    port map (
            O => \N__65658\,
            I => \N__65034\
        );

    \I__16245\ : ClkMux
    port map (
            O => \N__65657\,
            I => \N__65034\
        );

    \I__16244\ : ClkMux
    port map (
            O => \N__65656\,
            I => \N__65034\
        );

    \I__16243\ : ClkMux
    port map (
            O => \N__65655\,
            I => \N__65034\
        );

    \I__16242\ : ClkMux
    port map (
            O => \N__65654\,
            I => \N__65034\
        );

    \I__16241\ : ClkMux
    port map (
            O => \N__65653\,
            I => \N__65034\
        );

    \I__16240\ : ClkMux
    port map (
            O => \N__65652\,
            I => \N__65034\
        );

    \I__16239\ : ClkMux
    port map (
            O => \N__65651\,
            I => \N__65034\
        );

    \I__16238\ : ClkMux
    port map (
            O => \N__65650\,
            I => \N__65034\
        );

    \I__16237\ : ClkMux
    port map (
            O => \N__65649\,
            I => \N__65034\
        );

    \I__16236\ : ClkMux
    port map (
            O => \N__65648\,
            I => \N__65034\
        );

    \I__16235\ : ClkMux
    port map (
            O => \N__65647\,
            I => \N__65034\
        );

    \I__16234\ : ClkMux
    port map (
            O => \N__65646\,
            I => \N__65034\
        );

    \I__16233\ : ClkMux
    port map (
            O => \N__65645\,
            I => \N__65034\
        );

    \I__16232\ : ClkMux
    port map (
            O => \N__65644\,
            I => \N__65034\
        );

    \I__16231\ : ClkMux
    port map (
            O => \N__65643\,
            I => \N__65034\
        );

    \I__16230\ : ClkMux
    port map (
            O => \N__65642\,
            I => \N__65034\
        );

    \I__16229\ : ClkMux
    port map (
            O => \N__65641\,
            I => \N__65034\
        );

    \I__16228\ : ClkMux
    port map (
            O => \N__65640\,
            I => \N__65034\
        );

    \I__16227\ : ClkMux
    port map (
            O => \N__65639\,
            I => \N__65034\
        );

    \I__16226\ : ClkMux
    port map (
            O => \N__65638\,
            I => \N__65034\
        );

    \I__16225\ : ClkMux
    port map (
            O => \N__65637\,
            I => \N__65034\
        );

    \I__16224\ : ClkMux
    port map (
            O => \N__65636\,
            I => \N__65034\
        );

    \I__16223\ : ClkMux
    port map (
            O => \N__65635\,
            I => \N__65034\
        );

    \I__16222\ : ClkMux
    port map (
            O => \N__65634\,
            I => \N__65034\
        );

    \I__16221\ : ClkMux
    port map (
            O => \N__65633\,
            I => \N__65034\
        );

    \I__16220\ : ClkMux
    port map (
            O => \N__65632\,
            I => \N__65034\
        );

    \I__16219\ : ClkMux
    port map (
            O => \N__65631\,
            I => \N__65034\
        );

    \I__16218\ : ClkMux
    port map (
            O => \N__65630\,
            I => \N__65034\
        );

    \I__16217\ : ClkMux
    port map (
            O => \N__65629\,
            I => \N__65034\
        );

    \I__16216\ : ClkMux
    port map (
            O => \N__65628\,
            I => \N__65034\
        );

    \I__16215\ : ClkMux
    port map (
            O => \N__65627\,
            I => \N__65034\
        );

    \I__16214\ : ClkMux
    port map (
            O => \N__65626\,
            I => \N__65034\
        );

    \I__16213\ : ClkMux
    port map (
            O => \N__65625\,
            I => \N__65034\
        );

    \I__16212\ : ClkMux
    port map (
            O => \N__65624\,
            I => \N__65034\
        );

    \I__16211\ : ClkMux
    port map (
            O => \N__65623\,
            I => \N__65034\
        );

    \I__16210\ : ClkMux
    port map (
            O => \N__65622\,
            I => \N__65034\
        );

    \I__16209\ : ClkMux
    port map (
            O => \N__65621\,
            I => \N__65034\
        );

    \I__16208\ : ClkMux
    port map (
            O => \N__65620\,
            I => \N__65034\
        );

    \I__16207\ : ClkMux
    port map (
            O => \N__65619\,
            I => \N__65034\
        );

    \I__16206\ : ClkMux
    port map (
            O => \N__65618\,
            I => \N__65034\
        );

    \I__16205\ : ClkMux
    port map (
            O => \N__65617\,
            I => \N__65034\
        );

    \I__16204\ : ClkMux
    port map (
            O => \N__65616\,
            I => \N__65034\
        );

    \I__16203\ : ClkMux
    port map (
            O => \N__65615\,
            I => \N__65034\
        );

    \I__16202\ : ClkMux
    port map (
            O => \N__65614\,
            I => \N__65034\
        );

    \I__16201\ : ClkMux
    port map (
            O => \N__65613\,
            I => \N__65034\
        );

    \I__16200\ : ClkMux
    port map (
            O => \N__65612\,
            I => \N__65034\
        );

    \I__16199\ : ClkMux
    port map (
            O => \N__65611\,
            I => \N__65034\
        );

    \I__16198\ : ClkMux
    port map (
            O => \N__65610\,
            I => \N__65034\
        );

    \I__16197\ : ClkMux
    port map (
            O => \N__65609\,
            I => \N__65034\
        );

    \I__16196\ : ClkMux
    port map (
            O => \N__65608\,
            I => \N__65034\
        );

    \I__16195\ : ClkMux
    port map (
            O => \N__65607\,
            I => \N__65034\
        );

    \I__16194\ : ClkMux
    port map (
            O => \N__65606\,
            I => \N__65034\
        );

    \I__16193\ : ClkMux
    port map (
            O => \N__65605\,
            I => \N__65034\
        );

    \I__16192\ : ClkMux
    port map (
            O => \N__65604\,
            I => \N__65034\
        );

    \I__16191\ : ClkMux
    port map (
            O => \N__65603\,
            I => \N__65034\
        );

    \I__16190\ : ClkMux
    port map (
            O => \N__65602\,
            I => \N__65034\
        );

    \I__16189\ : ClkMux
    port map (
            O => \N__65601\,
            I => \N__65034\
        );

    \I__16188\ : ClkMux
    port map (
            O => \N__65600\,
            I => \N__65034\
        );

    \I__16187\ : ClkMux
    port map (
            O => \N__65599\,
            I => \N__65034\
        );

    \I__16186\ : ClkMux
    port map (
            O => \N__65598\,
            I => \N__65034\
        );

    \I__16185\ : ClkMux
    port map (
            O => \N__65597\,
            I => \N__65034\
        );

    \I__16184\ : ClkMux
    port map (
            O => \N__65596\,
            I => \N__65034\
        );

    \I__16183\ : ClkMux
    port map (
            O => \N__65595\,
            I => \N__65034\
        );

    \I__16182\ : ClkMux
    port map (
            O => \N__65594\,
            I => \N__65034\
        );

    \I__16181\ : ClkMux
    port map (
            O => \N__65593\,
            I => \N__65034\
        );

    \I__16180\ : ClkMux
    port map (
            O => \N__65592\,
            I => \N__65034\
        );

    \I__16179\ : ClkMux
    port map (
            O => \N__65591\,
            I => \N__65034\
        );

    \I__16178\ : ClkMux
    port map (
            O => \N__65590\,
            I => \N__65034\
        );

    \I__16177\ : ClkMux
    port map (
            O => \N__65589\,
            I => \N__65034\
        );

    \I__16176\ : ClkMux
    port map (
            O => \N__65588\,
            I => \N__65034\
        );

    \I__16175\ : ClkMux
    port map (
            O => \N__65587\,
            I => \N__65034\
        );

    \I__16174\ : ClkMux
    port map (
            O => \N__65586\,
            I => \N__65034\
        );

    \I__16173\ : ClkMux
    port map (
            O => \N__65585\,
            I => \N__65034\
        );

    \I__16172\ : ClkMux
    port map (
            O => \N__65584\,
            I => \N__65034\
        );

    \I__16171\ : ClkMux
    port map (
            O => \N__65583\,
            I => \N__65034\
        );

    \I__16170\ : ClkMux
    port map (
            O => \N__65582\,
            I => \N__65034\
        );

    \I__16169\ : ClkMux
    port map (
            O => \N__65581\,
            I => \N__65034\
        );

    \I__16168\ : ClkMux
    port map (
            O => \N__65580\,
            I => \N__65034\
        );

    \I__16167\ : ClkMux
    port map (
            O => \N__65579\,
            I => \N__65034\
        );

    \I__16166\ : ClkMux
    port map (
            O => \N__65578\,
            I => \N__65034\
        );

    \I__16165\ : ClkMux
    port map (
            O => \N__65577\,
            I => \N__65034\
        );

    \I__16164\ : ClkMux
    port map (
            O => \N__65576\,
            I => \N__65034\
        );

    \I__16163\ : ClkMux
    port map (
            O => \N__65575\,
            I => \N__65034\
        );

    \I__16162\ : ClkMux
    port map (
            O => \N__65574\,
            I => \N__65034\
        );

    \I__16161\ : ClkMux
    port map (
            O => \N__65573\,
            I => \N__65034\
        );

    \I__16160\ : ClkMux
    port map (
            O => \N__65572\,
            I => \N__65034\
        );

    \I__16159\ : ClkMux
    port map (
            O => \N__65571\,
            I => \N__65034\
        );

    \I__16158\ : ClkMux
    port map (
            O => \N__65570\,
            I => \N__65034\
        );

    \I__16157\ : ClkMux
    port map (
            O => \N__65569\,
            I => \N__65034\
        );

    \I__16156\ : ClkMux
    port map (
            O => \N__65568\,
            I => \N__65034\
        );

    \I__16155\ : ClkMux
    port map (
            O => \N__65567\,
            I => \N__65034\
        );

    \I__16154\ : ClkMux
    port map (
            O => \N__65566\,
            I => \N__65034\
        );

    \I__16153\ : ClkMux
    port map (
            O => \N__65565\,
            I => \N__65034\
        );

    \I__16152\ : ClkMux
    port map (
            O => \N__65564\,
            I => \N__65034\
        );

    \I__16151\ : ClkMux
    port map (
            O => \N__65563\,
            I => \N__65034\
        );

    \I__16150\ : ClkMux
    port map (
            O => \N__65562\,
            I => \N__65034\
        );

    \I__16149\ : ClkMux
    port map (
            O => \N__65561\,
            I => \N__65034\
        );

    \I__16148\ : ClkMux
    port map (
            O => \N__65560\,
            I => \N__65034\
        );

    \I__16147\ : ClkMux
    port map (
            O => \N__65559\,
            I => \N__65034\
        );

    \I__16146\ : ClkMux
    port map (
            O => \N__65558\,
            I => \N__65034\
        );

    \I__16145\ : ClkMux
    port map (
            O => \N__65557\,
            I => \N__65034\
        );

    \I__16144\ : ClkMux
    port map (
            O => \N__65556\,
            I => \N__65034\
        );

    \I__16143\ : ClkMux
    port map (
            O => \N__65555\,
            I => \N__65034\
        );

    \I__16142\ : ClkMux
    port map (
            O => \N__65554\,
            I => \N__65034\
        );

    \I__16141\ : ClkMux
    port map (
            O => \N__65553\,
            I => \N__65034\
        );

    \I__16140\ : ClkMux
    port map (
            O => \N__65552\,
            I => \N__65034\
        );

    \I__16139\ : ClkMux
    port map (
            O => \N__65551\,
            I => \N__65034\
        );

    \I__16138\ : ClkMux
    port map (
            O => \N__65550\,
            I => \N__65034\
        );

    \I__16137\ : ClkMux
    port map (
            O => \N__65549\,
            I => \N__65034\
        );

    \I__16136\ : ClkMux
    port map (
            O => \N__65548\,
            I => \N__65034\
        );

    \I__16135\ : ClkMux
    port map (
            O => \N__65547\,
            I => \N__65034\
        );

    \I__16134\ : ClkMux
    port map (
            O => \N__65546\,
            I => \N__65034\
        );

    \I__16133\ : ClkMux
    port map (
            O => \N__65545\,
            I => \N__65034\
        );

    \I__16132\ : ClkMux
    port map (
            O => \N__65544\,
            I => \N__65034\
        );

    \I__16131\ : ClkMux
    port map (
            O => \N__65543\,
            I => \N__65034\
        );

    \I__16130\ : ClkMux
    port map (
            O => \N__65542\,
            I => \N__65034\
        );

    \I__16129\ : ClkMux
    port map (
            O => \N__65541\,
            I => \N__65034\
        );

    \I__16128\ : ClkMux
    port map (
            O => \N__65540\,
            I => \N__65034\
        );

    \I__16127\ : ClkMux
    port map (
            O => \N__65539\,
            I => \N__65034\
        );

    \I__16126\ : ClkMux
    port map (
            O => \N__65538\,
            I => \N__65034\
        );

    \I__16125\ : ClkMux
    port map (
            O => \N__65537\,
            I => \N__65034\
        );

    \I__16124\ : ClkMux
    port map (
            O => \N__65536\,
            I => \N__65034\
        );

    \I__16123\ : ClkMux
    port map (
            O => \N__65535\,
            I => \N__65034\
        );

    \I__16122\ : ClkMux
    port map (
            O => \N__65534\,
            I => \N__65034\
        );

    \I__16121\ : ClkMux
    port map (
            O => \N__65533\,
            I => \N__65034\
        );

    \I__16120\ : ClkMux
    port map (
            O => \N__65532\,
            I => \N__65034\
        );

    \I__16119\ : ClkMux
    port map (
            O => \N__65531\,
            I => \N__65034\
        );

    \I__16118\ : ClkMux
    port map (
            O => \N__65530\,
            I => \N__65034\
        );

    \I__16117\ : ClkMux
    port map (
            O => \N__65529\,
            I => \N__65034\
        );

    \I__16116\ : ClkMux
    port map (
            O => \N__65528\,
            I => \N__65034\
        );

    \I__16115\ : ClkMux
    port map (
            O => \N__65527\,
            I => \N__65034\
        );

    \I__16114\ : ClkMux
    port map (
            O => \N__65526\,
            I => \N__65034\
        );

    \I__16113\ : ClkMux
    port map (
            O => \N__65525\,
            I => \N__65034\
        );

    \I__16112\ : ClkMux
    port map (
            O => \N__65524\,
            I => \N__65034\
        );

    \I__16111\ : ClkMux
    port map (
            O => \N__65523\,
            I => \N__65034\
        );

    \I__16110\ : ClkMux
    port map (
            O => \N__65522\,
            I => \N__65034\
        );

    \I__16109\ : ClkMux
    port map (
            O => \N__65521\,
            I => \N__65034\
        );

    \I__16108\ : ClkMux
    port map (
            O => \N__65520\,
            I => \N__65034\
        );

    \I__16107\ : ClkMux
    port map (
            O => \N__65519\,
            I => \N__65034\
        );

    \I__16106\ : ClkMux
    port map (
            O => \N__65518\,
            I => \N__65034\
        );

    \I__16105\ : ClkMux
    port map (
            O => \N__65517\,
            I => \N__65034\
        );

    \I__16104\ : ClkMux
    port map (
            O => \N__65516\,
            I => \N__65034\
        );

    \I__16103\ : ClkMux
    port map (
            O => \N__65515\,
            I => \N__65034\
        );

    \I__16102\ : ClkMux
    port map (
            O => \N__65514\,
            I => \N__65034\
        );

    \I__16101\ : ClkMux
    port map (
            O => \N__65513\,
            I => \N__65034\
        );

    \I__16100\ : GlobalMux
    port map (
            O => \N__65034\,
            I => \N__65031\
        );

    \I__16099\ : gio2CtrlBuf
    port map (
            O => \N__65031\,
            I => clock_c_g
        );

    \I__16098\ : SRMux
    port map (
            O => \N__65028\,
            I => \N__64830\
        );

    \I__16097\ : SRMux
    port map (
            O => \N__65027\,
            I => \N__64830\
        );

    \I__16096\ : SRMux
    port map (
            O => \N__65026\,
            I => \N__64830\
        );

    \I__16095\ : SRMux
    port map (
            O => \N__65025\,
            I => \N__64830\
        );

    \I__16094\ : SRMux
    port map (
            O => \N__65024\,
            I => \N__64830\
        );

    \I__16093\ : SRMux
    port map (
            O => \N__65023\,
            I => \N__64830\
        );

    \I__16092\ : SRMux
    port map (
            O => \N__65022\,
            I => \N__64830\
        );

    \I__16091\ : SRMux
    port map (
            O => \N__65021\,
            I => \N__64830\
        );

    \I__16090\ : SRMux
    port map (
            O => \N__65020\,
            I => \N__64830\
        );

    \I__16089\ : SRMux
    port map (
            O => \N__65019\,
            I => \N__64830\
        );

    \I__16088\ : SRMux
    port map (
            O => \N__65018\,
            I => \N__64830\
        );

    \I__16087\ : SRMux
    port map (
            O => \N__65017\,
            I => \N__64830\
        );

    \I__16086\ : SRMux
    port map (
            O => \N__65016\,
            I => \N__64830\
        );

    \I__16085\ : SRMux
    port map (
            O => \N__65015\,
            I => \N__64830\
        );

    \I__16084\ : SRMux
    port map (
            O => \N__65014\,
            I => \N__64830\
        );

    \I__16083\ : SRMux
    port map (
            O => \N__65013\,
            I => \N__64830\
        );

    \I__16082\ : SRMux
    port map (
            O => \N__65012\,
            I => \N__64830\
        );

    \I__16081\ : SRMux
    port map (
            O => \N__65011\,
            I => \N__64830\
        );

    \I__16080\ : SRMux
    port map (
            O => \N__65010\,
            I => \N__64830\
        );

    \I__16079\ : SRMux
    port map (
            O => \N__65009\,
            I => \N__64830\
        );

    \I__16078\ : SRMux
    port map (
            O => \N__65008\,
            I => \N__64830\
        );

    \I__16077\ : SRMux
    port map (
            O => \N__65007\,
            I => \N__64830\
        );

    \I__16076\ : SRMux
    port map (
            O => \N__65006\,
            I => \N__64830\
        );

    \I__16075\ : SRMux
    port map (
            O => \N__65005\,
            I => \N__64830\
        );

    \I__16074\ : SRMux
    port map (
            O => \N__65004\,
            I => \N__64830\
        );

    \I__16073\ : SRMux
    port map (
            O => \N__65003\,
            I => \N__64830\
        );

    \I__16072\ : SRMux
    port map (
            O => \N__65002\,
            I => \N__64830\
        );

    \I__16071\ : SRMux
    port map (
            O => \N__65001\,
            I => \N__64830\
        );

    \I__16070\ : SRMux
    port map (
            O => \N__65000\,
            I => \N__64830\
        );

    \I__16069\ : SRMux
    port map (
            O => \N__64999\,
            I => \N__64830\
        );

    \I__16068\ : SRMux
    port map (
            O => \N__64998\,
            I => \N__64830\
        );

    \I__16067\ : SRMux
    port map (
            O => \N__64997\,
            I => \N__64830\
        );

    \I__16066\ : SRMux
    port map (
            O => \N__64996\,
            I => \N__64830\
        );

    \I__16065\ : SRMux
    port map (
            O => \N__64995\,
            I => \N__64830\
        );

    \I__16064\ : SRMux
    port map (
            O => \N__64994\,
            I => \N__64830\
        );

    \I__16063\ : SRMux
    port map (
            O => \N__64993\,
            I => \N__64830\
        );

    \I__16062\ : SRMux
    port map (
            O => \N__64992\,
            I => \N__64830\
        );

    \I__16061\ : SRMux
    port map (
            O => \N__64991\,
            I => \N__64830\
        );

    \I__16060\ : SRMux
    port map (
            O => \N__64990\,
            I => \N__64830\
        );

    \I__16059\ : SRMux
    port map (
            O => \N__64989\,
            I => \N__64830\
        );

    \I__16058\ : SRMux
    port map (
            O => \N__64988\,
            I => \N__64830\
        );

    \I__16057\ : SRMux
    port map (
            O => \N__64987\,
            I => \N__64830\
        );

    \I__16056\ : SRMux
    port map (
            O => \N__64986\,
            I => \N__64830\
        );

    \I__16055\ : SRMux
    port map (
            O => \N__64985\,
            I => \N__64830\
        );

    \I__16054\ : SRMux
    port map (
            O => \N__64984\,
            I => \N__64830\
        );

    \I__16053\ : SRMux
    port map (
            O => \N__64983\,
            I => \N__64830\
        );

    \I__16052\ : SRMux
    port map (
            O => \N__64982\,
            I => \N__64830\
        );

    \I__16051\ : SRMux
    port map (
            O => \N__64981\,
            I => \N__64830\
        );

    \I__16050\ : SRMux
    port map (
            O => \N__64980\,
            I => \N__64830\
        );

    \I__16049\ : SRMux
    port map (
            O => \N__64979\,
            I => \N__64830\
        );

    \I__16048\ : SRMux
    port map (
            O => \N__64978\,
            I => \N__64830\
        );

    \I__16047\ : SRMux
    port map (
            O => \N__64977\,
            I => \N__64830\
        );

    \I__16046\ : SRMux
    port map (
            O => \N__64976\,
            I => \N__64830\
        );

    \I__16045\ : SRMux
    port map (
            O => \N__64975\,
            I => \N__64830\
        );

    \I__16044\ : SRMux
    port map (
            O => \N__64974\,
            I => \N__64830\
        );

    \I__16043\ : SRMux
    port map (
            O => \N__64973\,
            I => \N__64830\
        );

    \I__16042\ : SRMux
    port map (
            O => \N__64972\,
            I => \N__64830\
        );

    \I__16041\ : SRMux
    port map (
            O => \N__64971\,
            I => \N__64830\
        );

    \I__16040\ : SRMux
    port map (
            O => \N__64970\,
            I => \N__64830\
        );

    \I__16039\ : SRMux
    port map (
            O => \N__64969\,
            I => \N__64830\
        );

    \I__16038\ : SRMux
    port map (
            O => \N__64968\,
            I => \N__64830\
        );

    \I__16037\ : SRMux
    port map (
            O => \N__64967\,
            I => \N__64830\
        );

    \I__16036\ : SRMux
    port map (
            O => \N__64966\,
            I => \N__64830\
        );

    \I__16035\ : SRMux
    port map (
            O => \N__64965\,
            I => \N__64830\
        );

    \I__16034\ : SRMux
    port map (
            O => \N__64964\,
            I => \N__64830\
        );

    \I__16033\ : SRMux
    port map (
            O => \N__64963\,
            I => \N__64830\
        );

    \I__16032\ : GlobalMux
    port map (
            O => \N__64830\,
            I => \N__64827\
        );

    \I__16031\ : gio2CtrlBuf
    port map (
            O => \N__64827\,
            I => \I2C_top_level_inst1.c_state4_0_i_g\
        );

    \I__16030\ : CascadeMux
    port map (
            O => \N__64824\,
            I => \N__64821\
        );

    \I__16029\ : InMux
    port map (
            O => \N__64821\,
            I => \N__64818\
        );

    \I__16028\ : LocalMux
    port map (
            O => \N__64818\,
            I => \N__64815\
        );

    \I__16027\ : Span4Mux_h
    port map (
            O => \N__64815\,
            I => \N__64812\
        );

    \I__16026\ : Odrv4
    port map (
            O => \N__64812\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666\
        );

    \I__16025\ : InMux
    port map (
            O => \N__64809\,
            I => \N__64806\
        );

    \I__16024\ : LocalMux
    port map (
            O => \N__64806\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_1\
        );

    \I__16023\ : InMux
    port map (
            O => \N__64803\,
            I => \N__64798\
        );

    \I__16022\ : InMux
    port map (
            O => \N__64802\,
            I => \N__64795\
        );

    \I__16021\ : CascadeMux
    port map (
            O => \N__64801\,
            I => \N__64791\
        );

    \I__16020\ : LocalMux
    port map (
            O => \N__64798\,
            I => \N__64784\
        );

    \I__16019\ : LocalMux
    port map (
            O => \N__64795\,
            I => \N__64781\
        );

    \I__16018\ : InMux
    port map (
            O => \N__64794\,
            I => \N__64778\
        );

    \I__16017\ : InMux
    port map (
            O => \N__64791\,
            I => \N__64775\
        );

    \I__16016\ : InMux
    port map (
            O => \N__64790\,
            I => \N__64772\
        );

    \I__16015\ : CascadeMux
    port map (
            O => \N__64789\,
            I => \N__64769\
        );

    \I__16014\ : InMux
    port map (
            O => \N__64788\,
            I => \N__64766\
        );

    \I__16013\ : InMux
    port map (
            O => \N__64787\,
            I => \N__64763\
        );

    \I__16012\ : Span4Mux_v
    port map (
            O => \N__64784\,
            I => \N__64756\
        );

    \I__16011\ : Span4Mux_v
    port map (
            O => \N__64781\,
            I => \N__64756\
        );

    \I__16010\ : LocalMux
    port map (
            O => \N__64778\,
            I => \N__64756\
        );

    \I__16009\ : LocalMux
    port map (
            O => \N__64775\,
            I => \N__64751\
        );

    \I__16008\ : LocalMux
    port map (
            O => \N__64772\,
            I => \N__64751\
        );

    \I__16007\ : InMux
    port map (
            O => \N__64769\,
            I => \N__64748\
        );

    \I__16006\ : LocalMux
    port map (
            O => \N__64766\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\
        );

    \I__16005\ : LocalMux
    port map (
            O => \N__64763\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\
        );

    \I__16004\ : Odrv4
    port map (
            O => \N__64756\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\
        );

    \I__16003\ : Odrv4
    port map (
            O => \N__64751\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\
        );

    \I__16002\ : LocalMux
    port map (
            O => \N__64748\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\
        );

    \I__16001\ : CascadeMux
    port map (
            O => \N__64737\,
            I => \N__64734\
        );

    \I__16000\ : InMux
    port map (
            O => \N__64734\,
            I => \N__64731\
        );

    \I__15999\ : LocalMux
    port map (
            O => \N__64731\,
            I => \N__64728\
        );

    \I__15998\ : Span4Mux_h
    port map (
            O => \N__64728\,
            I => \N__64725\
        );

    \I__15997\ : Odrv4
    port map (
            O => \N__64725\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_2_1\
        );

    \I__15996\ : InMux
    port map (
            O => \N__64722\,
            I => \N__64716\
        );

    \I__15995\ : InMux
    port map (
            O => \N__64721\,
            I => \N__64716\
        );

    \I__15994\ : LocalMux
    port map (
            O => \N__64716\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0\
        );

    \I__15993\ : InMux
    port map (
            O => \N__64713\,
            I => \N__64709\
        );

    \I__15992\ : InMux
    port map (
            O => \N__64712\,
            I => \N__64701\
        );

    \I__15991\ : LocalMux
    port map (
            O => \N__64709\,
            I => \N__64698\
        );

    \I__15990\ : InMux
    port map (
            O => \N__64708\,
            I => \N__64693\
        );

    \I__15989\ : InMux
    port map (
            O => \N__64707\,
            I => \N__64688\
        );

    \I__15988\ : InMux
    port map (
            O => \N__64706\,
            I => \N__64688\
        );

    \I__15987\ : InMux
    port map (
            O => \N__64705\,
            I => \N__64680\
        );

    \I__15986\ : InMux
    port map (
            O => \N__64704\,
            I => \N__64680\
        );

    \I__15985\ : LocalMux
    port map (
            O => \N__64701\,
            I => \N__64674\
        );

    \I__15984\ : Span4Mux_h
    port map (
            O => \N__64698\,
            I => \N__64674\
        );

    \I__15983\ : InMux
    port map (
            O => \N__64697\,
            I => \N__64669\
        );

    \I__15982\ : InMux
    port map (
            O => \N__64696\,
            I => \N__64669\
        );

    \I__15981\ : LocalMux
    port map (
            O => \N__64693\,
            I => \N__64664\
        );

    \I__15980\ : LocalMux
    port map (
            O => \N__64688\,
            I => \N__64664\
        );

    \I__15979\ : InMux
    port map (
            O => \N__64687\,
            I => \N__64657\
        );

    \I__15978\ : InMux
    port map (
            O => \N__64686\,
            I => \N__64657\
        );

    \I__15977\ : InMux
    port map (
            O => \N__64685\,
            I => \N__64657\
        );

    \I__15976\ : LocalMux
    port map (
            O => \N__64680\,
            I => \N__64654\
        );

    \I__15975\ : InMux
    port map (
            O => \N__64679\,
            I => \N__64651\
        );

    \I__15974\ : Span4Mux_h
    port map (
            O => \N__64674\,
            I => \N__64648\
        );

    \I__15973\ : LocalMux
    port map (
            O => \N__64669\,
            I => \N__64641\
        );

    \I__15972\ : Span4Mux_v
    port map (
            O => \N__64664\,
            I => \N__64641\
        );

    \I__15971\ : LocalMux
    port map (
            O => \N__64657\,
            I => \N__64641\
        );

    \I__15970\ : Span4Mux_h
    port map (
            O => \N__64654\,
            I => \N__64638\
        );

    \I__15969\ : LocalMux
    port map (
            O => \N__64651\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7\
        );

    \I__15968\ : Odrv4
    port map (
            O => \N__64648\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7\
        );

    \I__15967\ : Odrv4
    port map (
            O => \N__64641\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7\
        );

    \I__15966\ : Odrv4
    port map (
            O => \N__64638\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7\
        );

    \I__15965\ : InMux
    port map (
            O => \N__64629\,
            I => \N__64626\
        );

    \I__15964\ : LocalMux
    port map (
            O => \N__64626\,
            I => \N__64623\
        );

    \I__15963\ : Span4Mux_h
    port map (
            O => \N__64623\,
            I => \N__64620\
        );

    \I__15962\ : Odrv4
    port map (
            O => \N__64620\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o3_1\
        );

    \I__15961\ : CascadeMux
    port map (
            O => \N__64617\,
            I => \N__64614\
        );

    \I__15960\ : InMux
    port map (
            O => \N__64614\,
            I => \N__64611\
        );

    \I__15959\ : LocalMux
    port map (
            O => \N__64611\,
            I => \N__64608\
        );

    \I__15958\ : Odrv4
    port map (
            O => \N__64608\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1802\
        );

    \I__15957\ : InMux
    port map (
            O => \N__64605\,
            I => \N__64602\
        );

    \I__15956\ : LocalMux
    port map (
            O => \N__64602\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1609_0\
        );

    \I__15955\ : InMux
    port map (
            O => \N__64599\,
            I => \N__64596\
        );

    \I__15954\ : LocalMux
    port map (
            O => \N__64596\,
            I => \N__64593\
        );

    \I__15953\ : Span4Mux_v
    port map (
            O => \N__64593\,
            I => \N__64590\
        );

    \I__15952\ : Span4Mux_h
    port map (
            O => \N__64590\,
            I => \N__64587\
        );

    \I__15951\ : Odrv4
    port map (
            O => \N__64587\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa\
        );

    \I__15950\ : CascadeMux
    port map (
            O => \N__64584\,
            I => \N__64578\
        );

    \I__15949\ : InMux
    port map (
            O => \N__64583\,
            I => \N__64561\
        );

    \I__15948\ : InMux
    port map (
            O => \N__64582\,
            I => \N__64561\
        );

    \I__15947\ : InMux
    port map (
            O => \N__64581\,
            I => \N__64561\
        );

    \I__15946\ : InMux
    port map (
            O => \N__64578\,
            I => \N__64561\
        );

    \I__15945\ : InMux
    port map (
            O => \N__64577\,
            I => \N__64552\
        );

    \I__15944\ : InMux
    port map (
            O => \N__64576\,
            I => \N__64552\
        );

    \I__15943\ : InMux
    port map (
            O => \N__64575\,
            I => \N__64552\
        );

    \I__15942\ : InMux
    port map (
            O => \N__64574\,
            I => \N__64552\
        );

    \I__15941\ : InMux
    port map (
            O => \N__64573\,
            I => \N__64542\
        );

    \I__15940\ : InMux
    port map (
            O => \N__64572\,
            I => \N__64542\
        );

    \I__15939\ : InMux
    port map (
            O => \N__64571\,
            I => \N__64542\
        );

    \I__15938\ : InMux
    port map (
            O => \N__64570\,
            I => \N__64542\
        );

    \I__15937\ : LocalMux
    port map (
            O => \N__64561\,
            I => \N__64539\
        );

    \I__15936\ : LocalMux
    port map (
            O => \N__64552\,
            I => \N__64536\
        );

    \I__15935\ : InMux
    port map (
            O => \N__64551\,
            I => \N__64533\
        );

    \I__15934\ : LocalMux
    port map (
            O => \N__64542\,
            I => \N__64526\
        );

    \I__15933\ : Span4Mux_v
    port map (
            O => \N__64539\,
            I => \N__64526\
        );

    \I__15932\ : Span4Mux_v
    port map (
            O => \N__64536\,
            I => \N__64526\
        );

    \I__15931\ : LocalMux
    port map (
            O => \N__64533\,
            I => \N__64523\
        );

    \I__15930\ : Span4Mux_h
    port map (
            O => \N__64526\,
            I => \N__64518\
        );

    \I__15929\ : Span4Mux_v
    port map (
            O => \N__64523\,
            I => \N__64518\
        );

    \I__15928\ : Odrv4
    port map (
            O => \N__64518\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0\
        );

    \I__15927\ : CascadeMux
    port map (
            O => \N__64515\,
            I => \N__64512\
        );

    \I__15926\ : InMux
    port map (
            O => \N__64512\,
            I => \N__64509\
        );

    \I__15925\ : LocalMux
    port map (
            O => \N__64509\,
            I => \N__64506\
        );

    \I__15924\ : Span4Mux_h
    port map (
            O => \N__64506\,
            I => \N__64503\
        );

    \I__15923\ : Span4Mux_h
    port map (
            O => \N__64503\,
            I => \N__64500\
        );

    \I__15922\ : Odrv4
    port map (
            O => \N__64500\,
            I => \I2C_top_level_inst1.s_addr0_o_0\
        );

    \I__15921\ : InMux
    port map (
            O => \N__64497\,
            I => \N__64493\
        );

    \I__15920\ : InMux
    port map (
            O => \N__64496\,
            I => \N__64490\
        );

    \I__15919\ : LocalMux
    port map (
            O => \N__64493\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_691\
        );

    \I__15918\ : LocalMux
    port map (
            O => \N__64490\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_691\
        );

    \I__15917\ : InMux
    port map (
            O => \N__64485\,
            I => \N__64482\
        );

    \I__15916\ : LocalMux
    port map (
            O => \N__64482\,
            I => \N__64479\
        );

    \I__15915\ : Odrv12
    port map (
            O => \N__64479\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_0\
        );

    \I__15914\ : CascadeMux
    port map (
            O => \N__64476\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_295_cascade_\
        );

    \I__15913\ : InMux
    port map (
            O => \N__64473\,
            I => \N__64469\
        );

    \I__15912\ : InMux
    port map (
            O => \N__64472\,
            I => \N__64466\
        );

    \I__15911\ : LocalMux
    port map (
            O => \N__64469\,
            I => \N__64462\
        );

    \I__15910\ : LocalMux
    port map (
            O => \N__64466\,
            I => \N__64459\
        );

    \I__15909\ : InMux
    port map (
            O => \N__64465\,
            I => \N__64454\
        );

    \I__15908\ : Span4Mux_v
    port map (
            O => \N__64462\,
            I => \N__64449\
        );

    \I__15907\ : Span4Mux_h
    port map (
            O => \N__64459\,
            I => \N__64449\
        );

    \I__15906\ : InMux
    port map (
            O => \N__64458\,
            I => \N__64444\
        );

    \I__15905\ : InMux
    port map (
            O => \N__64457\,
            I => \N__64444\
        );

    \I__15904\ : LocalMux
    port map (
            O => \N__64454\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3\
        );

    \I__15903\ : Odrv4
    port map (
            O => \N__64449\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3\
        );

    \I__15902\ : LocalMux
    port map (
            O => \N__64444\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3\
        );

    \I__15901\ : CascadeMux
    port map (
            O => \N__64437\,
            I => \N__64434\
        );

    \I__15900\ : InMux
    port map (
            O => \N__64434\,
            I => \N__64429\
        );

    \I__15899\ : InMux
    port map (
            O => \N__64433\,
            I => \N__64426\
        );

    \I__15898\ : InMux
    port map (
            O => \N__64432\,
            I => \N__64422\
        );

    \I__15897\ : LocalMux
    port map (
            O => \N__64429\,
            I => \N__64417\
        );

    \I__15896\ : LocalMux
    port map (
            O => \N__64426\,
            I => \N__64414\
        );

    \I__15895\ : InMux
    port map (
            O => \N__64425\,
            I => \N__64411\
        );

    \I__15894\ : LocalMux
    port map (
            O => \N__64422\,
            I => \N__64408\
        );

    \I__15893\ : InMux
    port map (
            O => \N__64421\,
            I => \N__64401\
        );

    \I__15892\ : InMux
    port map (
            O => \N__64420\,
            I => \N__64401\
        );

    \I__15891\ : Span4Mux_h
    port map (
            O => \N__64417\,
            I => \N__64398\
        );

    \I__15890\ : Span4Mux_h
    port map (
            O => \N__64414\,
            I => \N__64393\
        );

    \I__15889\ : LocalMux
    port map (
            O => \N__64411\,
            I => \N__64393\
        );

    \I__15888\ : Span4Mux_h
    port map (
            O => \N__64408\,
            I => \N__64390\
        );

    \I__15887\ : InMux
    port map (
            O => \N__64407\,
            I => \N__64385\
        );

    \I__15886\ : InMux
    port map (
            O => \N__64406\,
            I => \N__64385\
        );

    \I__15885\ : LocalMux
    port map (
            O => \N__64401\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\
        );

    \I__15884\ : Odrv4
    port map (
            O => \N__64398\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\
        );

    \I__15883\ : Odrv4
    port map (
            O => \N__64393\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\
        );

    \I__15882\ : Odrv4
    port map (
            O => \N__64390\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\
        );

    \I__15881\ : LocalMux
    port map (
            O => \N__64385\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\
        );

    \I__15880\ : InMux
    port map (
            O => \N__64374\,
            I => \N__64371\
        );

    \I__15879\ : LocalMux
    port map (
            O => \N__64371\,
            I => \N__64368\
        );

    \I__15878\ : Span4Mux_h
    port map (
            O => \N__64368\,
            I => \N__64365\
        );

    \I__15877\ : Span4Mux_h
    port map (
            O => \N__64365\,
            I => \N__64362\
        );

    \I__15876\ : Odrv4
    port map (
            O => \N__64362\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_6\
        );

    \I__15875\ : InMux
    port map (
            O => \N__64359\,
            I => \N__64356\
        );

    \I__15874\ : LocalMux
    port map (
            O => \N__64356\,
            I => \N__64352\
        );

    \I__15873\ : InMux
    port map (
            O => \N__64355\,
            I => \N__64349\
        );

    \I__15872\ : Odrv4
    port map (
            O => \N__64352\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0\
        );

    \I__15871\ : LocalMux
    port map (
            O => \N__64349\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0\
        );

    \I__15870\ : InMux
    port map (
            O => \N__64344\,
            I => \N__64340\
        );

    \I__15869\ : InMux
    port map (
            O => \N__64343\,
            I => \N__64337\
        );

    \I__15868\ : LocalMux
    port map (
            O => \N__64340\,
            I => \N__64334\
        );

    \I__15867\ : LocalMux
    port map (
            O => \N__64337\,
            I => \N__64331\
        );

    \I__15866\ : Span4Mux_h
    port map (
            O => \N__64334\,
            I => \N__64328\
        );

    \I__15865\ : Odrv4
    port map (
            O => \N__64331\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2\
        );

    \I__15864\ : Odrv4
    port map (
            O => \N__64328\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2\
        );

    \I__15863\ : InMux
    port map (
            O => \N__64323\,
            I => \N__64320\
        );

    \I__15862\ : LocalMux
    port map (
            O => \N__64320\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_277\
        );

    \I__15861\ : CascadeMux
    port map (
            O => \N__64317\,
            I => \N__64313\
        );

    \I__15860\ : InMux
    port map (
            O => \N__64316\,
            I => \N__64309\
        );

    \I__15859\ : InMux
    port map (
            O => \N__64313\,
            I => \N__64306\
        );

    \I__15858\ : InMux
    port map (
            O => \N__64312\,
            I => \N__64303\
        );

    \I__15857\ : LocalMux
    port map (
            O => \N__64309\,
            I => \N__64300\
        );

    \I__15856\ : LocalMux
    port map (
            O => \N__64306\,
            I => \N__64296\
        );

    \I__15855\ : LocalMux
    port map (
            O => \N__64303\,
            I => \N__64293\
        );

    \I__15854\ : Span4Mux_v
    port map (
            O => \N__64300\,
            I => \N__64290\
        );

    \I__15853\ : InMux
    port map (
            O => \N__64299\,
            I => \N__64287\
        );

    \I__15852\ : Span12Mux_h
    port map (
            O => \N__64296\,
            I => \N__64284\
        );

    \I__15851\ : Span4Mux_v
    port map (
            O => \N__64293\,
            I => \N__64281\
        );

    \I__15850\ : Sp12to4
    port map (
            O => \N__64290\,
            I => \N__64274\
        );

    \I__15849\ : LocalMux
    port map (
            O => \N__64287\,
            I => \N__64274\
        );

    \I__15848\ : Span12Mux_v
    port map (
            O => \N__64284\,
            I => \N__64274\
        );

    \I__15847\ : Odrv4
    port map (
            O => \N__64281\,
            I => \N_552_i\
        );

    \I__15846\ : Odrv12
    port map (
            O => \N__64274\,
            I => \N_552_i\
        );

    \I__15845\ : InMux
    port map (
            O => \N__64269\,
            I => \N__64262\
        );

    \I__15844\ : InMux
    port map (
            O => \N__64268\,
            I => \N__64256\
        );

    \I__15843\ : InMux
    port map (
            O => \N__64267\,
            I => \N__64253\
        );

    \I__15842\ : InMux
    port map (
            O => \N__64266\,
            I => \N__64240\
        );

    \I__15841\ : InMux
    port map (
            O => \N__64265\,
            I => \N__64237\
        );

    \I__15840\ : LocalMux
    port map (
            O => \N__64262\,
            I => \N__64231\
        );

    \I__15839\ : InMux
    port map (
            O => \N__64261\,
            I => \N__64225\
        );

    \I__15838\ : InMux
    port map (
            O => \N__64260\,
            I => \N__64220\
        );

    \I__15837\ : InMux
    port map (
            O => \N__64259\,
            I => \N__64220\
        );

    \I__15836\ : LocalMux
    port map (
            O => \N__64256\,
            I => \N__64210\
        );

    \I__15835\ : LocalMux
    port map (
            O => \N__64253\,
            I => \N__64198\
        );

    \I__15834\ : InMux
    port map (
            O => \N__64252\,
            I => \N__64193\
        );

    \I__15833\ : InMux
    port map (
            O => \N__64251\,
            I => \N__64193\
        );

    \I__15832\ : InMux
    port map (
            O => \N__64250\,
            I => \N__64190\
        );

    \I__15831\ : InMux
    port map (
            O => \N__64249\,
            I => \N__64175\
        );

    \I__15830\ : InMux
    port map (
            O => \N__64248\,
            I => \N__64175\
        );

    \I__15829\ : InMux
    port map (
            O => \N__64247\,
            I => \N__64175\
        );

    \I__15828\ : InMux
    port map (
            O => \N__64246\,
            I => \N__64175\
        );

    \I__15827\ : InMux
    port map (
            O => \N__64245\,
            I => \N__64175\
        );

    \I__15826\ : InMux
    port map (
            O => \N__64244\,
            I => \N__64175\
        );

    \I__15825\ : InMux
    port map (
            O => \N__64243\,
            I => \N__64175\
        );

    \I__15824\ : LocalMux
    port map (
            O => \N__64240\,
            I => \N__64169\
        );

    \I__15823\ : LocalMux
    port map (
            O => \N__64237\,
            I => \N__64166\
        );

    \I__15822\ : InMux
    port map (
            O => \N__64236\,
            I => \N__64161\
        );

    \I__15821\ : InMux
    port map (
            O => \N__64235\,
            I => \N__64161\
        );

    \I__15820\ : InMux
    port map (
            O => \N__64234\,
            I => \N__64158\
        );

    \I__15819\ : Span4Mux_h
    port map (
            O => \N__64231\,
            I => \N__64154\
        );

    \I__15818\ : InMux
    port map (
            O => \N__64230\,
            I => \N__64149\
        );

    \I__15817\ : InMux
    port map (
            O => \N__64229\,
            I => \N__64144\
        );

    \I__15816\ : InMux
    port map (
            O => \N__64228\,
            I => \N__64144\
        );

    \I__15815\ : LocalMux
    port map (
            O => \N__64225\,
            I => \N__64139\
        );

    \I__15814\ : LocalMux
    port map (
            O => \N__64220\,
            I => \N__64139\
        );

    \I__15813\ : InMux
    port map (
            O => \N__64219\,
            I => \N__64124\
        );

    \I__15812\ : InMux
    port map (
            O => \N__64218\,
            I => \N__64124\
        );

    \I__15811\ : InMux
    port map (
            O => \N__64217\,
            I => \N__64124\
        );

    \I__15810\ : InMux
    port map (
            O => \N__64216\,
            I => \N__64124\
        );

    \I__15809\ : InMux
    port map (
            O => \N__64215\,
            I => \N__64124\
        );

    \I__15808\ : InMux
    port map (
            O => \N__64214\,
            I => \N__64124\
        );

    \I__15807\ : InMux
    port map (
            O => \N__64213\,
            I => \N__64124\
        );

    \I__15806\ : Span4Mux_h
    port map (
            O => \N__64210\,
            I => \N__64121\
        );

    \I__15805\ : CascadeMux
    port map (
            O => \N__64209\,
            I => \N__64118\
        );

    \I__15804\ : InMux
    port map (
            O => \N__64208\,
            I => \N__64100\
        );

    \I__15803\ : InMux
    port map (
            O => \N__64207\,
            I => \N__64100\
        );

    \I__15802\ : InMux
    port map (
            O => \N__64206\,
            I => \N__64100\
        );

    \I__15801\ : InMux
    port map (
            O => \N__64205\,
            I => \N__64100\
        );

    \I__15800\ : InMux
    port map (
            O => \N__64204\,
            I => \N__64100\
        );

    \I__15799\ : InMux
    port map (
            O => \N__64203\,
            I => \N__64100\
        );

    \I__15798\ : InMux
    port map (
            O => \N__64202\,
            I => \N__64100\
        );

    \I__15797\ : InMux
    port map (
            O => \N__64201\,
            I => \N__64100\
        );

    \I__15796\ : Span4Mux_h
    port map (
            O => \N__64198\,
            I => \N__64095\
        );

    \I__15795\ : LocalMux
    port map (
            O => \N__64193\,
            I => \N__64095\
        );

    \I__15794\ : LocalMux
    port map (
            O => \N__64190\,
            I => \N__64092\
        );

    \I__15793\ : LocalMux
    port map (
            O => \N__64175\,
            I => \N__64089\
        );

    \I__15792\ : InMux
    port map (
            O => \N__64174\,
            I => \N__64082\
        );

    \I__15791\ : InMux
    port map (
            O => \N__64173\,
            I => \N__64082\
        );

    \I__15790\ : InMux
    port map (
            O => \N__64172\,
            I => \N__64082\
        );

    \I__15789\ : Span4Mux_h
    port map (
            O => \N__64169\,
            I => \N__64078\
        );

    \I__15788\ : Span4Mux_h
    port map (
            O => \N__64166\,
            I => \N__64075\
        );

    \I__15787\ : LocalMux
    port map (
            O => \N__64161\,
            I => \N__64061\
        );

    \I__15786\ : LocalMux
    port map (
            O => \N__64158\,
            I => \N__64061\
        );

    \I__15785\ : InMux
    port map (
            O => \N__64157\,
            I => \N__64058\
        );

    \I__15784\ : Span4Mux_h
    port map (
            O => \N__64154\,
            I => \N__64055\
        );

    \I__15783\ : InMux
    port map (
            O => \N__64153\,
            I => \N__64050\
        );

    \I__15782\ : InMux
    port map (
            O => \N__64152\,
            I => \N__64050\
        );

    \I__15781\ : LocalMux
    port map (
            O => \N__64149\,
            I => \N__64043\
        );

    \I__15780\ : LocalMux
    port map (
            O => \N__64144\,
            I => \N__64043\
        );

    \I__15779\ : Span4Mux_v
    port map (
            O => \N__64139\,
            I => \N__64043\
        );

    \I__15778\ : LocalMux
    port map (
            O => \N__64124\,
            I => \N__64038\
        );

    \I__15777\ : Span4Mux_v
    port map (
            O => \N__64121\,
            I => \N__64038\
        );

    \I__15776\ : InMux
    port map (
            O => \N__64118\,
            I => \N__64033\
        );

    \I__15775\ : InMux
    port map (
            O => \N__64117\,
            I => \N__64033\
        );

    \I__15774\ : LocalMux
    port map (
            O => \N__64100\,
            I => \N__64028\
        );

    \I__15773\ : Span4Mux_v
    port map (
            O => \N__64095\,
            I => \N__64028\
        );

    \I__15772\ : Span4Mux_h
    port map (
            O => \N__64092\,
            I => \N__64021\
        );

    \I__15771\ : Span4Mux_v
    port map (
            O => \N__64089\,
            I => \N__64021\
        );

    \I__15770\ : LocalMux
    port map (
            O => \N__64082\,
            I => \N__64021\
        );

    \I__15769\ : InMux
    port map (
            O => \N__64081\,
            I => \N__64018\
        );

    \I__15768\ : Span4Mux_h
    port map (
            O => \N__64078\,
            I => \N__64013\
        );

    \I__15767\ : Span4Mux_h
    port map (
            O => \N__64075\,
            I => \N__64013\
        );

    \I__15766\ : InMux
    port map (
            O => \N__64074\,
            I => \N__64010\
        );

    \I__15765\ : InMux
    port map (
            O => \N__64073\,
            I => \N__64007\
        );

    \I__15764\ : InMux
    port map (
            O => \N__64072\,
            I => \N__64000\
        );

    \I__15763\ : InMux
    port map (
            O => \N__64071\,
            I => \N__64000\
        );

    \I__15762\ : InMux
    port map (
            O => \N__64070\,
            I => \N__64000\
        );

    \I__15761\ : InMux
    port map (
            O => \N__64069\,
            I => \N__63991\
        );

    \I__15760\ : InMux
    port map (
            O => \N__64068\,
            I => \N__63991\
        );

    \I__15759\ : InMux
    port map (
            O => \N__64067\,
            I => \N__63991\
        );

    \I__15758\ : InMux
    port map (
            O => \N__64066\,
            I => \N__63991\
        );

    \I__15757\ : Span4Mux_v
    port map (
            O => \N__64061\,
            I => \N__63988\
        );

    \I__15756\ : LocalMux
    port map (
            O => \N__64058\,
            I => \N__63977\
        );

    \I__15755\ : Span4Mux_v
    port map (
            O => \N__64055\,
            I => \N__63977\
        );

    \I__15754\ : LocalMux
    port map (
            O => \N__64050\,
            I => \N__63977\
        );

    \I__15753\ : Span4Mux_h
    port map (
            O => \N__64043\,
            I => \N__63977\
        );

    \I__15752\ : Span4Mux_v
    port map (
            O => \N__64038\,
            I => \N__63977\
        );

    \I__15751\ : LocalMux
    port map (
            O => \N__64033\,
            I => \N__63970\
        );

    \I__15750\ : Span4Mux_h
    port map (
            O => \N__64028\,
            I => \N__63970\
        );

    \I__15749\ : Span4Mux_v
    port map (
            O => \N__64021\,
            I => \N__63970\
        );

    \I__15748\ : LocalMux
    port map (
            O => \N__64018\,
            I => \N_1838_0\
        );

    \I__15747\ : Odrv4
    port map (
            O => \N__64013\,
            I => \N_1838_0\
        );

    \I__15746\ : LocalMux
    port map (
            O => \N__64010\,
            I => \N_1838_0\
        );

    \I__15745\ : LocalMux
    port map (
            O => \N__64007\,
            I => \N_1838_0\
        );

    \I__15744\ : LocalMux
    port map (
            O => \N__64000\,
            I => \N_1838_0\
        );

    \I__15743\ : LocalMux
    port map (
            O => \N__63991\,
            I => \N_1838_0\
        );

    \I__15742\ : Odrv4
    port map (
            O => \N__63988\,
            I => \N_1838_0\
        );

    \I__15741\ : Odrv4
    port map (
            O => \N__63977\,
            I => \N_1838_0\
        );

    \I__15740\ : Odrv4
    port map (
            O => \N__63970\,
            I => \N_1838_0\
        );

    \I__15739\ : InMux
    port map (
            O => \N__63951\,
            I => \N__63948\
        );

    \I__15738\ : LocalMux
    port map (
            O => \N__63948\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_2\
        );

    \I__15737\ : InMux
    port map (
            O => \N__63945\,
            I => \N__63941\
        );

    \I__15736\ : InMux
    port map (
            O => \N__63944\,
            I => \N__63936\
        );

    \I__15735\ : LocalMux
    port map (
            O => \N__63941\,
            I => \N__63933\
        );

    \I__15734\ : InMux
    port map (
            O => \N__63940\,
            I => \N__63930\
        );

    \I__15733\ : InMux
    port map (
            O => \N__63939\,
            I => \N__63927\
        );

    \I__15732\ : LocalMux
    port map (
            O => \N__63936\,
            I => \N__63924\
        );

    \I__15731\ : Span4Mux_v
    port map (
            O => \N__63933\,
            I => \N__63918\
        );

    \I__15730\ : LocalMux
    port map (
            O => \N__63930\,
            I => \N__63918\
        );

    \I__15729\ : LocalMux
    port map (
            O => \N__63927\,
            I => \N__63915\
        );

    \I__15728\ : Span4Mux_v
    port map (
            O => \N__63924\,
            I => \N__63911\
        );

    \I__15727\ : InMux
    port map (
            O => \N__63923\,
            I => \N__63906\
        );

    \I__15726\ : Span4Mux_v
    port map (
            O => \N__63918\,
            I => \N__63902\
        );

    \I__15725\ : Span4Mux_v
    port map (
            O => \N__63915\,
            I => \N__63899\
        );

    \I__15724\ : InMux
    port map (
            O => \N__63914\,
            I => \N__63896\
        );

    \I__15723\ : Span4Mux_v
    port map (
            O => \N__63911\,
            I => \N__63893\
        );

    \I__15722\ : InMux
    port map (
            O => \N__63910\,
            I => \N__63890\
        );

    \I__15721\ : InMux
    port map (
            O => \N__63909\,
            I => \N__63887\
        );

    \I__15720\ : LocalMux
    port map (
            O => \N__63906\,
            I => \N__63884\
        );

    \I__15719\ : InMux
    port map (
            O => \N__63905\,
            I => \N__63881\
        );

    \I__15718\ : Span4Mux_h
    port map (
            O => \N__63902\,
            I => \N__63878\
        );

    \I__15717\ : Span4Mux_h
    port map (
            O => \N__63899\,
            I => \N__63873\
        );

    \I__15716\ : LocalMux
    port map (
            O => \N__63896\,
            I => \N__63873\
        );

    \I__15715\ : Sp12to4
    port map (
            O => \N__63893\,
            I => \N__63870\
        );

    \I__15714\ : LocalMux
    port map (
            O => \N__63890\,
            I => \N__63867\
        );

    \I__15713\ : LocalMux
    port map (
            O => \N__63887\,
            I => \N__63864\
        );

    \I__15712\ : Span4Mux_v
    port map (
            O => \N__63884\,
            I => \N__63859\
        );

    \I__15711\ : LocalMux
    port map (
            O => \N__63881\,
            I => \N__63859\
        );

    \I__15710\ : Span4Mux_h
    port map (
            O => \N__63878\,
            I => \N__63854\
        );

    \I__15709\ : Span4Mux_v
    port map (
            O => \N__63873\,
            I => \N__63854\
        );

    \I__15708\ : Span12Mux_h
    port map (
            O => \N__63870\,
            I => \N__63851\
        );

    \I__15707\ : Span4Mux_v
    port map (
            O => \N__63867\,
            I => \N__63844\
        );

    \I__15706\ : Span4Mux_v
    port map (
            O => \N__63864\,
            I => \N__63844\
        );

    \I__15705\ : Span4Mux_h
    port map (
            O => \N__63859\,
            I => \N__63844\
        );

    \I__15704\ : Odrv4
    port map (
            O => \N__63854\,
            I => \I2C_top_level_inst1_s_data_oreg_3\
        );

    \I__15703\ : Odrv12
    port map (
            O => \N__63851\,
            I => \I2C_top_level_inst1_s_data_oreg_3\
        );

    \I__15702\ : Odrv4
    port map (
            O => \N__63844\,
            I => \I2C_top_level_inst1_s_data_oreg_3\
        );

    \I__15701\ : InMux
    port map (
            O => \N__63837\,
            I => \N__63834\
        );

    \I__15700\ : LocalMux
    port map (
            O => \N__63834\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_3\
        );

    \I__15699\ : CascadeMux
    port map (
            O => \N__63831\,
            I => \N__63828\
        );

    \I__15698\ : InMux
    port map (
            O => \N__63828\,
            I => \N__63823\
        );

    \I__15697\ : InMux
    port map (
            O => \N__63827\,
            I => \N__63819\
        );

    \I__15696\ : InMux
    port map (
            O => \N__63826\,
            I => \N__63816\
        );

    \I__15695\ : LocalMux
    port map (
            O => \N__63823\,
            I => \N__63813\
        );

    \I__15694\ : InMux
    port map (
            O => \N__63822\,
            I => \N__63810\
        );

    \I__15693\ : LocalMux
    port map (
            O => \N__63819\,
            I => \N__63806\
        );

    \I__15692\ : LocalMux
    port map (
            O => \N__63816\,
            I => \N__63803\
        );

    \I__15691\ : Span4Mux_v
    port map (
            O => \N__63813\,
            I => \N__63800\
        );

    \I__15690\ : LocalMux
    port map (
            O => \N__63810\,
            I => \N__63796\
        );

    \I__15689\ : InMux
    port map (
            O => \N__63809\,
            I => \N__63793\
        );

    \I__15688\ : Span4Mux_v
    port map (
            O => \N__63806\,
            I => \N__63790\
        );

    \I__15687\ : Span4Mux_h
    port map (
            O => \N__63803\,
            I => \N__63786\
        );

    \I__15686\ : Span4Mux_h
    port map (
            O => \N__63800\,
            I => \N__63782\
        );

    \I__15685\ : InMux
    port map (
            O => \N__63799\,
            I => \N__63779\
        );

    \I__15684\ : Span4Mux_h
    port map (
            O => \N__63796\,
            I => \N__63776\
        );

    \I__15683\ : LocalMux
    port map (
            O => \N__63793\,
            I => \N__63770\
        );

    \I__15682\ : Span4Mux_h
    port map (
            O => \N__63790\,
            I => \N__63770\
        );

    \I__15681\ : InMux
    port map (
            O => \N__63789\,
            I => \N__63767\
        );

    \I__15680\ : Sp12to4
    port map (
            O => \N__63786\,
            I => \N__63764\
        );

    \I__15679\ : InMux
    port map (
            O => \N__63785\,
            I => \N__63761\
        );

    \I__15678\ : Span4Mux_h
    port map (
            O => \N__63782\,
            I => \N__63756\
        );

    \I__15677\ : LocalMux
    port map (
            O => \N__63779\,
            I => \N__63756\
        );

    \I__15676\ : Span4Mux_h
    port map (
            O => \N__63776\,
            I => \N__63753\
        );

    \I__15675\ : InMux
    port map (
            O => \N__63775\,
            I => \N__63750\
        );

    \I__15674\ : Span4Mux_v
    port map (
            O => \N__63770\,
            I => \N__63747\
        );

    \I__15673\ : LocalMux
    port map (
            O => \N__63767\,
            I => \N__63742\
        );

    \I__15672\ : Span12Mux_v
    port map (
            O => \N__63764\,
            I => \N__63742\
        );

    \I__15671\ : LocalMux
    port map (
            O => \N__63761\,
            I => \N__63739\
        );

    \I__15670\ : Span4Mux_v
    port map (
            O => \N__63756\,
            I => \N__63736\
        );

    \I__15669\ : Span4Mux_v
    port map (
            O => \N__63753\,
            I => \N__63733\
        );

    \I__15668\ : LocalMux
    port map (
            O => \N__63750\,
            I => \N__63730\
        );

    \I__15667\ : Span4Mux_h
    port map (
            O => \N__63747\,
            I => \N__63727\
        );

    \I__15666\ : Span12Mux_h
    port map (
            O => \N__63742\,
            I => \N__63724\
        );

    \I__15665\ : Span4Mux_v
    port map (
            O => \N__63739\,
            I => \N__63719\
        );

    \I__15664\ : Span4Mux_v
    port map (
            O => \N__63736\,
            I => \N__63719\
        );

    \I__15663\ : Odrv4
    port map (
            O => \N__63733\,
            I => \I2C_top_level_inst1_s_data_oreg_4\
        );

    \I__15662\ : Odrv4
    port map (
            O => \N__63730\,
            I => \I2C_top_level_inst1_s_data_oreg_4\
        );

    \I__15661\ : Odrv4
    port map (
            O => \N__63727\,
            I => \I2C_top_level_inst1_s_data_oreg_4\
        );

    \I__15660\ : Odrv12
    port map (
            O => \N__63724\,
            I => \I2C_top_level_inst1_s_data_oreg_4\
        );

    \I__15659\ : Odrv4
    port map (
            O => \N__63719\,
            I => \I2C_top_level_inst1_s_data_oreg_4\
        );

    \I__15658\ : InMux
    port map (
            O => \N__63708\,
            I => \N__63705\
        );

    \I__15657\ : LocalMux
    port map (
            O => \N__63705\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_4\
        );

    \I__15656\ : InMux
    port map (
            O => \N__63702\,
            I => \N__63698\
        );

    \I__15655\ : InMux
    port map (
            O => \N__63701\,
            I => \N__63694\
        );

    \I__15654\ : LocalMux
    port map (
            O => \N__63698\,
            I => \N__63691\
        );

    \I__15653\ : CascadeMux
    port map (
            O => \N__63697\,
            I => \N__63688\
        );

    \I__15652\ : LocalMux
    port map (
            O => \N__63694\,
            I => \N__63684\
        );

    \I__15651\ : Span4Mux_v
    port map (
            O => \N__63691\,
            I => \N__63681\
        );

    \I__15650\ : InMux
    port map (
            O => \N__63688\,
            I => \N__63678\
        );

    \I__15649\ : InMux
    port map (
            O => \N__63687\,
            I => \N__63674\
        );

    \I__15648\ : Span4Mux_h
    port map (
            O => \N__63684\,
            I => \N__63671\
        );

    \I__15647\ : Span4Mux_h
    port map (
            O => \N__63681\,
            I => \N__63665\
        );

    \I__15646\ : LocalMux
    port map (
            O => \N__63678\,
            I => \N__63665\
        );

    \I__15645\ : InMux
    port map (
            O => \N__63677\,
            I => \N__63662\
        );

    \I__15644\ : LocalMux
    port map (
            O => \N__63674\,
            I => \N__63658\
        );

    \I__15643\ : Span4Mux_v
    port map (
            O => \N__63671\,
            I => \N__63654\
        );

    \I__15642\ : CascadeMux
    port map (
            O => \N__63670\,
            I => \N__63651\
        );

    \I__15641\ : Span4Mux_v
    port map (
            O => \N__63665\,
            I => \N__63646\
        );

    \I__15640\ : LocalMux
    port map (
            O => \N__63662\,
            I => \N__63646\
        );

    \I__15639\ : InMux
    port map (
            O => \N__63661\,
            I => \N__63642\
        );

    \I__15638\ : Span4Mux_v
    port map (
            O => \N__63658\,
            I => \N__63639\
        );

    \I__15637\ : InMux
    port map (
            O => \N__63657\,
            I => \N__63636\
        );

    \I__15636\ : Sp12to4
    port map (
            O => \N__63654\,
            I => \N__63633\
        );

    \I__15635\ : InMux
    port map (
            O => \N__63651\,
            I => \N__63630\
        );

    \I__15634\ : Span4Mux_h
    port map (
            O => \N__63646\,
            I => \N__63627\
        );

    \I__15633\ : InMux
    port map (
            O => \N__63645\,
            I => \N__63624\
        );

    \I__15632\ : LocalMux
    port map (
            O => \N__63642\,
            I => \N__63621\
        );

    \I__15631\ : Sp12to4
    port map (
            O => \N__63639\,
            I => \N__63612\
        );

    \I__15630\ : LocalMux
    port map (
            O => \N__63636\,
            I => \N__63612\
        );

    \I__15629\ : Span12Mux_v
    port map (
            O => \N__63633\,
            I => \N__63612\
        );

    \I__15628\ : LocalMux
    port map (
            O => \N__63630\,
            I => \N__63612\
        );

    \I__15627\ : Span4Mux_h
    port map (
            O => \N__63627\,
            I => \N__63609\
        );

    \I__15626\ : LocalMux
    port map (
            O => \N__63624\,
            I => \N__63606\
        );

    \I__15625\ : Span4Mux_h
    port map (
            O => \N__63621\,
            I => \N__63603\
        );

    \I__15624\ : Span12Mux_h
    port map (
            O => \N__63612\,
            I => \N__63600\
        );

    \I__15623\ : Odrv4
    port map (
            O => \N__63609\,
            I => \I2C_top_level_inst1_s_data_oreg_5\
        );

    \I__15622\ : Odrv12
    port map (
            O => \N__63606\,
            I => \I2C_top_level_inst1_s_data_oreg_5\
        );

    \I__15621\ : Odrv4
    port map (
            O => \N__63603\,
            I => \I2C_top_level_inst1_s_data_oreg_5\
        );

    \I__15620\ : Odrv12
    port map (
            O => \N__63600\,
            I => \I2C_top_level_inst1_s_data_oreg_5\
        );

    \I__15619\ : InMux
    port map (
            O => \N__63591\,
            I => \N__63588\
        );

    \I__15618\ : LocalMux
    port map (
            O => \N__63588\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_5\
        );

    \I__15617\ : InMux
    port map (
            O => \N__63585\,
            I => \N__63577\
        );

    \I__15616\ : InMux
    port map (
            O => \N__63584\,
            I => \N__63574\
        );

    \I__15615\ : InMux
    port map (
            O => \N__63583\,
            I => \N__63569\
        );

    \I__15614\ : InMux
    port map (
            O => \N__63582\,
            I => \N__63569\
        );

    \I__15613\ : InMux
    port map (
            O => \N__63581\,
            I => \N__63565\
        );

    \I__15612\ : InMux
    port map (
            O => \N__63580\,
            I => \N__63562\
        );

    \I__15611\ : LocalMux
    port map (
            O => \N__63577\,
            I => \N__63559\
        );

    \I__15610\ : LocalMux
    port map (
            O => \N__63574\,
            I => \N__63556\
        );

    \I__15609\ : LocalMux
    port map (
            O => \N__63569\,
            I => \N__63553\
        );

    \I__15608\ : InMux
    port map (
            O => \N__63568\,
            I => \N__63550\
        );

    \I__15607\ : LocalMux
    port map (
            O => \N__63565\,
            I => \N__63547\
        );

    \I__15606\ : LocalMux
    port map (
            O => \N__63562\,
            I => \N__63544\
        );

    \I__15605\ : Span4Mux_v
    port map (
            O => \N__63559\,
            I => \N__63540\
        );

    \I__15604\ : Span4Mux_v
    port map (
            O => \N__63556\,
            I => \N__63537\
        );

    \I__15603\ : Span4Mux_h
    port map (
            O => \N__63553\,
            I => \N__63532\
        );

    \I__15602\ : LocalMux
    port map (
            O => \N__63550\,
            I => \N__63532\
        );

    \I__15601\ : Span4Mux_h
    port map (
            O => \N__63547\,
            I => \N__63527\
        );

    \I__15600\ : Span4Mux_v
    port map (
            O => \N__63544\,
            I => \N__63527\
        );

    \I__15599\ : InMux
    port map (
            O => \N__63543\,
            I => \N__63523\
        );

    \I__15598\ : Sp12to4
    port map (
            O => \N__63540\,
            I => \N__63520\
        );

    \I__15597\ : Span4Mux_h
    port map (
            O => \N__63537\,
            I => \N__63517\
        );

    \I__15596\ : Span4Mux_h
    port map (
            O => \N__63532\,
            I => \N__63514\
        );

    \I__15595\ : Span4Mux_h
    port map (
            O => \N__63527\,
            I => \N__63511\
        );

    \I__15594\ : InMux
    port map (
            O => \N__63526\,
            I => \N__63508\
        );

    \I__15593\ : LocalMux
    port map (
            O => \N__63523\,
            I => \N__63503\
        );

    \I__15592\ : Span12Mux_h
    port map (
            O => \N__63520\,
            I => \N__63503\
        );

    \I__15591\ : Span4Mux_v
    port map (
            O => \N__63517\,
            I => \N__63498\
        );

    \I__15590\ : Span4Mux_v
    port map (
            O => \N__63514\,
            I => \N__63498\
        );

    \I__15589\ : Odrv4
    port map (
            O => \N__63511\,
            I => \I2C_top_level_inst1_s_data_oreg_6\
        );

    \I__15588\ : LocalMux
    port map (
            O => \N__63508\,
            I => \I2C_top_level_inst1_s_data_oreg_6\
        );

    \I__15587\ : Odrv12
    port map (
            O => \N__63503\,
            I => \I2C_top_level_inst1_s_data_oreg_6\
        );

    \I__15586\ : Odrv4
    port map (
            O => \N__63498\,
            I => \I2C_top_level_inst1_s_data_oreg_6\
        );

    \I__15585\ : InMux
    port map (
            O => \N__63489\,
            I => \N__63486\
        );

    \I__15584\ : LocalMux
    port map (
            O => \N__63486\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_6\
        );

    \I__15583\ : InMux
    port map (
            O => \N__63483\,
            I => \N__63478\
        );

    \I__15582\ : InMux
    port map (
            O => \N__63482\,
            I => \N__63473\
        );

    \I__15581\ : InMux
    port map (
            O => \N__63481\,
            I => \N__63468\
        );

    \I__15580\ : LocalMux
    port map (
            O => \N__63478\,
            I => \N__63464\
        );

    \I__15579\ : InMux
    port map (
            O => \N__63477\,
            I => \N__63461\
        );

    \I__15578\ : InMux
    port map (
            O => \N__63476\,
            I => \N__63458\
        );

    \I__15577\ : LocalMux
    port map (
            O => \N__63473\,
            I => \N__63455\
        );

    \I__15576\ : CascadeMux
    port map (
            O => \N__63472\,
            I => \N__63452\
        );

    \I__15575\ : InMux
    port map (
            O => \N__63471\,
            I => \N__63449\
        );

    \I__15574\ : LocalMux
    port map (
            O => \N__63468\,
            I => \N__63445\
        );

    \I__15573\ : InMux
    port map (
            O => \N__63467\,
            I => \N__63442\
        );

    \I__15572\ : Span4Mux_v
    port map (
            O => \N__63464\,
            I => \N__63439\
        );

    \I__15571\ : LocalMux
    port map (
            O => \N__63461\,
            I => \N__63436\
        );

    \I__15570\ : LocalMux
    port map (
            O => \N__63458\,
            I => \N__63433\
        );

    \I__15569\ : Span4Mux_v
    port map (
            O => \N__63455\,
            I => \N__63430\
        );

    \I__15568\ : InMux
    port map (
            O => \N__63452\,
            I => \N__63427\
        );

    \I__15567\ : LocalMux
    port map (
            O => \N__63449\,
            I => \N__63424\
        );

    \I__15566\ : InMux
    port map (
            O => \N__63448\,
            I => \N__63421\
        );

    \I__15565\ : Span4Mux_v
    port map (
            O => \N__63445\,
            I => \N__63418\
        );

    \I__15564\ : LocalMux
    port map (
            O => \N__63442\,
            I => \N__63407\
        );

    \I__15563\ : Sp12to4
    port map (
            O => \N__63439\,
            I => \N__63407\
        );

    \I__15562\ : Span12Mux_v
    port map (
            O => \N__63436\,
            I => \N__63407\
        );

    \I__15561\ : Sp12to4
    port map (
            O => \N__63433\,
            I => \N__63407\
        );

    \I__15560\ : Sp12to4
    port map (
            O => \N__63430\,
            I => \N__63407\
        );

    \I__15559\ : LocalMux
    port map (
            O => \N__63427\,
            I => \N__63400\
        );

    \I__15558\ : Span12Mux_v
    port map (
            O => \N__63424\,
            I => \N__63400\
        );

    \I__15557\ : LocalMux
    port map (
            O => \N__63421\,
            I => \N__63400\
        );

    \I__15556\ : Span4Mux_h
    port map (
            O => \N__63418\,
            I => \N__63397\
        );

    \I__15555\ : Span12Mux_h
    port map (
            O => \N__63407\,
            I => \N__63394\
        );

    \I__15554\ : Span12Mux_h
    port map (
            O => \N__63400\,
            I => \N__63391\
        );

    \I__15553\ : Odrv4
    port map (
            O => \N__63397\,
            I => \I2C_top_level_inst1_s_data_oreg_7\
        );

    \I__15552\ : Odrv12
    port map (
            O => \N__63394\,
            I => \I2C_top_level_inst1_s_data_oreg_7\
        );

    \I__15551\ : Odrv12
    port map (
            O => \N__63391\,
            I => \I2C_top_level_inst1_s_data_oreg_7\
        );

    \I__15550\ : InMux
    port map (
            O => \N__63384\,
            I => \N__63359\
        );

    \I__15549\ : InMux
    port map (
            O => \N__63383\,
            I => \N__63359\
        );

    \I__15548\ : InMux
    port map (
            O => \N__63382\,
            I => \N__63359\
        );

    \I__15547\ : InMux
    port map (
            O => \N__63381\,
            I => \N__63359\
        );

    \I__15546\ : InMux
    port map (
            O => \N__63380\,
            I => \N__63359\
        );

    \I__15545\ : InMux
    port map (
            O => \N__63379\,
            I => \N__63359\
        );

    \I__15544\ : InMux
    port map (
            O => \N__63378\,
            I => \N__63359\
        );

    \I__15543\ : InMux
    port map (
            O => \N__63377\,
            I => \N__63359\
        );

    \I__15542\ : CascadeMux
    port map (
            O => \N__63376\,
            I => \N__63356\
        );

    \I__15541\ : LocalMux
    port map (
            O => \N__63359\,
            I => \N__63338\
        );

    \I__15540\ : InMux
    port map (
            O => \N__63356\,
            I => \N__63327\
        );

    \I__15539\ : InMux
    port map (
            O => \N__63355\,
            I => \N__63327\
        );

    \I__15538\ : InMux
    port map (
            O => \N__63354\,
            I => \N__63327\
        );

    \I__15537\ : InMux
    port map (
            O => \N__63353\,
            I => \N__63327\
        );

    \I__15536\ : InMux
    port map (
            O => \N__63352\,
            I => \N__63327\
        );

    \I__15535\ : InMux
    port map (
            O => \N__63351\,
            I => \N__63310\
        );

    \I__15534\ : InMux
    port map (
            O => \N__63350\,
            I => \N__63310\
        );

    \I__15533\ : InMux
    port map (
            O => \N__63349\,
            I => \N__63310\
        );

    \I__15532\ : InMux
    port map (
            O => \N__63348\,
            I => \N__63310\
        );

    \I__15531\ : InMux
    port map (
            O => \N__63347\,
            I => \N__63310\
        );

    \I__15530\ : InMux
    port map (
            O => \N__63346\,
            I => \N__63310\
        );

    \I__15529\ : InMux
    port map (
            O => \N__63345\,
            I => \N__63310\
        );

    \I__15528\ : InMux
    port map (
            O => \N__63344\,
            I => \N__63310\
        );

    \I__15527\ : InMux
    port map (
            O => \N__63343\,
            I => \N__63303\
        );

    \I__15526\ : InMux
    port map (
            O => \N__63342\,
            I => \N__63303\
        );

    \I__15525\ : InMux
    port map (
            O => \N__63341\,
            I => \N__63303\
        );

    \I__15524\ : Span4Mux_v
    port map (
            O => \N__63338\,
            I => \N__63285\
        );

    \I__15523\ : LocalMux
    port map (
            O => \N__63327\,
            I => \N__63285\
        );

    \I__15522\ : LocalMux
    port map (
            O => \N__63310\,
            I => \N__63285\
        );

    \I__15521\ : LocalMux
    port map (
            O => \N__63303\,
            I => \N__63282\
        );

    \I__15520\ : CascadeMux
    port map (
            O => \N__63302\,
            I => \N__63278\
        );

    \I__15519\ : CascadeMux
    port map (
            O => \N__63301\,
            I => \N__63275\
        );

    \I__15518\ : InMux
    port map (
            O => \N__63300\,
            I => \N__63270\
        );

    \I__15517\ : InMux
    port map (
            O => \N__63299\,
            I => \N__63255\
        );

    \I__15516\ : InMux
    port map (
            O => \N__63298\,
            I => \N__63255\
        );

    \I__15515\ : InMux
    port map (
            O => \N__63297\,
            I => \N__63255\
        );

    \I__15514\ : InMux
    port map (
            O => \N__63296\,
            I => \N__63255\
        );

    \I__15513\ : InMux
    port map (
            O => \N__63295\,
            I => \N__63255\
        );

    \I__15512\ : InMux
    port map (
            O => \N__63294\,
            I => \N__63255\
        );

    \I__15511\ : InMux
    port map (
            O => \N__63293\,
            I => \N__63255\
        );

    \I__15510\ : InMux
    port map (
            O => \N__63292\,
            I => \N__63252\
        );

    \I__15509\ : Span4Mux_v
    port map (
            O => \N__63285\,
            I => \N__63247\
        );

    \I__15508\ : Span4Mux_v
    port map (
            O => \N__63282\,
            I => \N__63247\
        );

    \I__15507\ : InMux
    port map (
            O => \N__63281\,
            I => \N__63243\
        );

    \I__15506\ : InMux
    port map (
            O => \N__63278\,
            I => \N__63238\
        );

    \I__15505\ : InMux
    port map (
            O => \N__63275\,
            I => \N__63238\
        );

    \I__15504\ : CascadeMux
    port map (
            O => \N__63274\,
            I => \N__63235\
        );

    \I__15503\ : CascadeMux
    port map (
            O => \N__63273\,
            I => \N__63232\
        );

    \I__15502\ : LocalMux
    port map (
            O => \N__63270\,
            I => \N__63225\
        );

    \I__15501\ : LocalMux
    port map (
            O => \N__63255\,
            I => \N__63225\
        );

    \I__15500\ : LocalMux
    port map (
            O => \N__63252\,
            I => \N__63222\
        );

    \I__15499\ : Span4Mux_h
    port map (
            O => \N__63247\,
            I => \N__63219\
        );

    \I__15498\ : InMux
    port map (
            O => \N__63246\,
            I => \N__63216\
        );

    \I__15497\ : LocalMux
    port map (
            O => \N__63243\,
            I => \N__63211\
        );

    \I__15496\ : LocalMux
    port map (
            O => \N__63238\,
            I => \N__63211\
        );

    \I__15495\ : InMux
    port map (
            O => \N__63235\,
            I => \N__63202\
        );

    \I__15494\ : InMux
    port map (
            O => \N__63232\,
            I => \N__63202\
        );

    \I__15493\ : InMux
    port map (
            O => \N__63231\,
            I => \N__63202\
        );

    \I__15492\ : InMux
    port map (
            O => \N__63230\,
            I => \N__63202\
        );

    \I__15491\ : Span4Mux_h
    port map (
            O => \N__63225\,
            I => \N__63199\
        );

    \I__15490\ : Span4Mux_v
    port map (
            O => \N__63222\,
            I => \N__63194\
        );

    \I__15489\ : Sp12to4
    port map (
            O => \N__63219\,
            I => \N__63191\
        );

    \I__15488\ : LocalMux
    port map (
            O => \N__63216\,
            I => \N__63188\
        );

    \I__15487\ : Span4Mux_h
    port map (
            O => \N__63211\,
            I => \N__63183\
        );

    \I__15486\ : LocalMux
    port map (
            O => \N__63202\,
            I => \N__63183\
        );

    \I__15485\ : Span4Mux_v
    port map (
            O => \N__63199\,
            I => \N__63180\
        );

    \I__15484\ : InMux
    port map (
            O => \N__63198\,
            I => \N__63175\
        );

    \I__15483\ : InMux
    port map (
            O => \N__63197\,
            I => \N__63175\
        );

    \I__15482\ : Sp12to4
    port map (
            O => \N__63194\,
            I => \N__63170\
        );

    \I__15481\ : Span12Mux_v
    port map (
            O => \N__63191\,
            I => \N__63170\
        );

    \I__15480\ : Span4Mux_v
    port map (
            O => \N__63188\,
            I => \N__63163\
        );

    \I__15479\ : Span4Mux_v
    port map (
            O => \N__63183\,
            I => \N__63163\
        );

    \I__15478\ : Span4Mux_h
    port map (
            O => \N__63180\,
            I => \N__63163\
        );

    \I__15477\ : LocalMux
    port map (
            O => \N__63175\,
            I => \I2C_top_level_inst1.s_enable_desp_tx\
        );

    \I__15476\ : Odrv12
    port map (
            O => \N__63170\,
            I => \I2C_top_level_inst1.s_enable_desp_tx\
        );

    \I__15475\ : Odrv4
    port map (
            O => \N__63163\,
            I => \I2C_top_level_inst1.s_enable_desp_tx\
        );

    \I__15474\ : InMux
    port map (
            O => \N__63156\,
            I => \N__63153\
        );

    \I__15473\ : LocalMux
    port map (
            O => \N__63153\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_7\
        );

    \I__15472\ : InMux
    port map (
            O => \N__63150\,
            I => \N__63146\
        );

    \I__15471\ : InMux
    port map (
            O => \N__63149\,
            I => \N__63141\
        );

    \I__15470\ : LocalMux
    port map (
            O => \N__63146\,
            I => \N__63138\
        );

    \I__15469\ : InMux
    port map (
            O => \N__63145\,
            I => \N__63135\
        );

    \I__15468\ : InMux
    port map (
            O => \N__63144\,
            I => \N__63131\
        );

    \I__15467\ : LocalMux
    port map (
            O => \N__63141\,
            I => \N__63128\
        );

    \I__15466\ : Span4Mux_v
    port map (
            O => \N__63138\,
            I => \N__63123\
        );

    \I__15465\ : LocalMux
    port map (
            O => \N__63135\,
            I => \N__63123\
        );

    \I__15464\ : CascadeMux
    port map (
            O => \N__63134\,
            I => \N__63120\
        );

    \I__15463\ : LocalMux
    port map (
            O => \N__63131\,
            I => \N__63115\
        );

    \I__15462\ : Span4Mux_v
    port map (
            O => \N__63128\,
            I => \N__63110\
        );

    \I__15461\ : Span4Mux_v
    port map (
            O => \N__63123\,
            I => \N__63110\
        );

    \I__15460\ : InMux
    port map (
            O => \N__63120\,
            I => \N__63107\
        );

    \I__15459\ : InMux
    port map (
            O => \N__63119\,
            I => \N__63104\
        );

    \I__15458\ : InMux
    port map (
            O => \N__63118\,
            I => \N__63099\
        );

    \I__15457\ : Span4Mux_v
    port map (
            O => \N__63115\,
            I => \N__63094\
        );

    \I__15456\ : Span4Mux_h
    port map (
            O => \N__63110\,
            I => \N__63094\
        );

    \I__15455\ : LocalMux
    port map (
            O => \N__63107\,
            I => \N__63091\
        );

    \I__15454\ : LocalMux
    port map (
            O => \N__63104\,
            I => \N__63088\
        );

    \I__15453\ : InMux
    port map (
            O => \N__63103\,
            I => \N__63083\
        );

    \I__15452\ : InMux
    port map (
            O => \N__63102\,
            I => \N__63083\
        );

    \I__15451\ : LocalMux
    port map (
            O => \N__63099\,
            I => \N__63080\
        );

    \I__15450\ : Span4Mux_h
    port map (
            O => \N__63094\,
            I => \N__63077\
        );

    \I__15449\ : Span4Mux_h
    port map (
            O => \N__63091\,
            I => \N__63074\
        );

    \I__15448\ : Span4Mux_v
    port map (
            O => \N__63088\,
            I => \N__63071\
        );

    \I__15447\ : LocalMux
    port map (
            O => \N__63083\,
            I => \N__63068\
        );

    \I__15446\ : Span12Mux_v
    port map (
            O => \N__63080\,
            I => \N__63065\
        );

    \I__15445\ : Span4Mux_v
    port map (
            O => \N__63077\,
            I => \N__63062\
        );

    \I__15444\ : Span4Mux_h
    port map (
            O => \N__63074\,
            I => \N__63059\
        );

    \I__15443\ : Span4Mux_h
    port map (
            O => \N__63071\,
            I => \N__63054\
        );

    \I__15442\ : Span4Mux_v
    port map (
            O => \N__63068\,
            I => \N__63054\
        );

    \I__15441\ : Odrv12
    port map (
            O => \N__63065\,
            I => \I2C_top_level_inst1_s_data_oreg_8\
        );

    \I__15440\ : Odrv4
    port map (
            O => \N__63062\,
            I => \I2C_top_level_inst1_s_data_oreg_8\
        );

    \I__15439\ : Odrv4
    port map (
            O => \N__63059\,
            I => \I2C_top_level_inst1_s_data_oreg_8\
        );

    \I__15438\ : Odrv4
    port map (
            O => \N__63054\,
            I => \I2C_top_level_inst1_s_data_oreg_8\
        );

    \I__15437\ : InMux
    port map (
            O => \N__63045\,
            I => \N__63042\
        );

    \I__15436\ : LocalMux
    port map (
            O => \N__63042\,
            I => \N__63039\
        );

    \I__15435\ : Span4Mux_h
    port map (
            O => \N__63039\,
            I => \N__63036\
        );

    \I__15434\ : Span4Mux_h
    port map (
            O => \N__63036\,
            I => \N__63033\
        );

    \I__15433\ : Odrv4
    port map (
            O => \N__63033\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_8\
        );

    \I__15432\ : CEMux
    port map (
            O => \N__63030\,
            I => \N__63026\
        );

    \I__15431\ : CEMux
    port map (
            O => \N__63029\,
            I => \N__63022\
        );

    \I__15430\ : LocalMux
    port map (
            O => \N__63026\,
            I => \N__63019\
        );

    \I__15429\ : CEMux
    port map (
            O => \N__63025\,
            I => \N__63016\
        );

    \I__15428\ : LocalMux
    port map (
            O => \N__63022\,
            I => \N__63012\
        );

    \I__15427\ : Span4Mux_h
    port map (
            O => \N__63019\,
            I => \N__63007\
        );

    \I__15426\ : LocalMux
    port map (
            O => \N__63016\,
            I => \N__63007\
        );

    \I__15425\ : CEMux
    port map (
            O => \N__63015\,
            I => \N__63004\
        );

    \I__15424\ : Span4Mux_v
    port map (
            O => \N__63012\,
            I => \N__62999\
        );

    \I__15423\ : Span4Mux_v
    port map (
            O => \N__63007\,
            I => \N__62994\
        );

    \I__15422\ : LocalMux
    port map (
            O => \N__63004\,
            I => \N__62994\
        );

    \I__15421\ : CEMux
    port map (
            O => \N__63003\,
            I => \N__62991\
        );

    \I__15420\ : CEMux
    port map (
            O => \N__63002\,
            I => \N__62988\
        );

    \I__15419\ : Span4Mux_h
    port map (
            O => \N__62999\,
            I => \N__62985\
        );

    \I__15418\ : Span4Mux_v
    port map (
            O => \N__62994\,
            I => \N__62980\
        );

    \I__15417\ : LocalMux
    port map (
            O => \N__62991\,
            I => \N__62980\
        );

    \I__15416\ : LocalMux
    port map (
            O => \N__62988\,
            I => \N__62977\
        );

    \I__15415\ : Span4Mux_v
    port map (
            O => \N__62985\,
            I => \N__62974\
        );

    \I__15414\ : Span4Mux_h
    port map (
            O => \N__62980\,
            I => \N__62971\
        );

    \I__15413\ : Span4Mux_v
    port map (
            O => \N__62977\,
            I => \N__62968\
        );

    \I__15412\ : Odrv4
    port map (
            O => \N__62974\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0\
        );

    \I__15411\ : Odrv4
    port map (
            O => \N__62971\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0\
        );

    \I__15410\ : Odrv4
    port map (
            O => \N__62968\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0\
        );

    \I__15409\ : SRMux
    port map (
            O => \N__62961\,
            I => \N__62487\
        );

    \I__15408\ : SRMux
    port map (
            O => \N__62960\,
            I => \N__62487\
        );

    \I__15407\ : SRMux
    port map (
            O => \N__62959\,
            I => \N__62487\
        );

    \I__15406\ : SRMux
    port map (
            O => \N__62958\,
            I => \N__62487\
        );

    \I__15405\ : SRMux
    port map (
            O => \N__62957\,
            I => \N__62487\
        );

    \I__15404\ : SRMux
    port map (
            O => \N__62956\,
            I => \N__62487\
        );

    \I__15403\ : SRMux
    port map (
            O => \N__62955\,
            I => \N__62487\
        );

    \I__15402\ : SRMux
    port map (
            O => \N__62954\,
            I => \N__62487\
        );

    \I__15401\ : SRMux
    port map (
            O => \N__62953\,
            I => \N__62487\
        );

    \I__15400\ : SRMux
    port map (
            O => \N__62952\,
            I => \N__62487\
        );

    \I__15399\ : SRMux
    port map (
            O => \N__62951\,
            I => \N__62487\
        );

    \I__15398\ : SRMux
    port map (
            O => \N__62950\,
            I => \N__62487\
        );

    \I__15397\ : SRMux
    port map (
            O => \N__62949\,
            I => \N__62487\
        );

    \I__15396\ : SRMux
    port map (
            O => \N__62948\,
            I => \N__62487\
        );

    \I__15395\ : SRMux
    port map (
            O => \N__62947\,
            I => \N__62487\
        );

    \I__15394\ : SRMux
    port map (
            O => \N__62946\,
            I => \N__62487\
        );

    \I__15393\ : SRMux
    port map (
            O => \N__62945\,
            I => \N__62487\
        );

    \I__15392\ : SRMux
    port map (
            O => \N__62944\,
            I => \N__62487\
        );

    \I__15391\ : SRMux
    port map (
            O => \N__62943\,
            I => \N__62487\
        );

    \I__15390\ : SRMux
    port map (
            O => \N__62942\,
            I => \N__62487\
        );

    \I__15389\ : SRMux
    port map (
            O => \N__62941\,
            I => \N__62487\
        );

    \I__15388\ : SRMux
    port map (
            O => \N__62940\,
            I => \N__62487\
        );

    \I__15387\ : SRMux
    port map (
            O => \N__62939\,
            I => \N__62487\
        );

    \I__15386\ : SRMux
    port map (
            O => \N__62938\,
            I => \N__62487\
        );

    \I__15385\ : SRMux
    port map (
            O => \N__62937\,
            I => \N__62487\
        );

    \I__15384\ : SRMux
    port map (
            O => \N__62936\,
            I => \N__62487\
        );

    \I__15383\ : SRMux
    port map (
            O => \N__62935\,
            I => \N__62487\
        );

    \I__15382\ : SRMux
    port map (
            O => \N__62934\,
            I => \N__62487\
        );

    \I__15381\ : SRMux
    port map (
            O => \N__62933\,
            I => \N__62487\
        );

    \I__15380\ : SRMux
    port map (
            O => \N__62932\,
            I => \N__62487\
        );

    \I__15379\ : SRMux
    port map (
            O => \N__62931\,
            I => \N__62487\
        );

    \I__15378\ : SRMux
    port map (
            O => \N__62930\,
            I => \N__62487\
        );

    \I__15377\ : SRMux
    port map (
            O => \N__62929\,
            I => \N__62487\
        );

    \I__15376\ : SRMux
    port map (
            O => \N__62928\,
            I => \N__62487\
        );

    \I__15375\ : SRMux
    port map (
            O => \N__62927\,
            I => \N__62487\
        );

    \I__15374\ : SRMux
    port map (
            O => \N__62926\,
            I => \N__62487\
        );

    \I__15373\ : SRMux
    port map (
            O => \N__62925\,
            I => \N__62487\
        );

    \I__15372\ : SRMux
    port map (
            O => \N__62924\,
            I => \N__62487\
        );

    \I__15371\ : SRMux
    port map (
            O => \N__62923\,
            I => \N__62487\
        );

    \I__15370\ : SRMux
    port map (
            O => \N__62922\,
            I => \N__62487\
        );

    \I__15369\ : SRMux
    port map (
            O => \N__62921\,
            I => \N__62487\
        );

    \I__15368\ : SRMux
    port map (
            O => \N__62920\,
            I => \N__62487\
        );

    \I__15367\ : SRMux
    port map (
            O => \N__62919\,
            I => \N__62487\
        );

    \I__15366\ : SRMux
    port map (
            O => \N__62918\,
            I => \N__62487\
        );

    \I__15365\ : SRMux
    port map (
            O => \N__62917\,
            I => \N__62487\
        );

    \I__15364\ : SRMux
    port map (
            O => \N__62916\,
            I => \N__62487\
        );

    \I__15363\ : SRMux
    port map (
            O => \N__62915\,
            I => \N__62487\
        );

    \I__15362\ : SRMux
    port map (
            O => \N__62914\,
            I => \N__62487\
        );

    \I__15361\ : SRMux
    port map (
            O => \N__62913\,
            I => \N__62487\
        );

    \I__15360\ : SRMux
    port map (
            O => \N__62912\,
            I => \N__62487\
        );

    \I__15359\ : SRMux
    port map (
            O => \N__62911\,
            I => \N__62487\
        );

    \I__15358\ : SRMux
    port map (
            O => \N__62910\,
            I => \N__62487\
        );

    \I__15357\ : SRMux
    port map (
            O => \N__62909\,
            I => \N__62487\
        );

    \I__15356\ : SRMux
    port map (
            O => \N__62908\,
            I => \N__62487\
        );

    \I__15355\ : SRMux
    port map (
            O => \N__62907\,
            I => \N__62487\
        );

    \I__15354\ : SRMux
    port map (
            O => \N__62906\,
            I => \N__62487\
        );

    \I__15353\ : SRMux
    port map (
            O => \N__62905\,
            I => \N__62487\
        );

    \I__15352\ : SRMux
    port map (
            O => \N__62904\,
            I => \N__62487\
        );

    \I__15351\ : SRMux
    port map (
            O => \N__62903\,
            I => \N__62487\
        );

    \I__15350\ : SRMux
    port map (
            O => \N__62902\,
            I => \N__62487\
        );

    \I__15349\ : SRMux
    port map (
            O => \N__62901\,
            I => \N__62487\
        );

    \I__15348\ : SRMux
    port map (
            O => \N__62900\,
            I => \N__62487\
        );

    \I__15347\ : SRMux
    port map (
            O => \N__62899\,
            I => \N__62487\
        );

    \I__15346\ : SRMux
    port map (
            O => \N__62898\,
            I => \N__62487\
        );

    \I__15345\ : SRMux
    port map (
            O => \N__62897\,
            I => \N__62487\
        );

    \I__15344\ : SRMux
    port map (
            O => \N__62896\,
            I => \N__62487\
        );

    \I__15343\ : SRMux
    port map (
            O => \N__62895\,
            I => \N__62487\
        );

    \I__15342\ : SRMux
    port map (
            O => \N__62894\,
            I => \N__62487\
        );

    \I__15341\ : SRMux
    port map (
            O => \N__62893\,
            I => \N__62487\
        );

    \I__15340\ : SRMux
    port map (
            O => \N__62892\,
            I => \N__62487\
        );

    \I__15339\ : SRMux
    port map (
            O => \N__62891\,
            I => \N__62487\
        );

    \I__15338\ : SRMux
    port map (
            O => \N__62890\,
            I => \N__62487\
        );

    \I__15337\ : SRMux
    port map (
            O => \N__62889\,
            I => \N__62487\
        );

    \I__15336\ : SRMux
    port map (
            O => \N__62888\,
            I => \N__62487\
        );

    \I__15335\ : SRMux
    port map (
            O => \N__62887\,
            I => \N__62487\
        );

    \I__15334\ : SRMux
    port map (
            O => \N__62886\,
            I => \N__62487\
        );

    \I__15333\ : SRMux
    port map (
            O => \N__62885\,
            I => \N__62487\
        );

    \I__15332\ : SRMux
    port map (
            O => \N__62884\,
            I => \N__62487\
        );

    \I__15331\ : SRMux
    port map (
            O => \N__62883\,
            I => \N__62487\
        );

    \I__15330\ : SRMux
    port map (
            O => \N__62882\,
            I => \N__62487\
        );

    \I__15329\ : SRMux
    port map (
            O => \N__62881\,
            I => \N__62487\
        );

    \I__15328\ : SRMux
    port map (
            O => \N__62880\,
            I => \N__62487\
        );

    \I__15327\ : SRMux
    port map (
            O => \N__62879\,
            I => \N__62487\
        );

    \I__15326\ : SRMux
    port map (
            O => \N__62878\,
            I => \N__62487\
        );

    \I__15325\ : SRMux
    port map (
            O => \N__62877\,
            I => \N__62487\
        );

    \I__15324\ : SRMux
    port map (
            O => \N__62876\,
            I => \N__62487\
        );

    \I__15323\ : SRMux
    port map (
            O => \N__62875\,
            I => \N__62487\
        );

    \I__15322\ : SRMux
    port map (
            O => \N__62874\,
            I => \N__62487\
        );

    \I__15321\ : SRMux
    port map (
            O => \N__62873\,
            I => \N__62487\
        );

    \I__15320\ : SRMux
    port map (
            O => \N__62872\,
            I => \N__62487\
        );

    \I__15319\ : SRMux
    port map (
            O => \N__62871\,
            I => \N__62487\
        );

    \I__15318\ : SRMux
    port map (
            O => \N__62870\,
            I => \N__62487\
        );

    \I__15317\ : SRMux
    port map (
            O => \N__62869\,
            I => \N__62487\
        );

    \I__15316\ : SRMux
    port map (
            O => \N__62868\,
            I => \N__62487\
        );

    \I__15315\ : SRMux
    port map (
            O => \N__62867\,
            I => \N__62487\
        );

    \I__15314\ : SRMux
    port map (
            O => \N__62866\,
            I => \N__62487\
        );

    \I__15313\ : SRMux
    port map (
            O => \N__62865\,
            I => \N__62487\
        );

    \I__15312\ : SRMux
    port map (
            O => \N__62864\,
            I => \N__62487\
        );

    \I__15311\ : SRMux
    port map (
            O => \N__62863\,
            I => \N__62487\
        );

    \I__15310\ : SRMux
    port map (
            O => \N__62862\,
            I => \N__62487\
        );

    \I__15309\ : SRMux
    port map (
            O => \N__62861\,
            I => \N__62487\
        );

    \I__15308\ : SRMux
    port map (
            O => \N__62860\,
            I => \N__62487\
        );

    \I__15307\ : SRMux
    port map (
            O => \N__62859\,
            I => \N__62487\
        );

    \I__15306\ : SRMux
    port map (
            O => \N__62858\,
            I => \N__62487\
        );

    \I__15305\ : SRMux
    port map (
            O => \N__62857\,
            I => \N__62487\
        );

    \I__15304\ : SRMux
    port map (
            O => \N__62856\,
            I => \N__62487\
        );

    \I__15303\ : SRMux
    port map (
            O => \N__62855\,
            I => \N__62487\
        );

    \I__15302\ : SRMux
    port map (
            O => \N__62854\,
            I => \N__62487\
        );

    \I__15301\ : SRMux
    port map (
            O => \N__62853\,
            I => \N__62487\
        );

    \I__15300\ : SRMux
    port map (
            O => \N__62852\,
            I => \N__62487\
        );

    \I__15299\ : SRMux
    port map (
            O => \N__62851\,
            I => \N__62487\
        );

    \I__15298\ : SRMux
    port map (
            O => \N__62850\,
            I => \N__62487\
        );

    \I__15297\ : SRMux
    port map (
            O => \N__62849\,
            I => \N__62487\
        );

    \I__15296\ : SRMux
    port map (
            O => \N__62848\,
            I => \N__62487\
        );

    \I__15295\ : SRMux
    port map (
            O => \N__62847\,
            I => \N__62487\
        );

    \I__15294\ : SRMux
    port map (
            O => \N__62846\,
            I => \N__62487\
        );

    \I__15293\ : SRMux
    port map (
            O => \N__62845\,
            I => \N__62487\
        );

    \I__15292\ : SRMux
    port map (
            O => \N__62844\,
            I => \N__62487\
        );

    \I__15291\ : SRMux
    port map (
            O => \N__62843\,
            I => \N__62487\
        );

    \I__15290\ : SRMux
    port map (
            O => \N__62842\,
            I => \N__62487\
        );

    \I__15289\ : SRMux
    port map (
            O => \N__62841\,
            I => \N__62487\
        );

    \I__15288\ : SRMux
    port map (
            O => \N__62840\,
            I => \N__62487\
        );

    \I__15287\ : SRMux
    port map (
            O => \N__62839\,
            I => \N__62487\
        );

    \I__15286\ : SRMux
    port map (
            O => \N__62838\,
            I => \N__62487\
        );

    \I__15285\ : SRMux
    port map (
            O => \N__62837\,
            I => \N__62487\
        );

    \I__15284\ : SRMux
    port map (
            O => \N__62836\,
            I => \N__62487\
        );

    \I__15283\ : SRMux
    port map (
            O => \N__62835\,
            I => \N__62487\
        );

    \I__15282\ : SRMux
    port map (
            O => \N__62834\,
            I => \N__62487\
        );

    \I__15281\ : SRMux
    port map (
            O => \N__62833\,
            I => \N__62487\
        );

    \I__15280\ : SRMux
    port map (
            O => \N__62832\,
            I => \N__62487\
        );

    \I__15279\ : SRMux
    port map (
            O => \N__62831\,
            I => \N__62487\
        );

    \I__15278\ : SRMux
    port map (
            O => \N__62830\,
            I => \N__62487\
        );

    \I__15277\ : SRMux
    port map (
            O => \N__62829\,
            I => \N__62487\
        );

    \I__15276\ : SRMux
    port map (
            O => \N__62828\,
            I => \N__62487\
        );

    \I__15275\ : SRMux
    port map (
            O => \N__62827\,
            I => \N__62487\
        );

    \I__15274\ : SRMux
    port map (
            O => \N__62826\,
            I => \N__62487\
        );

    \I__15273\ : SRMux
    port map (
            O => \N__62825\,
            I => \N__62487\
        );

    \I__15272\ : SRMux
    port map (
            O => \N__62824\,
            I => \N__62487\
        );

    \I__15271\ : SRMux
    port map (
            O => \N__62823\,
            I => \N__62487\
        );

    \I__15270\ : SRMux
    port map (
            O => \N__62822\,
            I => \N__62487\
        );

    \I__15269\ : SRMux
    port map (
            O => \N__62821\,
            I => \N__62487\
        );

    \I__15268\ : SRMux
    port map (
            O => \N__62820\,
            I => \N__62487\
        );

    \I__15267\ : SRMux
    port map (
            O => \N__62819\,
            I => \N__62487\
        );

    \I__15266\ : SRMux
    port map (
            O => \N__62818\,
            I => \N__62487\
        );

    \I__15265\ : SRMux
    port map (
            O => \N__62817\,
            I => \N__62487\
        );

    \I__15264\ : SRMux
    port map (
            O => \N__62816\,
            I => \N__62487\
        );

    \I__15263\ : SRMux
    port map (
            O => \N__62815\,
            I => \N__62487\
        );

    \I__15262\ : SRMux
    port map (
            O => \N__62814\,
            I => \N__62487\
        );

    \I__15261\ : SRMux
    port map (
            O => \N__62813\,
            I => \N__62487\
        );

    \I__15260\ : SRMux
    port map (
            O => \N__62812\,
            I => \N__62487\
        );

    \I__15259\ : SRMux
    port map (
            O => \N__62811\,
            I => \N__62487\
        );

    \I__15258\ : SRMux
    port map (
            O => \N__62810\,
            I => \N__62487\
        );

    \I__15257\ : SRMux
    port map (
            O => \N__62809\,
            I => \N__62487\
        );

    \I__15256\ : SRMux
    port map (
            O => \N__62808\,
            I => \N__62487\
        );

    \I__15255\ : SRMux
    port map (
            O => \N__62807\,
            I => \N__62487\
        );

    \I__15254\ : SRMux
    port map (
            O => \N__62806\,
            I => \N__62487\
        );

    \I__15253\ : SRMux
    port map (
            O => \N__62805\,
            I => \N__62487\
        );

    \I__15252\ : SRMux
    port map (
            O => \N__62804\,
            I => \N__62487\
        );

    \I__15251\ : GlobalMux
    port map (
            O => \N__62487\,
            I => \N__62484\
        );

    \I__15250\ : gio2CtrlBuf
    port map (
            O => \N__62484\,
            I => rst_n_c_i_g
        );

    \I__15249\ : InMux
    port map (
            O => \N__62481\,
            I => \N__62476\
        );

    \I__15248\ : InMux
    port map (
            O => \N__62480\,
            I => \N__62473\
        );

    \I__15247\ : InMux
    port map (
            O => \N__62479\,
            I => \N__62469\
        );

    \I__15246\ : LocalMux
    port map (
            O => \N__62476\,
            I => \N__62466\
        );

    \I__15245\ : LocalMux
    port map (
            O => \N__62473\,
            I => \N__62463\
        );

    \I__15244\ : InMux
    port map (
            O => \N__62472\,
            I => \N__62460\
        );

    \I__15243\ : LocalMux
    port map (
            O => \N__62469\,
            I => \N__62457\
        );

    \I__15242\ : Span4Mux_v
    port map (
            O => \N__62466\,
            I => \N__62452\
        );

    \I__15241\ : Span4Mux_v
    port map (
            O => \N__62463\,
            I => \N__62447\
        );

    \I__15240\ : LocalMux
    port map (
            O => \N__62460\,
            I => \N__62447\
        );

    \I__15239\ : Span4Mux_h
    port map (
            O => \N__62457\,
            I => \N__62444\
        );

    \I__15238\ : InMux
    port map (
            O => \N__62456\,
            I => \N__62441\
        );

    \I__15237\ : InMux
    port map (
            O => \N__62455\,
            I => \N__62438\
        );

    \I__15236\ : Span4Mux_h
    port map (
            O => \N__62452\,
            I => \N__62433\
        );

    \I__15235\ : Span4Mux_h
    port map (
            O => \N__62447\,
            I => \N__62433\
        );

    \I__15234\ : Span4Mux_v
    port map (
            O => \N__62444\,
            I => \N__62428\
        );

    \I__15233\ : LocalMux
    port map (
            O => \N__62441\,
            I => \N__62428\
        );

    \I__15232\ : LocalMux
    port map (
            O => \N__62438\,
            I => \c_state_RNIEVJ7_22\
        );

    \I__15231\ : Odrv4
    port map (
            O => \N__62433\,
            I => \c_state_RNIEVJ7_22\
        );

    \I__15230\ : Odrv4
    port map (
            O => \N__62428\,
            I => \c_state_RNIEVJ7_22\
        );

    \I__15229\ : InMux
    port map (
            O => \N__62421\,
            I => \N__62417\
        );

    \I__15228\ : InMux
    port map (
            O => \N__62420\,
            I => \N__62414\
        );

    \I__15227\ : LocalMux
    port map (
            O => \N__62417\,
            I => \N__62411\
        );

    \I__15226\ : LocalMux
    port map (
            O => \N__62414\,
            I => \I2C_top_level_inst1.s_load_rdata2\
        );

    \I__15225\ : Odrv4
    port map (
            O => \N__62411\,
            I => \I2C_top_level_inst1.s_load_rdata2\
        );

    \I__15224\ : InMux
    port map (
            O => \N__62406\,
            I => \N__62403\
        );

    \I__15223\ : LocalMux
    port map (
            O => \N__62403\,
            I => \N__62399\
        );

    \I__15222\ : InMux
    port map (
            O => \N__62402\,
            I => \N__62396\
        );

    \I__15221\ : Span4Mux_v
    port map (
            O => \N__62399\,
            I => \N__62393\
        );

    \I__15220\ : LocalMux
    port map (
            O => \N__62396\,
            I => \N__62390\
        );

    \I__15219\ : Span4Mux_h
    port map (
            O => \N__62393\,
            I => \N__62387\
        );

    \I__15218\ : Odrv4
    port map (
            O => \N__62390\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0\
        );

    \I__15217\ : Odrv4
    port map (
            O => \N__62387\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0\
        );

    \I__15216\ : InMux
    port map (
            O => \N__62382\,
            I => \N__62379\
        );

    \I__15215\ : LocalMux
    port map (
            O => \N__62379\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_27\
        );

    \I__15214\ : CascadeMux
    port map (
            O => \N__62376\,
            I => \N__62373\
        );

    \I__15213\ : InMux
    port map (
            O => \N__62373\,
            I => \N__62370\
        );

    \I__15212\ : LocalMux
    port map (
            O => \N__62370\,
            I => \N__62364\
        );

    \I__15211\ : InMux
    port map (
            O => \N__62369\,
            I => \N__62361\
        );

    \I__15210\ : InMux
    port map (
            O => \N__62368\,
            I => \N__62358\
        );

    \I__15209\ : InMux
    port map (
            O => \N__62367\,
            I => \N__62353\
        );

    \I__15208\ : Span4Mux_v
    port map (
            O => \N__62364\,
            I => \N__62350\
        );

    \I__15207\ : LocalMux
    port map (
            O => \N__62361\,
            I => \N__62347\
        );

    \I__15206\ : LocalMux
    port map (
            O => \N__62358\,
            I => \N__62344\
        );

    \I__15205\ : InMux
    port map (
            O => \N__62357\,
            I => \N__62341\
        );

    \I__15204\ : InMux
    port map (
            O => \N__62356\,
            I => \N__62338\
        );

    \I__15203\ : LocalMux
    port map (
            O => \N__62353\,
            I => \N__62333\
        );

    \I__15202\ : Span4Mux_v
    port map (
            O => \N__62350\,
            I => \N__62330\
        );

    \I__15201\ : Span4Mux_h
    port map (
            O => \N__62347\,
            I => \N__62327\
        );

    \I__15200\ : Span4Mux_v
    port map (
            O => \N__62344\,
            I => \N__62320\
        );

    \I__15199\ : LocalMux
    port map (
            O => \N__62341\,
            I => \N__62320\
        );

    \I__15198\ : LocalMux
    port map (
            O => \N__62338\,
            I => \N__62320\
        );

    \I__15197\ : InMux
    port map (
            O => \N__62337\,
            I => \N__62317\
        );

    \I__15196\ : InMux
    port map (
            O => \N__62336\,
            I => \N__62314\
        );

    \I__15195\ : Span4Mux_v
    port map (
            O => \N__62333\,
            I => \N__62311\
        );

    \I__15194\ : Span4Mux_h
    port map (
            O => \N__62330\,
            I => \N__62306\
        );

    \I__15193\ : Span4Mux_v
    port map (
            O => \N__62327\,
            I => \N__62306\
        );

    \I__15192\ : Span4Mux_h
    port map (
            O => \N__62320\,
            I => \N__62303\
        );

    \I__15191\ : LocalMux
    port map (
            O => \N__62317\,
            I => \N__62300\
        );

    \I__15190\ : LocalMux
    port map (
            O => \N__62314\,
            I => \N__62295\
        );

    \I__15189\ : Sp12to4
    port map (
            O => \N__62311\,
            I => \N__62295\
        );

    \I__15188\ : Span4Mux_h
    port map (
            O => \N__62306\,
            I => \N__62292\
        );

    \I__15187\ : Span4Mux_v
    port map (
            O => \N__62303\,
            I => \N__62289\
        );

    \I__15186\ : Span4Mux_v
    port map (
            O => \N__62300\,
            I => \N__62286\
        );

    \I__15185\ : Span12Mux_h
    port map (
            O => \N__62295\,
            I => \N__62281\
        );

    \I__15184\ : Sp12to4
    port map (
            O => \N__62292\,
            I => \N__62281\
        );

    \I__15183\ : Span4Mux_h
    port map (
            O => \N__62289\,
            I => \N__62276\
        );

    \I__15182\ : Span4Mux_h
    port map (
            O => \N__62286\,
            I => \N__62276\
        );

    \I__15181\ : Odrv12
    port map (
            O => \N__62281\,
            I => \I2C_top_level_inst1_s_data_oreg_28\
        );

    \I__15180\ : Odrv4
    port map (
            O => \N__62276\,
            I => \I2C_top_level_inst1_s_data_oreg_28\
        );

    \I__15179\ : InMux
    port map (
            O => \N__62271\,
            I => \N__62268\
        );

    \I__15178\ : LocalMux
    port map (
            O => \N__62268\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_28\
        );

    \I__15177\ : InMux
    port map (
            O => \N__62265\,
            I => \N__62256\
        );

    \I__15176\ : InMux
    port map (
            O => \N__62264\,
            I => \N__62253\
        );

    \I__15175\ : InMux
    port map (
            O => \N__62263\,
            I => \N__62250\
        );

    \I__15174\ : InMux
    port map (
            O => \N__62262\,
            I => \N__62247\
        );

    \I__15173\ : InMux
    port map (
            O => \N__62261\,
            I => \N__62243\
        );

    \I__15172\ : InMux
    port map (
            O => \N__62260\,
            I => \N__62240\
        );

    \I__15171\ : InMux
    port map (
            O => \N__62259\,
            I => \N__62237\
        );

    \I__15170\ : LocalMux
    port map (
            O => \N__62256\,
            I => \N__62234\
        );

    \I__15169\ : LocalMux
    port map (
            O => \N__62253\,
            I => \N__62231\
        );

    \I__15168\ : LocalMux
    port map (
            O => \N__62250\,
            I => \N__62226\
        );

    \I__15167\ : LocalMux
    port map (
            O => \N__62247\,
            I => \N__62226\
        );

    \I__15166\ : InMux
    port map (
            O => \N__62246\,
            I => \N__62223\
        );

    \I__15165\ : LocalMux
    port map (
            O => \N__62243\,
            I => \N__62218\
        );

    \I__15164\ : LocalMux
    port map (
            O => \N__62240\,
            I => \N__62218\
        );

    \I__15163\ : LocalMux
    port map (
            O => \N__62237\,
            I => \N__62215\
        );

    \I__15162\ : Sp12to4
    port map (
            O => \N__62234\,
            I => \N__62212\
        );

    \I__15161\ : Span4Mux_v
    port map (
            O => \N__62231\,
            I => \N__62209\
        );

    \I__15160\ : Span4Mux_v
    port map (
            O => \N__62226\,
            I => \N__62206\
        );

    \I__15159\ : LocalMux
    port map (
            O => \N__62223\,
            I => \N__62197\
        );

    \I__15158\ : Span12Mux_v
    port map (
            O => \N__62218\,
            I => \N__62197\
        );

    \I__15157\ : Span12Mux_v
    port map (
            O => \N__62215\,
            I => \N__62197\
        );

    \I__15156\ : Span12Mux_s11_h
    port map (
            O => \N__62212\,
            I => \N__62197\
        );

    \I__15155\ : Odrv4
    port map (
            O => \N__62209\,
            I => \I2C_top_level_inst1_s_data_oreg_29\
        );

    \I__15154\ : Odrv4
    port map (
            O => \N__62206\,
            I => \I2C_top_level_inst1_s_data_oreg_29\
        );

    \I__15153\ : Odrv12
    port map (
            O => \N__62197\,
            I => \I2C_top_level_inst1_s_data_oreg_29\
        );

    \I__15152\ : InMux
    port map (
            O => \N__62190\,
            I => \N__62187\
        );

    \I__15151\ : LocalMux
    port map (
            O => \N__62187\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_29\
        );

    \I__15150\ : InMux
    port map (
            O => \N__62184\,
            I => \N__62180\
        );

    \I__15149\ : CascadeMux
    port map (
            O => \N__62183\,
            I => \N__62176\
        );

    \I__15148\ : LocalMux
    port map (
            O => \N__62180\,
            I => \N__62173\
        );

    \I__15147\ : InMux
    port map (
            O => \N__62179\,
            I => \N__62170\
        );

    \I__15146\ : InMux
    port map (
            O => \N__62176\,
            I => \N__62166\
        );

    \I__15145\ : Span4Mux_v
    port map (
            O => \N__62173\,
            I => \N__62160\
        );

    \I__15144\ : LocalMux
    port map (
            O => \N__62170\,
            I => \N__62160\
        );

    \I__15143\ : InMux
    port map (
            O => \N__62169\,
            I => \N__62157\
        );

    \I__15142\ : LocalMux
    port map (
            O => \N__62166\,
            I => \N__62154\
        );

    \I__15141\ : InMux
    port map (
            O => \N__62165\,
            I => \N__62151\
        );

    \I__15140\ : Span4Mux_h
    port map (
            O => \N__62160\,
            I => \N__62148\
        );

    \I__15139\ : LocalMux
    port map (
            O => \N__62157\,
            I => \N__62144\
        );

    \I__15138\ : Span4Mux_h
    port map (
            O => \N__62154\,
            I => \N__62139\
        );

    \I__15137\ : LocalMux
    port map (
            O => \N__62151\,
            I => \N__62139\
        );

    \I__15136\ : Span4Mux_v
    port map (
            O => \N__62148\,
            I => \N__62136\
        );

    \I__15135\ : InMux
    port map (
            O => \N__62147\,
            I => \N__62133\
        );

    \I__15134\ : Span4Mux_v
    port map (
            O => \N__62144\,
            I => \N__62129\
        );

    \I__15133\ : Span4Mux_v
    port map (
            O => \N__62139\,
            I => \N__62126\
        );

    \I__15132\ : Span4Mux_h
    port map (
            O => \N__62136\,
            I => \N__62120\
        );

    \I__15131\ : LocalMux
    port map (
            O => \N__62133\,
            I => \N__62120\
        );

    \I__15130\ : InMux
    port map (
            O => \N__62132\,
            I => \N__62117\
        );

    \I__15129\ : Span4Mux_v
    port map (
            O => \N__62129\,
            I => \N__62114\
        );

    \I__15128\ : Span4Mux_v
    port map (
            O => \N__62126\,
            I => \N__62111\
        );

    \I__15127\ : InMux
    port map (
            O => \N__62125\,
            I => \N__62108\
        );

    \I__15126\ : Span4Mux_h
    port map (
            O => \N__62120\,
            I => \N__62105\
        );

    \I__15125\ : LocalMux
    port map (
            O => \N__62117\,
            I => \N__62102\
        );

    \I__15124\ : Sp12to4
    port map (
            O => \N__62114\,
            I => \N__62097\
        );

    \I__15123\ : Sp12to4
    port map (
            O => \N__62111\,
            I => \N__62097\
        );

    \I__15122\ : LocalMux
    port map (
            O => \N__62108\,
            I => \N__62090\
        );

    \I__15121\ : Span4Mux_v
    port map (
            O => \N__62105\,
            I => \N__62090\
        );

    \I__15120\ : Span4Mux_v
    port map (
            O => \N__62102\,
            I => \N__62090\
        );

    \I__15119\ : Span12Mux_h
    port map (
            O => \N__62097\,
            I => \N__62087\
        );

    \I__15118\ : Span4Mux_h
    port map (
            O => \N__62090\,
            I => \N__62084\
        );

    \I__15117\ : Odrv12
    port map (
            O => \N__62087\,
            I => \I2C_top_level_inst1_s_data_oreg_30\
        );

    \I__15116\ : Odrv4
    port map (
            O => \N__62084\,
            I => \I2C_top_level_inst1_s_data_oreg_30\
        );

    \I__15115\ : InMux
    port map (
            O => \N__62079\,
            I => \N__62076\
        );

    \I__15114\ : LocalMux
    port map (
            O => \N__62076\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_30\
        );

    \I__15113\ : InMux
    port map (
            O => \N__62073\,
            I => \N__62067\
        );

    \I__15112\ : InMux
    port map (
            O => \N__62072\,
            I => \N__62064\
        );

    \I__15111\ : InMux
    port map (
            O => \N__62071\,
            I => \N__62061\
        );

    \I__15110\ : InMux
    port map (
            O => \N__62070\,
            I => \N__62056\
        );

    \I__15109\ : LocalMux
    port map (
            O => \N__62067\,
            I => \N__62051\
        );

    \I__15108\ : LocalMux
    port map (
            O => \N__62064\,
            I => \N__62051\
        );

    \I__15107\ : LocalMux
    port map (
            O => \N__62061\,
            I => \N__62048\
        );

    \I__15106\ : CascadeMux
    port map (
            O => \N__62060\,
            I => \N__62045\
        );

    \I__15105\ : InMux
    port map (
            O => \N__62059\,
            I => \N__62041\
        );

    \I__15104\ : LocalMux
    port map (
            O => \N__62056\,
            I => \N__62038\
        );

    \I__15103\ : Span4Mux_v
    port map (
            O => \N__62051\,
            I => \N__62033\
        );

    \I__15102\ : Span4Mux_h
    port map (
            O => \N__62048\,
            I => \N__62033\
        );

    \I__15101\ : InMux
    port map (
            O => \N__62045\,
            I => \N__62028\
        );

    \I__15100\ : InMux
    port map (
            O => \N__62044\,
            I => \N__62028\
        );

    \I__15099\ : LocalMux
    port map (
            O => \N__62041\,
            I => \N__62025\
        );

    \I__15098\ : Span4Mux_v
    port map (
            O => \N__62038\,
            I => \N__62019\
        );

    \I__15097\ : Span4Mux_h
    port map (
            O => \N__62033\,
            I => \N__62019\
        );

    \I__15096\ : LocalMux
    port map (
            O => \N__62028\,
            I => \N__62016\
        );

    \I__15095\ : Span12Mux_v
    port map (
            O => \N__62025\,
            I => \N__62013\
        );

    \I__15094\ : InMux
    port map (
            O => \N__62024\,
            I => \N__62010\
        );

    \I__15093\ : Span4Mux_h
    port map (
            O => \N__62019\,
            I => \N__62007\
        );

    \I__15092\ : Span4Mux_h
    port map (
            O => \N__62016\,
            I => \N__62004\
        );

    \I__15091\ : Span12Mux_h
    port map (
            O => \N__62013\,
            I => \N__62001\
        );

    \I__15090\ : LocalMux
    port map (
            O => \N__62010\,
            I => \N__61994\
        );

    \I__15089\ : Span4Mux_v
    port map (
            O => \N__62007\,
            I => \N__61994\
        );

    \I__15088\ : Span4Mux_v
    port map (
            O => \N__62004\,
            I => \N__61994\
        );

    \I__15087\ : Odrv12
    port map (
            O => \N__62001\,
            I => \I2C_top_level_inst1_s_data_oreg_31\
        );

    \I__15086\ : Odrv4
    port map (
            O => \N__61994\,
            I => \I2C_top_level_inst1_s_data_oreg_31\
        );

    \I__15085\ : InMux
    port map (
            O => \N__61989\,
            I => \N__61986\
        );

    \I__15084\ : LocalMux
    port map (
            O => \N__61986\,
            I => \N__61983\
        );

    \I__15083\ : Span4Mux_v
    port map (
            O => \N__61983\,
            I => \N__61980\
        );

    \I__15082\ : Span4Mux_h
    port map (
            O => \N__61980\,
            I => \N__61977\
        );

    \I__15081\ : Span4Mux_h
    port map (
            O => \N__61977\,
            I => \N__61974\
        );

    \I__15080\ : Odrv4
    port map (
            O => \N__61974\,
            I => \I2C_top_level_inst1.s_sda_o_reg\
        );

    \I__15079\ : InMux
    port map (
            O => \N__61971\,
            I => \N__61965\
        );

    \I__15078\ : InMux
    port map (
            O => \N__61970\,
            I => \N__61960\
        );

    \I__15077\ : InMux
    port map (
            O => \N__61969\,
            I => \N__61956\
        );

    \I__15076\ : InMux
    port map (
            O => \N__61968\,
            I => \N__61953\
        );

    \I__15075\ : LocalMux
    port map (
            O => \N__61965\,
            I => \N__61950\
        );

    \I__15074\ : InMux
    port map (
            O => \N__61964\,
            I => \N__61947\
        );

    \I__15073\ : InMux
    port map (
            O => \N__61963\,
            I => \N__61944\
        );

    \I__15072\ : LocalMux
    port map (
            O => \N__61960\,
            I => \N__61940\
        );

    \I__15071\ : InMux
    port map (
            O => \N__61959\,
            I => \N__61937\
        );

    \I__15070\ : LocalMux
    port map (
            O => \N__61956\,
            I => \N__61934\
        );

    \I__15069\ : LocalMux
    port map (
            O => \N__61953\,
            I => \N__61931\
        );

    \I__15068\ : Span4Mux_v
    port map (
            O => \N__61950\,
            I => \N__61927\
        );

    \I__15067\ : LocalMux
    port map (
            O => \N__61947\,
            I => \N__61922\
        );

    \I__15066\ : LocalMux
    port map (
            O => \N__61944\,
            I => \N__61922\
        );

    \I__15065\ : InMux
    port map (
            O => \N__61943\,
            I => \N__61919\
        );

    \I__15064\ : Span4Mux_v
    port map (
            O => \N__61940\,
            I => \N__61910\
        );

    \I__15063\ : LocalMux
    port map (
            O => \N__61937\,
            I => \N__61910\
        );

    \I__15062\ : Span4Mux_h
    port map (
            O => \N__61934\,
            I => \N__61910\
        );

    \I__15061\ : Span4Mux_v
    port map (
            O => \N__61931\,
            I => \N__61910\
        );

    \I__15060\ : InMux
    port map (
            O => \N__61930\,
            I => \N__61907\
        );

    \I__15059\ : Sp12to4
    port map (
            O => \N__61927\,
            I => \N__61904\
        );

    \I__15058\ : Span12Mux_s9_v
    port map (
            O => \N__61922\,
            I => \N__61901\
        );

    \I__15057\ : LocalMux
    port map (
            O => \N__61919\,
            I => \N__61898\
        );

    \I__15056\ : Span4Mux_v
    port map (
            O => \N__61910\,
            I => \N__61895\
        );

    \I__15055\ : LocalMux
    port map (
            O => \N__61907\,
            I => \N__61890\
        );

    \I__15054\ : Span12Mux_h
    port map (
            O => \N__61904\,
            I => \N__61890\
        );

    \I__15053\ : Span12Mux_h
    port map (
            O => \N__61901\,
            I => \N__61887\
        );

    \I__15052\ : Odrv4
    port map (
            O => \N__61898\,
            I => \I2C_top_level_inst1_s_data_oreg_0\
        );

    \I__15051\ : Odrv4
    port map (
            O => \N__61895\,
            I => \I2C_top_level_inst1_s_data_oreg_0\
        );

    \I__15050\ : Odrv12
    port map (
            O => \N__61890\,
            I => \I2C_top_level_inst1_s_data_oreg_0\
        );

    \I__15049\ : Odrv12
    port map (
            O => \N__61887\,
            I => \I2C_top_level_inst1_s_data_oreg_0\
        );

    \I__15048\ : InMux
    port map (
            O => \N__61878\,
            I => \N__61875\
        );

    \I__15047\ : LocalMux
    port map (
            O => \N__61875\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_0\
        );

    \I__15046\ : InMux
    port map (
            O => \N__61872\,
            I => \N__61868\
        );

    \I__15045\ : InMux
    port map (
            O => \N__61871\,
            I => \N__61864\
        );

    \I__15044\ : LocalMux
    port map (
            O => \N__61868\,
            I => \N__61856\
        );

    \I__15043\ : InMux
    port map (
            O => \N__61867\,
            I => \N__61853\
        );

    \I__15042\ : LocalMux
    port map (
            O => \N__61864\,
            I => \N__61850\
        );

    \I__15041\ : InMux
    port map (
            O => \N__61863\,
            I => \N__61847\
        );

    \I__15040\ : CascadeMux
    port map (
            O => \N__61862\,
            I => \N__61844\
        );

    \I__15039\ : InMux
    port map (
            O => \N__61861\,
            I => \N__61841\
        );

    \I__15038\ : InMux
    port map (
            O => \N__61860\,
            I => \N__61838\
        );

    \I__15037\ : InMux
    port map (
            O => \N__61859\,
            I => \N__61835\
        );

    \I__15036\ : Span4Mux_v
    port map (
            O => \N__61856\,
            I => \N__61832\
        );

    \I__15035\ : LocalMux
    port map (
            O => \N__61853\,
            I => \N__61827\
        );

    \I__15034\ : Span4Mux_v
    port map (
            O => \N__61850\,
            I => \N__61827\
        );

    \I__15033\ : LocalMux
    port map (
            O => \N__61847\,
            I => \N__61824\
        );

    \I__15032\ : InMux
    port map (
            O => \N__61844\,
            I => \N__61821\
        );

    \I__15031\ : LocalMux
    port map (
            O => \N__61841\,
            I => \N__61817\
        );

    \I__15030\ : LocalMux
    port map (
            O => \N__61838\,
            I => \N__61814\
        );

    \I__15029\ : LocalMux
    port map (
            O => \N__61835\,
            I => \N__61811\
        );

    \I__15028\ : Span4Mux_v
    port map (
            O => \N__61832\,
            I => \N__61808\
        );

    \I__15027\ : Span4Mux_h
    port map (
            O => \N__61827\,
            I => \N__61803\
        );

    \I__15026\ : Span4Mux_v
    port map (
            O => \N__61824\,
            I => \N__61803\
        );

    \I__15025\ : LocalMux
    port map (
            O => \N__61821\,
            I => \N__61800\
        );

    \I__15024\ : InMux
    port map (
            O => \N__61820\,
            I => \N__61797\
        );

    \I__15023\ : Span4Mux_v
    port map (
            O => \N__61817\,
            I => \N__61794\
        );

    \I__15022\ : Span4Mux_v
    port map (
            O => \N__61814\,
            I => \N__61791\
        );

    \I__15021\ : Span4Mux_v
    port map (
            O => \N__61811\,
            I => \N__61788\
        );

    \I__15020\ : Sp12to4
    port map (
            O => \N__61808\,
            I => \N__61785\
        );

    \I__15019\ : Span4Mux_h
    port map (
            O => \N__61803\,
            I => \N__61782\
        );

    \I__15018\ : Span4Mux_h
    port map (
            O => \N__61800\,
            I => \N__61779\
        );

    \I__15017\ : LocalMux
    port map (
            O => \N__61797\,
            I => \N__61776\
        );

    \I__15016\ : Span4Mux_h
    port map (
            O => \N__61794\,
            I => \N__61773\
        );

    \I__15015\ : Sp12to4
    port map (
            O => \N__61791\,
            I => \N__61766\
        );

    \I__15014\ : Sp12to4
    port map (
            O => \N__61788\,
            I => \N__61766\
        );

    \I__15013\ : Span12Mux_s10_h
    port map (
            O => \N__61785\,
            I => \N__61766\
        );

    \I__15012\ : Span4Mux_v
    port map (
            O => \N__61782\,
            I => \N__61759\
        );

    \I__15011\ : Span4Mux_v
    port map (
            O => \N__61779\,
            I => \N__61759\
        );

    \I__15010\ : Span4Mux_h
    port map (
            O => \N__61776\,
            I => \N__61759\
        );

    \I__15009\ : Odrv4
    port map (
            O => \N__61773\,
            I => \I2C_top_level_inst1_s_data_oreg_1\
        );

    \I__15008\ : Odrv12
    port map (
            O => \N__61766\,
            I => \I2C_top_level_inst1_s_data_oreg_1\
        );

    \I__15007\ : Odrv4
    port map (
            O => \N__61759\,
            I => \I2C_top_level_inst1_s_data_oreg_1\
        );

    \I__15006\ : InMux
    port map (
            O => \N__61752\,
            I => \N__61749\
        );

    \I__15005\ : LocalMux
    port map (
            O => \N__61749\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_1\
        );

    \I__15004\ : InMux
    port map (
            O => \N__61746\,
            I => \N__61742\
        );

    \I__15003\ : InMux
    port map (
            O => \N__61745\,
            I => \N__61739\
        );

    \I__15002\ : LocalMux
    port map (
            O => \N__61742\,
            I => \N__61734\
        );

    \I__15001\ : LocalMux
    port map (
            O => \N__61739\,
            I => \N__61731\
        );

    \I__15000\ : InMux
    port map (
            O => \N__61738\,
            I => \N__61726\
        );

    \I__14999\ : InMux
    port map (
            O => \N__61737\,
            I => \N__61723\
        );

    \I__14998\ : Span4Mux_v
    port map (
            O => \N__61734\,
            I => \N__61720\
        );

    \I__14997\ : Span4Mux_h
    port map (
            O => \N__61731\,
            I => \N__61716\
        );

    \I__14996\ : InMux
    port map (
            O => \N__61730\,
            I => \N__61713\
        );

    \I__14995\ : InMux
    port map (
            O => \N__61729\,
            I => \N__61708\
        );

    \I__14994\ : LocalMux
    port map (
            O => \N__61726\,
            I => \N__61705\
        );

    \I__14993\ : LocalMux
    port map (
            O => \N__61723\,
            I => \N__61700\
        );

    \I__14992\ : Span4Mux_h
    port map (
            O => \N__61720\,
            I => \N__61700\
        );

    \I__14991\ : InMux
    port map (
            O => \N__61719\,
            I => \N__61697\
        );

    \I__14990\ : Span4Mux_v
    port map (
            O => \N__61716\,
            I => \N__61694\
        );

    \I__14989\ : LocalMux
    port map (
            O => \N__61713\,
            I => \N__61691\
        );

    \I__14988\ : CascadeMux
    port map (
            O => \N__61712\,
            I => \N__61688\
        );

    \I__14987\ : InMux
    port map (
            O => \N__61711\,
            I => \N__61685\
        );

    \I__14986\ : LocalMux
    port map (
            O => \N__61708\,
            I => \N__61682\
        );

    \I__14985\ : Sp12to4
    port map (
            O => \N__61705\,
            I => \N__61675\
        );

    \I__14984\ : Sp12to4
    port map (
            O => \N__61700\,
            I => \N__61675\
        );

    \I__14983\ : LocalMux
    port map (
            O => \N__61697\,
            I => \N__61675\
        );

    \I__14982\ : Span4Mux_h
    port map (
            O => \N__61694\,
            I => \N__61670\
        );

    \I__14981\ : Span4Mux_h
    port map (
            O => \N__61691\,
            I => \N__61670\
        );

    \I__14980\ : InMux
    port map (
            O => \N__61688\,
            I => \N__61667\
        );

    \I__14979\ : LocalMux
    port map (
            O => \N__61685\,
            I => \N__61662\
        );

    \I__14978\ : Sp12to4
    port map (
            O => \N__61682\,
            I => \N__61662\
        );

    \I__14977\ : Span12Mux_v
    port map (
            O => \N__61675\,
            I => \N__61659\
        );

    \I__14976\ : Span4Mux_h
    port map (
            O => \N__61670\,
            I => \N__61656\
        );

    \I__14975\ : LocalMux
    port map (
            O => \N__61667\,
            I => \I2C_top_level_inst1_s_data_oreg_2\
        );

    \I__14974\ : Odrv12
    port map (
            O => \N__61662\,
            I => \I2C_top_level_inst1_s_data_oreg_2\
        );

    \I__14973\ : Odrv12
    port map (
            O => \N__61659\,
            I => \I2C_top_level_inst1_s_data_oreg_2\
        );

    \I__14972\ : Odrv4
    port map (
            O => \N__61656\,
            I => \I2C_top_level_inst1_s_data_oreg_2\
        );

    \I__14971\ : InMux
    port map (
            O => \N__61647\,
            I => \N__61641\
        );

    \I__14970\ : InMux
    port map (
            O => \N__61646\,
            I => \N__61636\
        );

    \I__14969\ : InMux
    port map (
            O => \N__61645\,
            I => \N__61633\
        );

    \I__14968\ : InMux
    port map (
            O => \N__61644\,
            I => \N__61628\
        );

    \I__14967\ : LocalMux
    port map (
            O => \N__61641\,
            I => \N__61625\
        );

    \I__14966\ : InMux
    port map (
            O => \N__61640\,
            I => \N__61622\
        );

    \I__14965\ : InMux
    port map (
            O => \N__61639\,
            I => \N__61619\
        );

    \I__14964\ : LocalMux
    port map (
            O => \N__61636\,
            I => \N__61614\
        );

    \I__14963\ : LocalMux
    port map (
            O => \N__61633\,
            I => \N__61614\
        );

    \I__14962\ : CascadeMux
    port map (
            O => \N__61632\,
            I => \N__61610\
        );

    \I__14961\ : InMux
    port map (
            O => \N__61631\,
            I => \N__61607\
        );

    \I__14960\ : LocalMux
    port map (
            O => \N__61628\,
            I => \N__61604\
        );

    \I__14959\ : Span4Mux_v
    port map (
            O => \N__61625\,
            I => \N__61599\
        );

    \I__14958\ : LocalMux
    port map (
            O => \N__61622\,
            I => \N__61599\
        );

    \I__14957\ : LocalMux
    port map (
            O => \N__61619\,
            I => \N__61596\
        );

    \I__14956\ : Span4Mux_v
    port map (
            O => \N__61614\,
            I => \N__61593\
        );

    \I__14955\ : InMux
    port map (
            O => \N__61613\,
            I => \N__61590\
        );

    \I__14954\ : InMux
    port map (
            O => \N__61610\,
            I => \N__61587\
        );

    \I__14953\ : LocalMux
    port map (
            O => \N__61607\,
            I => \N__61580\
        );

    \I__14952\ : Span4Mux_v
    port map (
            O => \N__61604\,
            I => \N__61580\
        );

    \I__14951\ : Span4Mux_v
    port map (
            O => \N__61599\,
            I => \N__61580\
        );

    \I__14950\ : Span4Mux_v
    port map (
            O => \N__61596\,
            I => \N__61575\
        );

    \I__14949\ : Span4Mux_h
    port map (
            O => \N__61593\,
            I => \N__61575\
        );

    \I__14948\ : LocalMux
    port map (
            O => \N__61590\,
            I => \N__61572\
        );

    \I__14947\ : LocalMux
    port map (
            O => \N__61587\,
            I => \N__61569\
        );

    \I__14946\ : Span4Mux_h
    port map (
            O => \N__61580\,
            I => \N__61566\
        );

    \I__14945\ : Span4Mux_h
    port map (
            O => \N__61575\,
            I => \N__61559\
        );

    \I__14944\ : Span4Mux_v
    port map (
            O => \N__61572\,
            I => \N__61559\
        );

    \I__14943\ : Span4Mux_v
    port map (
            O => \N__61569\,
            I => \N__61559\
        );

    \I__14942\ : Sp12to4
    port map (
            O => \N__61566\,
            I => \N__61554\
        );

    \I__14941\ : Sp12to4
    port map (
            O => \N__61559\,
            I => \N__61554\
        );

    \I__14940\ : Odrv12
    port map (
            O => \N__61554\,
            I => \I2C_top_level_inst1_s_data_oreg_19\
        );

    \I__14939\ : InMux
    port map (
            O => \N__61551\,
            I => \N__61548\
        );

    \I__14938\ : LocalMux
    port map (
            O => \N__61548\,
            I => \N__61541\
        );

    \I__14937\ : InMux
    port map (
            O => \N__61547\,
            I => \N__61538\
        );

    \I__14936\ : InMux
    port map (
            O => \N__61546\,
            I => \N__61535\
        );

    \I__14935\ : InMux
    port map (
            O => \N__61545\,
            I => \N__61532\
        );

    \I__14934\ : InMux
    port map (
            O => \N__61544\,
            I => \N__61527\
        );

    \I__14933\ : Span4Mux_v
    port map (
            O => \N__61541\,
            I => \N__61522\
        );

    \I__14932\ : LocalMux
    port map (
            O => \N__61538\,
            I => \N__61517\
        );

    \I__14931\ : LocalMux
    port map (
            O => \N__61535\,
            I => \N__61517\
        );

    \I__14930\ : LocalMux
    port map (
            O => \N__61532\,
            I => \N__61514\
        );

    \I__14929\ : InMux
    port map (
            O => \N__61531\,
            I => \N__61511\
        );

    \I__14928\ : InMux
    port map (
            O => \N__61530\,
            I => \N__61508\
        );

    \I__14927\ : LocalMux
    port map (
            O => \N__61527\,
            I => \N__61505\
        );

    \I__14926\ : InMux
    port map (
            O => \N__61526\,
            I => \N__61502\
        );

    \I__14925\ : InMux
    port map (
            O => \N__61525\,
            I => \N__61499\
        );

    \I__14924\ : Span4Mux_h
    port map (
            O => \N__61522\,
            I => \N__61494\
        );

    \I__14923\ : Span4Mux_v
    port map (
            O => \N__61517\,
            I => \N__61494\
        );

    \I__14922\ : Span4Mux_v
    port map (
            O => \N__61514\,
            I => \N__61491\
        );

    \I__14921\ : LocalMux
    port map (
            O => \N__61511\,
            I => \N__61486\
        );

    \I__14920\ : LocalMux
    port map (
            O => \N__61508\,
            I => \N__61486\
        );

    \I__14919\ : Span4Mux_v
    port map (
            O => \N__61505\,
            I => \N__61483\
        );

    \I__14918\ : LocalMux
    port map (
            O => \N__61502\,
            I => \N__61478\
        );

    \I__14917\ : LocalMux
    port map (
            O => \N__61499\,
            I => \N__61478\
        );

    \I__14916\ : Sp12to4
    port map (
            O => \N__61494\,
            I => \N__61473\
        );

    \I__14915\ : Sp12to4
    port map (
            O => \N__61491\,
            I => \N__61473\
        );

    \I__14914\ : Span4Mux_v
    port map (
            O => \N__61486\,
            I => \N__61468\
        );

    \I__14913\ : Span4Mux_h
    port map (
            O => \N__61483\,
            I => \N__61468\
        );

    \I__14912\ : Odrv4
    port map (
            O => \N__61478\,
            I => \I2C_top_level_inst1_s_data_oreg_20\
        );

    \I__14911\ : Odrv12
    port map (
            O => \N__61473\,
            I => \I2C_top_level_inst1_s_data_oreg_20\
        );

    \I__14910\ : Odrv4
    port map (
            O => \N__61468\,
            I => \I2C_top_level_inst1_s_data_oreg_20\
        );

    \I__14909\ : InMux
    port map (
            O => \N__61461\,
            I => \N__61458\
        );

    \I__14908\ : LocalMux
    port map (
            O => \N__61458\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_19\
        );

    \I__14907\ : InMux
    port map (
            O => \N__61455\,
            I => \N__61452\
        );

    \I__14906\ : LocalMux
    port map (
            O => \N__61452\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_20\
        );

    \I__14905\ : InMux
    port map (
            O => \N__61449\,
            I => \N__61444\
        );

    \I__14904\ : CascadeMux
    port map (
            O => \N__61448\,
            I => \N__61441\
        );

    \I__14903\ : InMux
    port map (
            O => \N__61447\,
            I => \N__61438\
        );

    \I__14902\ : LocalMux
    port map (
            O => \N__61444\,
            I => \N__61431\
        );

    \I__14901\ : InMux
    port map (
            O => \N__61441\,
            I => \N__61428\
        );

    \I__14900\ : LocalMux
    port map (
            O => \N__61438\,
            I => \N__61425\
        );

    \I__14899\ : InMux
    port map (
            O => \N__61437\,
            I => \N__61422\
        );

    \I__14898\ : InMux
    port map (
            O => \N__61436\,
            I => \N__61418\
        );

    \I__14897\ : InMux
    port map (
            O => \N__61435\,
            I => \N__61415\
        );

    \I__14896\ : InMux
    port map (
            O => \N__61434\,
            I => \N__61412\
        );

    \I__14895\ : Span4Mux_v
    port map (
            O => \N__61431\,
            I => \N__61407\
        );

    \I__14894\ : LocalMux
    port map (
            O => \N__61428\,
            I => \N__61407\
        );

    \I__14893\ : Span4Mux_h
    port map (
            O => \N__61425\,
            I => \N__61401\
        );

    \I__14892\ : LocalMux
    port map (
            O => \N__61422\,
            I => \N__61401\
        );

    \I__14891\ : InMux
    port map (
            O => \N__61421\,
            I => \N__61398\
        );

    \I__14890\ : LocalMux
    port map (
            O => \N__61418\,
            I => \N__61395\
        );

    \I__14889\ : LocalMux
    port map (
            O => \N__61415\,
            I => \N__61390\
        );

    \I__14888\ : LocalMux
    port map (
            O => \N__61412\,
            I => \N__61390\
        );

    \I__14887\ : Span4Mux_h
    port map (
            O => \N__61407\,
            I => \N__61387\
        );

    \I__14886\ : InMux
    port map (
            O => \N__61406\,
            I => \N__61384\
        );

    \I__14885\ : Span4Mux_h
    port map (
            O => \N__61401\,
            I => \N__61381\
        );

    \I__14884\ : LocalMux
    port map (
            O => \N__61398\,
            I => \N__61376\
        );

    \I__14883\ : Span4Mux_h
    port map (
            O => \N__61395\,
            I => \N__61376\
        );

    \I__14882\ : Span4Mux_v
    port map (
            O => \N__61390\,
            I => \N__61371\
        );

    \I__14881\ : Span4Mux_h
    port map (
            O => \N__61387\,
            I => \N__61371\
        );

    \I__14880\ : LocalMux
    port map (
            O => \N__61384\,
            I => \I2C_top_level_inst1_s_data_oreg_21\
        );

    \I__14879\ : Odrv4
    port map (
            O => \N__61381\,
            I => \I2C_top_level_inst1_s_data_oreg_21\
        );

    \I__14878\ : Odrv4
    port map (
            O => \N__61376\,
            I => \I2C_top_level_inst1_s_data_oreg_21\
        );

    \I__14877\ : Odrv4
    port map (
            O => \N__61371\,
            I => \I2C_top_level_inst1_s_data_oreg_21\
        );

    \I__14876\ : InMux
    port map (
            O => \N__61362\,
            I => \N__61359\
        );

    \I__14875\ : LocalMux
    port map (
            O => \N__61359\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_21\
        );

    \I__14874\ : InMux
    port map (
            O => \N__61356\,
            I => \N__61349\
        );

    \I__14873\ : InMux
    port map (
            O => \N__61355\,
            I => \N__61345\
        );

    \I__14872\ : InMux
    port map (
            O => \N__61354\,
            I => \N__61342\
        );

    \I__14871\ : InMux
    port map (
            O => \N__61353\,
            I => \N__61339\
        );

    \I__14870\ : InMux
    port map (
            O => \N__61352\,
            I => \N__61336\
        );

    \I__14869\ : LocalMux
    port map (
            O => \N__61349\,
            I => \N__61333\
        );

    \I__14868\ : InMux
    port map (
            O => \N__61348\,
            I => \N__61330\
        );

    \I__14867\ : LocalMux
    port map (
            O => \N__61345\,
            I => \N__61327\
        );

    \I__14866\ : LocalMux
    port map (
            O => \N__61342\,
            I => \N__61320\
        );

    \I__14865\ : LocalMux
    port map (
            O => \N__61339\,
            I => \N__61320\
        );

    \I__14864\ : LocalMux
    port map (
            O => \N__61336\,
            I => \N__61320\
        );

    \I__14863\ : Span4Mux_v
    port map (
            O => \N__61333\,
            I => \N__61311\
        );

    \I__14862\ : LocalMux
    port map (
            O => \N__61330\,
            I => \N__61311\
        );

    \I__14861\ : Span4Mux_v
    port map (
            O => \N__61327\,
            I => \N__61311\
        );

    \I__14860\ : Span4Mux_v
    port map (
            O => \N__61320\,
            I => \N__61307\
        );

    \I__14859\ : InMux
    port map (
            O => \N__61319\,
            I => \N__61304\
        );

    \I__14858\ : InMux
    port map (
            O => \N__61318\,
            I => \N__61301\
        );

    \I__14857\ : Span4Mux_h
    port map (
            O => \N__61311\,
            I => \N__61298\
        );

    \I__14856\ : InMux
    port map (
            O => \N__61310\,
            I => \N__61295\
        );

    \I__14855\ : Span4Mux_h
    port map (
            O => \N__61307\,
            I => \N__61290\
        );

    \I__14854\ : LocalMux
    port map (
            O => \N__61304\,
            I => \N__61290\
        );

    \I__14853\ : LocalMux
    port map (
            O => \N__61301\,
            I => \N__61287\
        );

    \I__14852\ : Span4Mux_h
    port map (
            O => \N__61298\,
            I => \N__61284\
        );

    \I__14851\ : LocalMux
    port map (
            O => \N__61295\,
            I => \N__61281\
        );

    \I__14850\ : Span4Mux_v
    port map (
            O => \N__61290\,
            I => \N__61276\
        );

    \I__14849\ : Span4Mux_h
    port map (
            O => \N__61287\,
            I => \N__61276\
        );

    \I__14848\ : Span4Mux_v
    port map (
            O => \N__61284\,
            I => \N__61273\
        );

    \I__14847\ : Span4Mux_h
    port map (
            O => \N__61281\,
            I => \N__61270\
        );

    \I__14846\ : Span4Mux_v
    port map (
            O => \N__61276\,
            I => \N__61267\
        );

    \I__14845\ : Odrv4
    port map (
            O => \N__61273\,
            I => \I2C_top_level_inst1_s_data_oreg_22\
        );

    \I__14844\ : Odrv4
    port map (
            O => \N__61270\,
            I => \I2C_top_level_inst1_s_data_oreg_22\
        );

    \I__14843\ : Odrv4
    port map (
            O => \N__61267\,
            I => \I2C_top_level_inst1_s_data_oreg_22\
        );

    \I__14842\ : InMux
    port map (
            O => \N__61260\,
            I => \N__61257\
        );

    \I__14841\ : LocalMux
    port map (
            O => \N__61257\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_22\
        );

    \I__14840\ : InMux
    port map (
            O => \N__61254\,
            I => \N__61249\
        );

    \I__14839\ : InMux
    port map (
            O => \N__61253\,
            I => \N__61243\
        );

    \I__14838\ : CascadeMux
    port map (
            O => \N__61252\,
            I => \N__61239\
        );

    \I__14837\ : LocalMux
    port map (
            O => \N__61249\,
            I => \N__61236\
        );

    \I__14836\ : InMux
    port map (
            O => \N__61248\,
            I => \N__61233\
        );

    \I__14835\ : InMux
    port map (
            O => \N__61247\,
            I => \N__61230\
        );

    \I__14834\ : InMux
    port map (
            O => \N__61246\,
            I => \N__61226\
        );

    \I__14833\ : LocalMux
    port map (
            O => \N__61243\,
            I => \N__61223\
        );

    \I__14832\ : InMux
    port map (
            O => \N__61242\,
            I => \N__61220\
        );

    \I__14831\ : InMux
    port map (
            O => \N__61239\,
            I => \N__61217\
        );

    \I__14830\ : Span4Mux_v
    port map (
            O => \N__61236\,
            I => \N__61212\
        );

    \I__14829\ : LocalMux
    port map (
            O => \N__61233\,
            I => \N__61212\
        );

    \I__14828\ : LocalMux
    port map (
            O => \N__61230\,
            I => \N__61209\
        );

    \I__14827\ : InMux
    port map (
            O => \N__61229\,
            I => \N__61206\
        );

    \I__14826\ : LocalMux
    port map (
            O => \N__61226\,
            I => \N__61203\
        );

    \I__14825\ : Span4Mux_v
    port map (
            O => \N__61223\,
            I => \N__61200\
        );

    \I__14824\ : LocalMux
    port map (
            O => \N__61220\,
            I => \N__61197\
        );

    \I__14823\ : LocalMux
    port map (
            O => \N__61217\,
            I => \N__61194\
        );

    \I__14822\ : Span4Mux_v
    port map (
            O => \N__61212\,
            I => \N__61188\
        );

    \I__14821\ : Span4Mux_v
    port map (
            O => \N__61209\,
            I => \N__61188\
        );

    \I__14820\ : LocalMux
    port map (
            O => \N__61206\,
            I => \N__61185\
        );

    \I__14819\ : Span4Mux_v
    port map (
            O => \N__61203\,
            I => \N__61182\
        );

    \I__14818\ : Span4Mux_h
    port map (
            O => \N__61200\,
            I => \N__61177\
        );

    \I__14817\ : Span4Mux_v
    port map (
            O => \N__61197\,
            I => \N__61177\
        );

    \I__14816\ : Span4Mux_v
    port map (
            O => \N__61194\,
            I => \N__61174\
        );

    \I__14815\ : InMux
    port map (
            O => \N__61193\,
            I => \N__61171\
        );

    \I__14814\ : Span4Mux_h
    port map (
            O => \N__61188\,
            I => \N__61166\
        );

    \I__14813\ : Span4Mux_v
    port map (
            O => \N__61185\,
            I => \N__61166\
        );

    \I__14812\ : Span4Mux_h
    port map (
            O => \N__61182\,
            I => \N__61163\
        );

    \I__14811\ : Span4Mux_h
    port map (
            O => \N__61177\,
            I => \N__61158\
        );

    \I__14810\ : Span4Mux_h
    port map (
            O => \N__61174\,
            I => \N__61158\
        );

    \I__14809\ : LocalMux
    port map (
            O => \N__61171\,
            I => \N__61155\
        );

    \I__14808\ : Sp12to4
    port map (
            O => \N__61166\,
            I => \N__61152\
        );

    \I__14807\ : Span4Mux_h
    port map (
            O => \N__61163\,
            I => \N__61149\
        );

    \I__14806\ : Span4Mux_h
    port map (
            O => \N__61158\,
            I => \N__61146\
        );

    \I__14805\ : Odrv12
    port map (
            O => \N__61155\,
            I => \I2C_top_level_inst1_s_data_oreg_23\
        );

    \I__14804\ : Odrv12
    port map (
            O => \N__61152\,
            I => \I2C_top_level_inst1_s_data_oreg_23\
        );

    \I__14803\ : Odrv4
    port map (
            O => \N__61149\,
            I => \I2C_top_level_inst1_s_data_oreg_23\
        );

    \I__14802\ : Odrv4
    port map (
            O => \N__61146\,
            I => \I2C_top_level_inst1_s_data_oreg_23\
        );

    \I__14801\ : InMux
    port map (
            O => \N__61137\,
            I => \N__61134\
        );

    \I__14800\ : LocalMux
    port map (
            O => \N__61134\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_23\
        );

    \I__14799\ : InMux
    port map (
            O => \N__61131\,
            I => \N__61127\
        );

    \I__14798\ : InMux
    port map (
            O => \N__61130\,
            I => \N__61121\
        );

    \I__14797\ : LocalMux
    port map (
            O => \N__61127\,
            I => \N__61118\
        );

    \I__14796\ : InMux
    port map (
            O => \N__61126\,
            I => \N__61114\
        );

    \I__14795\ : InMux
    port map (
            O => \N__61125\,
            I => \N__61110\
        );

    \I__14794\ : InMux
    port map (
            O => \N__61124\,
            I => \N__61107\
        );

    \I__14793\ : LocalMux
    port map (
            O => \N__61121\,
            I => \N__61104\
        );

    \I__14792\ : Span4Mux_v
    port map (
            O => \N__61118\,
            I => \N__61100\
        );

    \I__14791\ : InMux
    port map (
            O => \N__61117\,
            I => \N__61097\
        );

    \I__14790\ : LocalMux
    port map (
            O => \N__61114\,
            I => \N__61094\
        );

    \I__14789\ : InMux
    port map (
            O => \N__61113\,
            I => \N__61091\
        );

    \I__14788\ : LocalMux
    port map (
            O => \N__61110\,
            I => \N__61088\
        );

    \I__14787\ : LocalMux
    port map (
            O => \N__61107\,
            I => \N__61085\
        );

    \I__14786\ : Span4Mux_h
    port map (
            O => \N__61104\,
            I => \N__61082\
        );

    \I__14785\ : InMux
    port map (
            O => \N__61103\,
            I => \N__61079\
        );

    \I__14784\ : Span4Mux_h
    port map (
            O => \N__61100\,
            I => \N__61076\
        );

    \I__14783\ : LocalMux
    port map (
            O => \N__61097\,
            I => \N__61073\
        );

    \I__14782\ : Span4Mux_v
    port map (
            O => \N__61094\,
            I => \N__61070\
        );

    \I__14781\ : LocalMux
    port map (
            O => \N__61091\,
            I => \N__61063\
        );

    \I__14780\ : Span4Mux_v
    port map (
            O => \N__61088\,
            I => \N__61063\
        );

    \I__14779\ : Span4Mux_v
    port map (
            O => \N__61085\,
            I => \N__61063\
        );

    \I__14778\ : Span4Mux_h
    port map (
            O => \N__61082\,
            I => \N__61060\
        );

    \I__14777\ : LocalMux
    port map (
            O => \N__61079\,
            I => \N__61057\
        );

    \I__14776\ : Sp12to4
    port map (
            O => \N__61076\,
            I => \N__61054\
        );

    \I__14775\ : Span4Mux_v
    port map (
            O => \N__61073\,
            I => \N__61051\
        );

    \I__14774\ : Span4Mux_h
    port map (
            O => \N__61070\,
            I => \N__61048\
        );

    \I__14773\ : Span4Mux_h
    port map (
            O => \N__61063\,
            I => \N__61045\
        );

    \I__14772\ : Sp12to4
    port map (
            O => \N__61060\,
            I => \N__61038\
        );

    \I__14771\ : Sp12to4
    port map (
            O => \N__61057\,
            I => \N__61038\
        );

    \I__14770\ : Span12Mux_v
    port map (
            O => \N__61054\,
            I => \N__61038\
        );

    \I__14769\ : Span4Mux_v
    port map (
            O => \N__61051\,
            I => \N__61033\
        );

    \I__14768\ : Span4Mux_h
    port map (
            O => \N__61048\,
            I => \N__61033\
        );

    \I__14767\ : Odrv4
    port map (
            O => \N__61045\,
            I => \I2C_top_level_inst1_s_data_oreg_24\
        );

    \I__14766\ : Odrv12
    port map (
            O => \N__61038\,
            I => \I2C_top_level_inst1_s_data_oreg_24\
        );

    \I__14765\ : Odrv4
    port map (
            O => \N__61033\,
            I => \I2C_top_level_inst1_s_data_oreg_24\
        );

    \I__14764\ : InMux
    port map (
            O => \N__61026\,
            I => \N__61023\
        );

    \I__14763\ : LocalMux
    port map (
            O => \N__61023\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_24\
        );

    \I__14762\ : CascadeMux
    port map (
            O => \N__61020\,
            I => \N__61015\
        );

    \I__14761\ : InMux
    port map (
            O => \N__61019\,
            I => \N__61010\
        );

    \I__14760\ : InMux
    port map (
            O => \N__61018\,
            I => \N__61007\
        );

    \I__14759\ : InMux
    port map (
            O => \N__61015\,
            I => \N__61004\
        );

    \I__14758\ : InMux
    port map (
            O => \N__61014\,
            I => \N__61001\
        );

    \I__14757\ : InMux
    port map (
            O => \N__61013\,
            I => \N__60997\
        );

    \I__14756\ : LocalMux
    port map (
            O => \N__61010\,
            I => \N__60994\
        );

    \I__14755\ : LocalMux
    port map (
            O => \N__61007\,
            I => \N__60991\
        );

    \I__14754\ : LocalMux
    port map (
            O => \N__61004\,
            I => \N__60988\
        );

    \I__14753\ : LocalMux
    port map (
            O => \N__61001\,
            I => \N__60985\
        );

    \I__14752\ : InMux
    port map (
            O => \N__61000\,
            I => \N__60982\
        );

    \I__14751\ : LocalMux
    port map (
            O => \N__60997\,
            I => \N__60977\
        );

    \I__14750\ : Span4Mux_v
    port map (
            O => \N__60994\,
            I => \N__60972\
        );

    \I__14749\ : Span4Mux_v
    port map (
            O => \N__60991\,
            I => \N__60972\
        );

    \I__14748\ : Span4Mux_v
    port map (
            O => \N__60988\,
            I => \N__60967\
        );

    \I__14747\ : Span4Mux_v
    port map (
            O => \N__60985\,
            I => \N__60967\
        );

    \I__14746\ : LocalMux
    port map (
            O => \N__60982\,
            I => \N__60964\
        );

    \I__14745\ : InMux
    port map (
            O => \N__60981\,
            I => \N__60961\
        );

    \I__14744\ : InMux
    port map (
            O => \N__60980\,
            I => \N__60958\
        );

    \I__14743\ : Span4Mux_h
    port map (
            O => \N__60977\,
            I => \N__60955\
        );

    \I__14742\ : Span4Mux_h
    port map (
            O => \N__60972\,
            I => \N__60952\
        );

    \I__14741\ : Sp12to4
    port map (
            O => \N__60967\,
            I => \N__60949\
        );

    \I__14740\ : Span4Mux_v
    port map (
            O => \N__60964\,
            I => \N__60946\
        );

    \I__14739\ : LocalMux
    port map (
            O => \N__60961\,
            I => \N__60939\
        );

    \I__14738\ : LocalMux
    port map (
            O => \N__60958\,
            I => \N__60939\
        );

    \I__14737\ : Span4Mux_v
    port map (
            O => \N__60955\,
            I => \N__60939\
        );

    \I__14736\ : Sp12to4
    port map (
            O => \N__60952\,
            I => \N__60934\
        );

    \I__14735\ : Span12Mux_h
    port map (
            O => \N__60949\,
            I => \N__60934\
        );

    \I__14734\ : Odrv4
    port map (
            O => \N__60946\,
            I => \I2C_top_level_inst1_s_data_oreg_25\
        );

    \I__14733\ : Odrv4
    port map (
            O => \N__60939\,
            I => \I2C_top_level_inst1_s_data_oreg_25\
        );

    \I__14732\ : Odrv12
    port map (
            O => \N__60934\,
            I => \I2C_top_level_inst1_s_data_oreg_25\
        );

    \I__14731\ : InMux
    port map (
            O => \N__60927\,
            I => \N__60924\
        );

    \I__14730\ : LocalMux
    port map (
            O => \N__60924\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_25\
        );

    \I__14729\ : InMux
    port map (
            O => \N__60921\,
            I => \N__60918\
        );

    \I__14728\ : LocalMux
    port map (
            O => \N__60918\,
            I => \N__60915\
        );

    \I__14727\ : Span4Mux_h
    port map (
            O => \N__60915\,
            I => \N__60909\
        );

    \I__14726\ : InMux
    port map (
            O => \N__60914\,
            I => \N__60906\
        );

    \I__14725\ : InMux
    port map (
            O => \N__60913\,
            I => \N__60902\
        );

    \I__14724\ : InMux
    port map (
            O => \N__60912\,
            I => \N__60898\
        );

    \I__14723\ : Span4Mux_h
    port map (
            O => \N__60909\,
            I => \N__60892\
        );

    \I__14722\ : LocalMux
    port map (
            O => \N__60906\,
            I => \N__60892\
        );

    \I__14721\ : InMux
    port map (
            O => \N__60905\,
            I => \N__60889\
        );

    \I__14720\ : LocalMux
    port map (
            O => \N__60902\,
            I => \N__60886\
        );

    \I__14719\ : InMux
    port map (
            O => \N__60901\,
            I => \N__60883\
        );

    \I__14718\ : LocalMux
    port map (
            O => \N__60898\,
            I => \N__60880\
        );

    \I__14717\ : InMux
    port map (
            O => \N__60897\,
            I => \N__60877\
        );

    \I__14716\ : Span4Mux_v
    port map (
            O => \N__60892\,
            I => \N__60872\
        );

    \I__14715\ : LocalMux
    port map (
            O => \N__60889\,
            I => \N__60872\
        );

    \I__14714\ : Span4Mux_h
    port map (
            O => \N__60886\,
            I => \N__60869\
        );

    \I__14713\ : LocalMux
    port map (
            O => \N__60883\,
            I => \N__60866\
        );

    \I__14712\ : Span4Mux_v
    port map (
            O => \N__60880\,
            I => \N__60863\
        );

    \I__14711\ : LocalMux
    port map (
            O => \N__60877\,
            I => \N__60860\
        );

    \I__14710\ : Span4Mux_h
    port map (
            O => \N__60872\,
            I => \N__60857\
        );

    \I__14709\ : Span4Mux_v
    port map (
            O => \N__60869\,
            I => \N__60850\
        );

    \I__14708\ : Span4Mux_v
    port map (
            O => \N__60866\,
            I => \N__60850\
        );

    \I__14707\ : Span4Mux_v
    port map (
            O => \N__60863\,
            I => \N__60850\
        );

    \I__14706\ : Span4Mux_h
    port map (
            O => \N__60860\,
            I => \N__60846\
        );

    \I__14705\ : Sp12to4
    port map (
            O => \N__60857\,
            I => \N__60843\
        );

    \I__14704\ : Sp12to4
    port map (
            O => \N__60850\,
            I => \N__60840\
        );

    \I__14703\ : InMux
    port map (
            O => \N__60849\,
            I => \N__60837\
        );

    \I__14702\ : Span4Mux_v
    port map (
            O => \N__60846\,
            I => \N__60834\
        );

    \I__14701\ : Span12Mux_v
    port map (
            O => \N__60843\,
            I => \N__60829\
        );

    \I__14700\ : Span12Mux_h
    port map (
            O => \N__60840\,
            I => \N__60829\
        );

    \I__14699\ : LocalMux
    port map (
            O => \N__60837\,
            I => \I2C_top_level_inst1_s_data_oreg_26\
        );

    \I__14698\ : Odrv4
    port map (
            O => \N__60834\,
            I => \I2C_top_level_inst1_s_data_oreg_26\
        );

    \I__14697\ : Odrv12
    port map (
            O => \N__60829\,
            I => \I2C_top_level_inst1_s_data_oreg_26\
        );

    \I__14696\ : InMux
    port map (
            O => \N__60822\,
            I => \N__60819\
        );

    \I__14695\ : LocalMux
    port map (
            O => \N__60819\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_26\
        );

    \I__14694\ : CascadeMux
    port map (
            O => \N__60816\,
            I => \N__60813\
        );

    \I__14693\ : InMux
    port map (
            O => \N__60813\,
            I => \N__60810\
        );

    \I__14692\ : LocalMux
    port map (
            O => \N__60810\,
            I => \N__60807\
        );

    \I__14691\ : Span4Mux_v
    port map (
            O => \N__60807\,
            I => \N__60802\
        );

    \I__14690\ : InMux
    port map (
            O => \N__60806\,
            I => \N__60799\
        );

    \I__14689\ : InMux
    port map (
            O => \N__60805\,
            I => \N__60794\
        );

    \I__14688\ : Span4Mux_h
    port map (
            O => \N__60802\,
            I => \N__60791\
        );

    \I__14687\ : LocalMux
    port map (
            O => \N__60799\,
            I => \N__60788\
        );

    \I__14686\ : InMux
    port map (
            O => \N__60798\,
            I => \N__60783\
        );

    \I__14685\ : InMux
    port map (
            O => \N__60797\,
            I => \N__60780\
        );

    \I__14684\ : LocalMux
    port map (
            O => \N__60794\,
            I => \N__60777\
        );

    \I__14683\ : Span4Mux_v
    port map (
            O => \N__60791\,
            I => \N__60771\
        );

    \I__14682\ : Span4Mux_h
    port map (
            O => \N__60788\,
            I => \N__60771\
        );

    \I__14681\ : InMux
    port map (
            O => \N__60787\,
            I => \N__60768\
        );

    \I__14680\ : InMux
    port map (
            O => \N__60786\,
            I => \N__60765\
        );

    \I__14679\ : LocalMux
    port map (
            O => \N__60783\,
            I => \N__60762\
        );

    \I__14678\ : LocalMux
    port map (
            O => \N__60780\,
            I => \N__60759\
        );

    \I__14677\ : Span4Mux_v
    port map (
            O => \N__60777\,
            I => \N__60756\
        );

    \I__14676\ : InMux
    port map (
            O => \N__60776\,
            I => \N__60753\
        );

    \I__14675\ : Span4Mux_v
    port map (
            O => \N__60771\,
            I => \N__60746\
        );

    \I__14674\ : LocalMux
    port map (
            O => \N__60768\,
            I => \N__60746\
        );

    \I__14673\ : LocalMux
    port map (
            O => \N__60765\,
            I => \N__60746\
        );

    \I__14672\ : Span4Mux_h
    port map (
            O => \N__60762\,
            I => \N__60743\
        );

    \I__14671\ : Span4Mux_v
    port map (
            O => \N__60759\,
            I => \N__60740\
        );

    \I__14670\ : Span4Mux_h
    port map (
            O => \N__60756\,
            I => \N__60737\
        );

    \I__14669\ : LocalMux
    port map (
            O => \N__60753\,
            I => \N__60734\
        );

    \I__14668\ : Span4Mux_h
    port map (
            O => \N__60746\,
            I => \N__60731\
        );

    \I__14667\ : Span4Mux_v
    port map (
            O => \N__60743\,
            I => \N__60728\
        );

    \I__14666\ : Span4Mux_v
    port map (
            O => \N__60740\,
            I => \N__60723\
        );

    \I__14665\ : Span4Mux_h
    port map (
            O => \N__60737\,
            I => \N__60723\
        );

    \I__14664\ : Odrv4
    port map (
            O => \N__60734\,
            I => \I2C_top_level_inst1_s_data_oreg_27\
        );

    \I__14663\ : Odrv4
    port map (
            O => \N__60731\,
            I => \I2C_top_level_inst1_s_data_oreg_27\
        );

    \I__14662\ : Odrv4
    port map (
            O => \N__60728\,
            I => \I2C_top_level_inst1_s_data_oreg_27\
        );

    \I__14661\ : Odrv4
    port map (
            O => \N__60723\,
            I => \I2C_top_level_inst1_s_data_oreg_27\
        );

    \I__14660\ : InMux
    port map (
            O => \N__60714\,
            I => \N__60711\
        );

    \I__14659\ : LocalMux
    port map (
            O => \N__60711\,
            I => \N__60706\
        );

    \I__14658\ : InMux
    port map (
            O => \N__60710\,
            I => \N__60703\
        );

    \I__14657\ : CascadeMux
    port map (
            O => \N__60709\,
            I => \N__60700\
        );

    \I__14656\ : Span4Mux_h
    port map (
            O => \N__60706\,
            I => \N__60697\
        );

    \I__14655\ : LocalMux
    port map (
            O => \N__60703\,
            I => \N__60694\
        );

    \I__14654\ : InMux
    port map (
            O => \N__60700\,
            I => \N__60691\
        );

    \I__14653\ : Span4Mux_h
    port map (
            O => \N__60697\,
            I => \N__60688\
        );

    \I__14652\ : Span4Mux_h
    port map (
            O => \N__60694\,
            I => \N__60683\
        );

    \I__14651\ : LocalMux
    port map (
            O => \N__60691\,
            I => \N__60683\
        );

    \I__14650\ : Odrv4
    port map (
            O => \N__60688\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_1
        );

    \I__14649\ : Odrv4
    port map (
            O => \N__60683\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_1
        );

    \I__14648\ : CascadeMux
    port map (
            O => \N__60678\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_1_cascade_\
        );

    \I__14647\ : InMux
    port map (
            O => \N__60675\,
            I => \N__60672\
        );

    \I__14646\ : LocalMux
    port map (
            O => \N__60672\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_1\
        );

    \I__14645\ : CascadeMux
    port map (
            O => \N__60669\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2QZ0Z5_cascade_\
        );

    \I__14644\ : InMux
    port map (
            O => \N__60666\,
            I => \N__60663\
        );

    \I__14643\ : LocalMux
    port map (
            O => \N__60663\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1\
        );

    \I__14642\ : CascadeMux
    port map (
            O => \N__60660\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_cascade_\
        );

    \I__14641\ : InMux
    port map (
            O => \N__60657\,
            I => \N__60654\
        );

    \I__14640\ : LocalMux
    port map (
            O => \N__60654\,
            I => \N__60651\
        );

    \I__14639\ : Span4Mux_h
    port map (
            O => \N__60651\,
            I => \N__60648\
        );

    \I__14638\ : Odrv4
    port map (
            O => \N__60648\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_1\
        );

    \I__14637\ : InMux
    port map (
            O => \N__60645\,
            I => \N__60642\
        );

    \I__14636\ : LocalMux
    port map (
            O => \N__60642\,
            I => \N__60637\
        );

    \I__14635\ : InMux
    port map (
            O => \N__60641\,
            I => \N__60634\
        );

    \I__14634\ : InMux
    port map (
            O => \N__60640\,
            I => \N__60631\
        );

    \I__14633\ : Span4Mux_v
    port map (
            O => \N__60637\,
            I => \N__60626\
        );

    \I__14632\ : LocalMux
    port map (
            O => \N__60634\,
            I => \N__60626\
        );

    \I__14631\ : LocalMux
    port map (
            O => \N__60631\,
            I => \N__60623\
        );

    \I__14630\ : Odrv4
    port map (
            O => \N__60626\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_0
        );

    \I__14629\ : Odrv4
    port map (
            O => \N__60623\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_0
        );

    \I__14628\ : InMux
    port map (
            O => \N__60618\,
            I => \N__60609\
        );

    \I__14627\ : InMux
    port map (
            O => \N__60617\,
            I => \N__60606\
        );

    \I__14626\ : InMux
    port map (
            O => \N__60616\,
            I => \N__60599\
        );

    \I__14625\ : InMux
    port map (
            O => \N__60615\,
            I => \N__60599\
        );

    \I__14624\ : InMux
    port map (
            O => \N__60614\,
            I => \N__60592\
        );

    \I__14623\ : InMux
    port map (
            O => \N__60613\,
            I => \N__60592\
        );

    \I__14622\ : InMux
    port map (
            O => \N__60612\,
            I => \N__60586\
        );

    \I__14621\ : LocalMux
    port map (
            O => \N__60609\,
            I => \N__60581\
        );

    \I__14620\ : LocalMux
    port map (
            O => \N__60606\,
            I => \N__60581\
        );

    \I__14619\ : InMux
    port map (
            O => \N__60605\,
            I => \N__60578\
        );

    \I__14618\ : InMux
    port map (
            O => \N__60604\,
            I => \N__60575\
        );

    \I__14617\ : LocalMux
    port map (
            O => \N__60599\,
            I => \N__60572\
        );

    \I__14616\ : InMux
    port map (
            O => \N__60598\,
            I => \N__60569\
        );

    \I__14615\ : InMux
    port map (
            O => \N__60597\,
            I => \N__60566\
        );

    \I__14614\ : LocalMux
    port map (
            O => \N__60592\,
            I => \N__60562\
        );

    \I__14613\ : InMux
    port map (
            O => \N__60591\,
            I => \N__60559\
        );

    \I__14612\ : InMux
    port map (
            O => \N__60590\,
            I => \N__60552\
        );

    \I__14611\ : InMux
    port map (
            O => \N__60589\,
            I => \N__60552\
        );

    \I__14610\ : LocalMux
    port map (
            O => \N__60586\,
            I => \N__60549\
        );

    \I__14609\ : Span4Mux_h
    port map (
            O => \N__60581\,
            I => \N__60544\
        );

    \I__14608\ : LocalMux
    port map (
            O => \N__60578\,
            I => \N__60544\
        );

    \I__14607\ : LocalMux
    port map (
            O => \N__60575\,
            I => \N__60541\
        );

    \I__14606\ : Span4Mux_v
    port map (
            O => \N__60572\,
            I => \N__60535\
        );

    \I__14605\ : LocalMux
    port map (
            O => \N__60569\,
            I => \N__60535\
        );

    \I__14604\ : LocalMux
    port map (
            O => \N__60566\,
            I => \N__60532\
        );

    \I__14603\ : InMux
    port map (
            O => \N__60565\,
            I => \N__60529\
        );

    \I__14602\ : Span4Mux_h
    port map (
            O => \N__60562\,
            I => \N__60524\
        );

    \I__14601\ : LocalMux
    port map (
            O => \N__60559\,
            I => \N__60524\
        );

    \I__14600\ : InMux
    port map (
            O => \N__60558\,
            I => \N__60521\
        );

    \I__14599\ : InMux
    port map (
            O => \N__60557\,
            I => \N__60518\
        );

    \I__14598\ : LocalMux
    port map (
            O => \N__60552\,
            I => \N__60512\
        );

    \I__14597\ : Span4Mux_v
    port map (
            O => \N__60549\,
            I => \N__60507\
        );

    \I__14596\ : Span4Mux_v
    port map (
            O => \N__60544\,
            I => \N__60507\
        );

    \I__14595\ : Span4Mux_h
    port map (
            O => \N__60541\,
            I => \N__60504\
        );

    \I__14594\ : InMux
    port map (
            O => \N__60540\,
            I => \N__60501\
        );

    \I__14593\ : Span4Mux_h
    port map (
            O => \N__60535\,
            I => \N__60496\
        );

    \I__14592\ : Span4Mux_v
    port map (
            O => \N__60532\,
            I => \N__60496\
        );

    \I__14591\ : LocalMux
    port map (
            O => \N__60529\,
            I => \N__60489\
        );

    \I__14590\ : Span4Mux_h
    port map (
            O => \N__60524\,
            I => \N__60489\
        );

    \I__14589\ : LocalMux
    port map (
            O => \N__60521\,
            I => \N__60489\
        );

    \I__14588\ : LocalMux
    port map (
            O => \N__60518\,
            I => \N__60486\
        );

    \I__14587\ : InMux
    port map (
            O => \N__60517\,
            I => \N__60483\
        );

    \I__14586\ : InMux
    port map (
            O => \N__60516\,
            I => \N__60478\
        );

    \I__14585\ : InMux
    port map (
            O => \N__60515\,
            I => \N__60478\
        );

    \I__14584\ : Span4Mux_v
    port map (
            O => \N__60512\,
            I => \N__60475\
        );

    \I__14583\ : Span4Mux_h
    port map (
            O => \N__60507\,
            I => \N__60469\
        );

    \I__14582\ : Span4Mux_h
    port map (
            O => \N__60504\,
            I => \N__60464\
        );

    \I__14581\ : LocalMux
    port map (
            O => \N__60501\,
            I => \N__60464\
        );

    \I__14580\ : Span4Mux_h
    port map (
            O => \N__60496\,
            I => \N__60461\
        );

    \I__14579\ : Span4Mux_v
    port map (
            O => \N__60489\,
            I => \N__60456\
        );

    \I__14578\ : Span4Mux_h
    port map (
            O => \N__60486\,
            I => \N__60456\
        );

    \I__14577\ : LocalMux
    port map (
            O => \N__60483\,
            I => \N__60451\
        );

    \I__14576\ : LocalMux
    port map (
            O => \N__60478\,
            I => \N__60451\
        );

    \I__14575\ : Sp12to4
    port map (
            O => \N__60475\,
            I => \N__60448\
        );

    \I__14574\ : InMux
    port map (
            O => \N__60474\,
            I => \N__60445\
        );

    \I__14573\ : InMux
    port map (
            O => \N__60473\,
            I => \N__60440\
        );

    \I__14572\ : InMux
    port map (
            O => \N__60472\,
            I => \N__60440\
        );

    \I__14571\ : Span4Mux_h
    port map (
            O => \N__60469\,
            I => \N__60435\
        );

    \I__14570\ : Span4Mux_v
    port map (
            O => \N__60464\,
            I => \N__60435\
        );

    \I__14569\ : Span4Mux_h
    port map (
            O => \N__60461\,
            I => \N__60430\
        );

    \I__14568\ : Span4Mux_h
    port map (
            O => \N__60456\,
            I => \N__60430\
        );

    \I__14567\ : Span12Mux_v
    port map (
            O => \N__60451\,
            I => \N__60427\
        );

    \I__14566\ : Span12Mux_h
    port map (
            O => \N__60448\,
            I => \N__60420\
        );

    \I__14565\ : LocalMux
    port map (
            O => \N__60445\,
            I => \N__60420\
        );

    \I__14564\ : LocalMux
    port map (
            O => \N__60440\,
            I => \N__60420\
        );

    \I__14563\ : Odrv4
    port map (
            O => \N__60435\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340\
        );

    \I__14562\ : Odrv4
    port map (
            O => \N__60430\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340\
        );

    \I__14561\ : Odrv12
    port map (
            O => \N__60427\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340\
        );

    \I__14560\ : Odrv12
    port map (
            O => \N__60420\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340\
        );

    \I__14559\ : CascadeMux
    port map (
            O => \N__60411\,
            I => \N__60408\
        );

    \I__14558\ : InMux
    port map (
            O => \N__60408\,
            I => \N__60405\
        );

    \I__14557\ : LocalMux
    port map (
            O => \N__60405\,
            I => \N__60402\
        );

    \I__14556\ : Span4Mux_v
    port map (
            O => \N__60402\,
            I => \N__60399\
        );

    \I__14555\ : Span4Mux_h
    port map (
            O => \N__60399\,
            I => \N__60396\
        );

    \I__14554\ : Odrv4
    port map (
            O => \N__60396\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_0\
        );

    \I__14553\ : InMux
    port map (
            O => \N__60393\,
            I => \N__60390\
        );

    \I__14552\ : LocalMux
    port map (
            O => \N__60390\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_0\
        );

    \I__14551\ : InMux
    port map (
            O => \N__60387\,
            I => \N__60369\
        );

    \I__14550\ : InMux
    port map (
            O => \N__60386\,
            I => \N__60369\
        );

    \I__14549\ : InMux
    port map (
            O => \N__60385\,
            I => \N__60364\
        );

    \I__14548\ : InMux
    port map (
            O => \N__60384\,
            I => \N__60364\
        );

    \I__14547\ : InMux
    port map (
            O => \N__60383\,
            I => \N__60359\
        );

    \I__14546\ : InMux
    port map (
            O => \N__60382\,
            I => \N__60359\
        );

    \I__14545\ : InMux
    port map (
            O => \N__60381\,
            I => \N__60350\
        );

    \I__14544\ : InMux
    port map (
            O => \N__60380\,
            I => \N__60347\
        );

    \I__14543\ : InMux
    port map (
            O => \N__60379\,
            I => \N__60340\
        );

    \I__14542\ : InMux
    port map (
            O => \N__60378\,
            I => \N__60340\
        );

    \I__14541\ : InMux
    port map (
            O => \N__60377\,
            I => \N__60335\
        );

    \I__14540\ : InMux
    port map (
            O => \N__60376\,
            I => \N__60335\
        );

    \I__14539\ : InMux
    port map (
            O => \N__60375\,
            I => \N__60330\
        );

    \I__14538\ : InMux
    port map (
            O => \N__60374\,
            I => \N__60330\
        );

    \I__14537\ : LocalMux
    port map (
            O => \N__60369\,
            I => \N__60325\
        );

    \I__14536\ : LocalMux
    port map (
            O => \N__60364\,
            I => \N__60320\
        );

    \I__14535\ : LocalMux
    port map (
            O => \N__60359\,
            I => \N__60320\
        );

    \I__14534\ : InMux
    port map (
            O => \N__60358\,
            I => \N__60317\
        );

    \I__14533\ : InMux
    port map (
            O => \N__60357\,
            I => \N__60312\
        );

    \I__14532\ : InMux
    port map (
            O => \N__60356\,
            I => \N__60312\
        );

    \I__14531\ : InMux
    port map (
            O => \N__60355\,
            I => \N__60307\
        );

    \I__14530\ : InMux
    port map (
            O => \N__60354\,
            I => \N__60307\
        );

    \I__14529\ : InMux
    port map (
            O => \N__60353\,
            I => \N__60304\
        );

    \I__14528\ : LocalMux
    port map (
            O => \N__60350\,
            I => \N__60299\
        );

    \I__14527\ : LocalMux
    port map (
            O => \N__60347\,
            I => \N__60299\
        );

    \I__14526\ : InMux
    port map (
            O => \N__60346\,
            I => \N__60294\
        );

    \I__14525\ : InMux
    port map (
            O => \N__60345\,
            I => \N__60294\
        );

    \I__14524\ : LocalMux
    port map (
            O => \N__60340\,
            I => \N__60287\
        );

    \I__14523\ : LocalMux
    port map (
            O => \N__60335\,
            I => \N__60287\
        );

    \I__14522\ : LocalMux
    port map (
            O => \N__60330\,
            I => \N__60287\
        );

    \I__14521\ : InMux
    port map (
            O => \N__60329\,
            I => \N__60282\
        );

    \I__14520\ : InMux
    port map (
            O => \N__60328\,
            I => \N__60282\
        );

    \I__14519\ : Span4Mux_h
    port map (
            O => \N__60325\,
            I => \N__60277\
        );

    \I__14518\ : Span4Mux_v
    port map (
            O => \N__60320\,
            I => \N__60277\
        );

    \I__14517\ : LocalMux
    port map (
            O => \N__60317\,
            I => \N__60272\
        );

    \I__14516\ : LocalMux
    port map (
            O => \N__60312\,
            I => \N__60272\
        );

    \I__14515\ : LocalMux
    port map (
            O => \N__60307\,
            I => \N__60269\
        );

    \I__14514\ : LocalMux
    port map (
            O => \N__60304\,
            I => \N__60266\
        );

    \I__14513\ : Span4Mux_v
    port map (
            O => \N__60299\,
            I => \N__60263\
        );

    \I__14512\ : LocalMux
    port map (
            O => \N__60294\,
            I => \N__60260\
        );

    \I__14511\ : Span4Mux_v
    port map (
            O => \N__60287\,
            I => \N__60257\
        );

    \I__14510\ : LocalMux
    port map (
            O => \N__60282\,
            I => \N__60254\
        );

    \I__14509\ : Span4Mux_h
    port map (
            O => \N__60277\,
            I => \N__60249\
        );

    \I__14508\ : Span4Mux_v
    port map (
            O => \N__60272\,
            I => \N__60249\
        );

    \I__14507\ : Sp12to4
    port map (
            O => \N__60269\,
            I => \N__60246\
        );

    \I__14506\ : Span12Mux_v
    port map (
            O => \N__60266\,
            I => \N__60243\
        );

    \I__14505\ : Span4Mux_v
    port map (
            O => \N__60263\,
            I => \N__60240\
        );

    \I__14504\ : Sp12to4
    port map (
            O => \N__60260\,
            I => \N__60235\
        );

    \I__14503\ : Sp12to4
    port map (
            O => \N__60257\,
            I => \N__60235\
        );

    \I__14502\ : Span4Mux_h
    port map (
            O => \N__60254\,
            I => \N__60230\
        );

    \I__14501\ : Span4Mux_h
    port map (
            O => \N__60249\,
            I => \N__60230\
        );

    \I__14500\ : Odrv12
    port map (
            O => \N__60246\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\
        );

    \I__14499\ : Odrv12
    port map (
            O => \N__60243\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\
        );

    \I__14498\ : Odrv4
    port map (
            O => \N__60240\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\
        );

    \I__14497\ : Odrv12
    port map (
            O => \N__60235\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\
        );

    \I__14496\ : Odrv4
    port map (
            O => \N__60230\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\
        );

    \I__14495\ : CascadeMux
    port map (
            O => \N__60219\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2QZ0Z5_cascade_\
        );

    \I__14494\ : InMux
    port map (
            O => \N__60216\,
            I => \N__60213\
        );

    \I__14493\ : LocalMux
    port map (
            O => \N__60213\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0\
        );

    \I__14492\ : CascadeMux
    port map (
            O => \N__60210\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0_cascade_\
        );

    \I__14491\ : InMux
    port map (
            O => \N__60207\,
            I => \N__60197\
        );

    \I__14490\ : InMux
    port map (
            O => \N__60206\,
            I => \N__60197\
        );

    \I__14489\ : InMux
    port map (
            O => \N__60205\,
            I => \N__60188\
        );

    \I__14488\ : InMux
    port map (
            O => \N__60204\,
            I => \N__60188\
        );

    \I__14487\ : InMux
    port map (
            O => \N__60203\,
            I => \N__60181\
        );

    \I__14486\ : InMux
    port map (
            O => \N__60202\,
            I => \N__60181\
        );

    \I__14485\ : LocalMux
    port map (
            O => \N__60197\,
            I => \N__60178\
        );

    \I__14484\ : InMux
    port map (
            O => \N__60196\,
            I => \N__60173\
        );

    \I__14483\ : InMux
    port map (
            O => \N__60195\,
            I => \N__60173\
        );

    \I__14482\ : InMux
    port map (
            O => \N__60194\,
            I => \N__60168\
        );

    \I__14481\ : InMux
    port map (
            O => \N__60193\,
            I => \N__60168\
        );

    \I__14480\ : LocalMux
    port map (
            O => \N__60188\,
            I => \N__60159\
        );

    \I__14479\ : InMux
    port map (
            O => \N__60187\,
            I => \N__60152\
        );

    \I__14478\ : InMux
    port map (
            O => \N__60186\,
            I => \N__60152\
        );

    \I__14477\ : LocalMux
    port map (
            O => \N__60181\,
            I => \N__60145\
        );

    \I__14476\ : Span4Mux_v
    port map (
            O => \N__60178\,
            I => \N__60138\
        );

    \I__14475\ : LocalMux
    port map (
            O => \N__60173\,
            I => \N__60138\
        );

    \I__14474\ : LocalMux
    port map (
            O => \N__60168\,
            I => \N__60138\
        );

    \I__14473\ : InMux
    port map (
            O => \N__60167\,
            I => \N__60133\
        );

    \I__14472\ : InMux
    port map (
            O => \N__60166\,
            I => \N__60133\
        );

    \I__14471\ : InMux
    port map (
            O => \N__60165\,
            I => \N__60128\
        );

    \I__14470\ : InMux
    port map (
            O => \N__60164\,
            I => \N__60128\
        );

    \I__14469\ : InMux
    port map (
            O => \N__60163\,
            I => \N__60122\
        );

    \I__14468\ : InMux
    port map (
            O => \N__60162\,
            I => \N__60122\
        );

    \I__14467\ : Span4Mux_v
    port map (
            O => \N__60159\,
            I => \N__60119\
        );

    \I__14466\ : InMux
    port map (
            O => \N__60158\,
            I => \N__60114\
        );

    \I__14465\ : InMux
    port map (
            O => \N__60157\,
            I => \N__60114\
        );

    \I__14464\ : LocalMux
    port map (
            O => \N__60152\,
            I => \N__60111\
        );

    \I__14463\ : InMux
    port map (
            O => \N__60151\,
            I => \N__60106\
        );

    \I__14462\ : InMux
    port map (
            O => \N__60150\,
            I => \N__60106\
        );

    \I__14461\ : InMux
    port map (
            O => \N__60149\,
            I => \N__60101\
        );

    \I__14460\ : InMux
    port map (
            O => \N__60148\,
            I => \N__60101\
        );

    \I__14459\ : Span4Mux_v
    port map (
            O => \N__60145\,
            I => \N__60098\
        );

    \I__14458\ : Span4Mux_v
    port map (
            O => \N__60138\,
            I => \N__60093\
        );

    \I__14457\ : LocalMux
    port map (
            O => \N__60133\,
            I => \N__60093\
        );

    \I__14456\ : LocalMux
    port map (
            O => \N__60128\,
            I => \N__60090\
        );

    \I__14455\ : InMux
    port map (
            O => \N__60127\,
            I => \N__60087\
        );

    \I__14454\ : LocalMux
    port map (
            O => \N__60122\,
            I => \N__60084\
        );

    \I__14453\ : Span4Mux_h
    port map (
            O => \N__60119\,
            I => \N__60081\
        );

    \I__14452\ : LocalMux
    port map (
            O => \N__60114\,
            I => \N__60078\
        );

    \I__14451\ : Span4Mux_h
    port map (
            O => \N__60111\,
            I => \N__60073\
        );

    \I__14450\ : LocalMux
    port map (
            O => \N__60106\,
            I => \N__60073\
        );

    \I__14449\ : LocalMux
    port map (
            O => \N__60101\,
            I => \N__60070\
        );

    \I__14448\ : Span4Mux_v
    port map (
            O => \N__60098\,
            I => \N__60063\
        );

    \I__14447\ : Span4Mux_h
    port map (
            O => \N__60093\,
            I => \N__60063\
        );

    \I__14446\ : Span4Mux_v
    port map (
            O => \N__60090\,
            I => \N__60063\
        );

    \I__14445\ : LocalMux
    port map (
            O => \N__60087\,
            I => \N__60060\
        );

    \I__14444\ : Span12Mux_v
    port map (
            O => \N__60084\,
            I => \N__60057\
        );

    \I__14443\ : Span4Mux_h
    port map (
            O => \N__60081\,
            I => \N__60054\
        );

    \I__14442\ : Span4Mux_v
    port map (
            O => \N__60078\,
            I => \N__60051\
        );

    \I__14441\ : Span4Mux_v
    port map (
            O => \N__60073\,
            I => \N__60046\
        );

    \I__14440\ : Span4Mux_h
    port map (
            O => \N__60070\,
            I => \N__60046\
        );

    \I__14439\ : Span4Mux_h
    port map (
            O => \N__60063\,
            I => \N__60041\
        );

    \I__14438\ : Span4Mux_h
    port map (
            O => \N__60060\,
            I => \N__60041\
        );

    \I__14437\ : Odrv12
    port map (
            O => \N__60057\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\
        );

    \I__14436\ : Odrv4
    port map (
            O => \N__60054\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\
        );

    \I__14435\ : Odrv4
    port map (
            O => \N__60051\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\
        );

    \I__14434\ : Odrv4
    port map (
            O => \N__60046\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\
        );

    \I__14433\ : Odrv4
    port map (
            O => \N__60041\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\
        );

    \I__14432\ : InMux
    port map (
            O => \N__60030\,
            I => \N__60027\
        );

    \I__14431\ : LocalMux
    port map (
            O => \N__60027\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_0\
        );

    \I__14430\ : CEMux
    port map (
            O => \N__60024\,
            I => \N__60019\
        );

    \I__14429\ : CEMux
    port map (
            O => \N__60023\,
            I => \N__60013\
        );

    \I__14428\ : CEMux
    port map (
            O => \N__60022\,
            I => \N__60010\
        );

    \I__14427\ : LocalMux
    port map (
            O => \N__60019\,
            I => \N__60006\
        );

    \I__14426\ : CEMux
    port map (
            O => \N__60018\,
            I => \N__60001\
        );

    \I__14425\ : CEMux
    port map (
            O => \N__60017\,
            I => \N__59998\
        );

    \I__14424\ : CEMux
    port map (
            O => \N__60016\,
            I => \N__59995\
        );

    \I__14423\ : LocalMux
    port map (
            O => \N__60013\,
            I => \N__59991\
        );

    \I__14422\ : LocalMux
    port map (
            O => \N__60010\,
            I => \N__59988\
        );

    \I__14421\ : CEMux
    port map (
            O => \N__60009\,
            I => \N__59985\
        );

    \I__14420\ : Span4Mux_h
    port map (
            O => \N__60006\,
            I => \N__59981\
        );

    \I__14419\ : CEMux
    port map (
            O => \N__60005\,
            I => \N__59978\
        );

    \I__14418\ : CEMux
    port map (
            O => \N__60004\,
            I => \N__59975\
        );

    \I__14417\ : LocalMux
    port map (
            O => \N__60001\,
            I => \N__59972\
        );

    \I__14416\ : LocalMux
    port map (
            O => \N__59998\,
            I => \N__59969\
        );

    \I__14415\ : LocalMux
    port map (
            O => \N__59995\,
            I => \N__59966\
        );

    \I__14414\ : CEMux
    port map (
            O => \N__59994\,
            I => \N__59963\
        );

    \I__14413\ : Span4Mux_v
    port map (
            O => \N__59991\,
            I => \N__59958\
        );

    \I__14412\ : Span4Mux_v
    port map (
            O => \N__59988\,
            I => \N__59958\
        );

    \I__14411\ : LocalMux
    port map (
            O => \N__59985\,
            I => \N__59955\
        );

    \I__14410\ : CEMux
    port map (
            O => \N__59984\,
            I => \N__59952\
        );

    \I__14409\ : Span4Mux_h
    port map (
            O => \N__59981\,
            I => \N__59947\
        );

    \I__14408\ : LocalMux
    port map (
            O => \N__59978\,
            I => \N__59947\
        );

    \I__14407\ : LocalMux
    port map (
            O => \N__59975\,
            I => \N__59944\
        );

    \I__14406\ : Span4Mux_h
    port map (
            O => \N__59972\,
            I => \N__59941\
        );

    \I__14405\ : Span4Mux_v
    port map (
            O => \N__59969\,
            I => \N__59935\
        );

    \I__14404\ : Span4Mux_v
    port map (
            O => \N__59966\,
            I => \N__59935\
        );

    \I__14403\ : LocalMux
    port map (
            O => \N__59963\,
            I => \N__59932\
        );

    \I__14402\ : Span4Mux_h
    port map (
            O => \N__59958\,
            I => \N__59929\
        );

    \I__14401\ : Span4Mux_v
    port map (
            O => \N__59955\,
            I => \N__59926\
        );

    \I__14400\ : LocalMux
    port map (
            O => \N__59952\,
            I => \N__59923\
        );

    \I__14399\ : Span4Mux_h
    port map (
            O => \N__59947\,
            I => \N__59920\
        );

    \I__14398\ : Span4Mux_v
    port map (
            O => \N__59944\,
            I => \N__59917\
        );

    \I__14397\ : Span4Mux_h
    port map (
            O => \N__59941\,
            I => \N__59914\
        );

    \I__14396\ : CEMux
    port map (
            O => \N__59940\,
            I => \N__59911\
        );

    \I__14395\ : Sp12to4
    port map (
            O => \N__59935\,
            I => \N__59906\
        );

    \I__14394\ : Sp12to4
    port map (
            O => \N__59932\,
            I => \N__59906\
        );

    \I__14393\ : Span4Mux_h
    port map (
            O => \N__59929\,
            I => \N__59901\
        );

    \I__14392\ : Span4Mux_v
    port map (
            O => \N__59926\,
            I => \N__59901\
        );

    \I__14391\ : Span4Mux_h
    port map (
            O => \N__59923\,
            I => \N__59896\
        );

    \I__14390\ : Span4Mux_v
    port map (
            O => \N__59920\,
            I => \N__59896\
        );

    \I__14389\ : Span4Mux_h
    port map (
            O => \N__59917\,
            I => \N__59893\
        );

    \I__14388\ : Span4Mux_h
    port map (
            O => \N__59914\,
            I => \N__59888\
        );

    \I__14387\ : LocalMux
    port map (
            O => \N__59911\,
            I => \N__59888\
        );

    \I__14386\ : Span12Mux_h
    port map (
            O => \N__59906\,
            I => \N__59885\
        );

    \I__14385\ : Span4Mux_h
    port map (
            O => \N__59901\,
            I => \N__59882\
        );

    \I__14384\ : Span4Mux_h
    port map (
            O => \N__59896\,
            I => \N__59879\
        );

    \I__14383\ : Span4Mux_v
    port map (
            O => \N__59893\,
            I => \N__59874\
        );

    \I__14382\ : Span4Mux_v
    port map (
            O => \N__59888\,
            I => \N__59874\
        );

    \I__14381\ : Odrv12
    port map (
            O => \N__59885\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i\
        );

    \I__14380\ : Odrv4
    port map (
            O => \N__59882\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i\
        );

    \I__14379\ : Odrv4
    port map (
            O => \N__59879\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i\
        );

    \I__14378\ : Odrv4
    port map (
            O => \N__59874\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i\
        );

    \I__14377\ : InMux
    port map (
            O => \N__59865\,
            I => \N__59860\
        );

    \I__14376\ : InMux
    port map (
            O => \N__59864\,
            I => \N__59857\
        );

    \I__14375\ : InMux
    port map (
            O => \N__59863\,
            I => \N__59854\
        );

    \I__14374\ : LocalMux
    port map (
            O => \N__59860\,
            I => \N__59845\
        );

    \I__14373\ : LocalMux
    port map (
            O => \N__59857\,
            I => \N__59845\
        );

    \I__14372\ : LocalMux
    port map (
            O => \N__59854\,
            I => \N__59841\
        );

    \I__14371\ : InMux
    port map (
            O => \N__59853\,
            I => \N__59838\
        );

    \I__14370\ : InMux
    port map (
            O => \N__59852\,
            I => \N__59835\
        );

    \I__14369\ : InMux
    port map (
            O => \N__59851\,
            I => \N__59831\
        );

    \I__14368\ : InMux
    port map (
            O => \N__59850\,
            I => \N__59828\
        );

    \I__14367\ : Span4Mux_v
    port map (
            O => \N__59845\,
            I => \N__59825\
        );

    \I__14366\ : InMux
    port map (
            O => \N__59844\,
            I => \N__59822\
        );

    \I__14365\ : Span4Mux_h
    port map (
            O => \N__59841\,
            I => \N__59817\
        );

    \I__14364\ : LocalMux
    port map (
            O => \N__59838\,
            I => \N__59817\
        );

    \I__14363\ : LocalMux
    port map (
            O => \N__59835\,
            I => \N__59814\
        );

    \I__14362\ : InMux
    port map (
            O => \N__59834\,
            I => \N__59811\
        );

    \I__14361\ : LocalMux
    port map (
            O => \N__59831\,
            I => \N__59808\
        );

    \I__14360\ : LocalMux
    port map (
            O => \N__59828\,
            I => \N__59805\
        );

    \I__14359\ : Span4Mux_h
    port map (
            O => \N__59825\,
            I => \N__59802\
        );

    \I__14358\ : LocalMux
    port map (
            O => \N__59822\,
            I => \N__59797\
        );

    \I__14357\ : Span4Mux_v
    port map (
            O => \N__59817\,
            I => \N__59797\
        );

    \I__14356\ : Span4Mux_h
    port map (
            O => \N__59814\,
            I => \N__59794\
        );

    \I__14355\ : LocalMux
    port map (
            O => \N__59811\,
            I => \N__59791\
        );

    \I__14354\ : Span4Mux_v
    port map (
            O => \N__59808\,
            I => \N__59788\
        );

    \I__14353\ : Span4Mux_v
    port map (
            O => \N__59805\,
            I => \N__59783\
        );

    \I__14352\ : Span4Mux_h
    port map (
            O => \N__59802\,
            I => \N__59783\
        );

    \I__14351\ : Span4Mux_h
    port map (
            O => \N__59797\,
            I => \N__59780\
        );

    \I__14350\ : Span4Mux_h
    port map (
            O => \N__59794\,
            I => \N__59775\
        );

    \I__14349\ : Span4Mux_h
    port map (
            O => \N__59791\,
            I => \N__59775\
        );

    \I__14348\ : Span4Mux_h
    port map (
            O => \N__59788\,
            I => \N__59772\
        );

    \I__14347\ : Odrv4
    port map (
            O => \N__59783\,
            I => \I2C_top_level_inst1_s_data_oreg_18\
        );

    \I__14346\ : Odrv4
    port map (
            O => \N__59780\,
            I => \I2C_top_level_inst1_s_data_oreg_18\
        );

    \I__14345\ : Odrv4
    port map (
            O => \N__59775\,
            I => \I2C_top_level_inst1_s_data_oreg_18\
        );

    \I__14344\ : Odrv4
    port map (
            O => \N__59772\,
            I => \I2C_top_level_inst1_s_data_oreg_18\
        );

    \I__14343\ : InMux
    port map (
            O => \N__59763\,
            I => \N__59760\
        );

    \I__14342\ : LocalMux
    port map (
            O => \N__59760\,
            I => \N__59757\
        );

    \I__14341\ : Odrv12
    port map (
            O => \N__59757\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_17\
        );

    \I__14340\ : InMux
    port map (
            O => \N__59754\,
            I => \N__59751\
        );

    \I__14339\ : LocalMux
    port map (
            O => \N__59751\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_18\
        );

    \I__14338\ : CascadeMux
    port map (
            O => \N__59748\,
            I => \N__59745\
        );

    \I__14337\ : InMux
    port map (
            O => \N__59745\,
            I => \N__59742\
        );

    \I__14336\ : LocalMux
    port map (
            O => \N__59742\,
            I => \N__59739\
        );

    \I__14335\ : Span4Mux_h
    port map (
            O => \N__59739\,
            I => \N__59736\
        );

    \I__14334\ : Span4Mux_h
    port map (
            O => \N__59736\,
            I => \N__59733\
        );

    \I__14333\ : Odrv4
    port map (
            O => \N__59733\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_29\
        );

    \I__14332\ : CascadeMux
    port map (
            O => \N__59730\,
            I => \N__59723\
        );

    \I__14331\ : CascadeMux
    port map (
            O => \N__59729\,
            I => \N__59720\
        );

    \I__14330\ : CascadeMux
    port map (
            O => \N__59728\,
            I => \N__59699\
        );

    \I__14329\ : InMux
    port map (
            O => \N__59727\,
            I => \N__59690\
        );

    \I__14328\ : InMux
    port map (
            O => \N__59726\,
            I => \N__59690\
        );

    \I__14327\ : InMux
    port map (
            O => \N__59723\,
            I => \N__59677\
        );

    \I__14326\ : InMux
    port map (
            O => \N__59720\,
            I => \N__59677\
        );

    \I__14325\ : InMux
    port map (
            O => \N__59719\,
            I => \N__59677\
        );

    \I__14324\ : InMux
    port map (
            O => \N__59718\,
            I => \N__59677\
        );

    \I__14323\ : InMux
    port map (
            O => \N__59717\,
            I => \N__59677\
        );

    \I__14322\ : InMux
    port map (
            O => \N__59716\,
            I => \N__59677\
        );

    \I__14321\ : InMux
    port map (
            O => \N__59715\,
            I => \N__59654\
        );

    \I__14320\ : InMux
    port map (
            O => \N__59714\,
            I => \N__59654\
        );

    \I__14319\ : InMux
    port map (
            O => \N__59713\,
            I => \N__59654\
        );

    \I__14318\ : InMux
    port map (
            O => \N__59712\,
            I => \N__59654\
        );

    \I__14317\ : InMux
    port map (
            O => \N__59711\,
            I => \N__59654\
        );

    \I__14316\ : InMux
    port map (
            O => \N__59710\,
            I => \N__59654\
        );

    \I__14315\ : InMux
    port map (
            O => \N__59709\,
            I => \N__59654\
        );

    \I__14314\ : InMux
    port map (
            O => \N__59708\,
            I => \N__59654\
        );

    \I__14313\ : InMux
    port map (
            O => \N__59707\,
            I => \N__59625\
        );

    \I__14312\ : InMux
    port map (
            O => \N__59706\,
            I => \N__59625\
        );

    \I__14311\ : InMux
    port map (
            O => \N__59705\,
            I => \N__59625\
        );

    \I__14310\ : InMux
    port map (
            O => \N__59704\,
            I => \N__59608\
        );

    \I__14309\ : InMux
    port map (
            O => \N__59703\,
            I => \N__59608\
        );

    \I__14308\ : InMux
    port map (
            O => \N__59702\,
            I => \N__59608\
        );

    \I__14307\ : InMux
    port map (
            O => \N__59699\,
            I => \N__59608\
        );

    \I__14306\ : InMux
    port map (
            O => \N__59698\,
            I => \N__59608\
        );

    \I__14305\ : InMux
    port map (
            O => \N__59697\,
            I => \N__59608\
        );

    \I__14304\ : InMux
    port map (
            O => \N__59696\,
            I => \N__59608\
        );

    \I__14303\ : InMux
    port map (
            O => \N__59695\,
            I => \N__59608\
        );

    \I__14302\ : LocalMux
    port map (
            O => \N__59690\,
            I => \N__59582\
        );

    \I__14301\ : LocalMux
    port map (
            O => \N__59677\,
            I => \N__59582\
        );

    \I__14300\ : InMux
    port map (
            O => \N__59676\,
            I => \N__59569\
        );

    \I__14299\ : InMux
    port map (
            O => \N__59675\,
            I => \N__59569\
        );

    \I__14298\ : InMux
    port map (
            O => \N__59674\,
            I => \N__59569\
        );

    \I__14297\ : InMux
    port map (
            O => \N__59673\,
            I => \N__59569\
        );

    \I__14296\ : InMux
    port map (
            O => \N__59672\,
            I => \N__59569\
        );

    \I__14295\ : InMux
    port map (
            O => \N__59671\,
            I => \N__59569\
        );

    \I__14294\ : LocalMux
    port map (
            O => \N__59654\,
            I => \N__59566\
        );

    \I__14293\ : InMux
    port map (
            O => \N__59653\,
            I => \N__59559\
        );

    \I__14292\ : InMux
    port map (
            O => \N__59652\,
            I => \N__59559\
        );

    \I__14291\ : InMux
    port map (
            O => \N__59651\,
            I => \N__59559\
        );

    \I__14290\ : InMux
    port map (
            O => \N__59650\,
            I => \N__59524\
        );

    \I__14289\ : InMux
    port map (
            O => \N__59649\,
            I => \N__59524\
        );

    \I__14288\ : InMux
    port map (
            O => \N__59648\,
            I => \N__59524\
        );

    \I__14287\ : InMux
    port map (
            O => \N__59647\,
            I => \N__59524\
        );

    \I__14286\ : InMux
    port map (
            O => \N__59646\,
            I => \N__59524\
        );

    \I__14285\ : InMux
    port map (
            O => \N__59645\,
            I => \N__59524\
        );

    \I__14284\ : InMux
    port map (
            O => \N__59644\,
            I => \N__59524\
        );

    \I__14283\ : InMux
    port map (
            O => \N__59643\,
            I => \N__59524\
        );

    \I__14282\ : InMux
    port map (
            O => \N__59642\,
            I => \N__59517\
        );

    \I__14281\ : InMux
    port map (
            O => \N__59641\,
            I => \N__59517\
        );

    \I__14280\ : InMux
    port map (
            O => \N__59640\,
            I => \N__59517\
        );

    \I__14279\ : InMux
    port map (
            O => \N__59639\,
            I => \N__59487\
        );

    \I__14278\ : InMux
    port map (
            O => \N__59638\,
            I => \N__59487\
        );

    \I__14277\ : InMux
    port map (
            O => \N__59637\,
            I => \N__59487\
        );

    \I__14276\ : InMux
    port map (
            O => \N__59636\,
            I => \N__59487\
        );

    \I__14275\ : InMux
    port map (
            O => \N__59635\,
            I => \N__59487\
        );

    \I__14274\ : InMux
    port map (
            O => \N__59634\,
            I => \N__59487\
        );

    \I__14273\ : InMux
    port map (
            O => \N__59633\,
            I => \N__59487\
        );

    \I__14272\ : InMux
    port map (
            O => \N__59632\,
            I => \N__59487\
        );

    \I__14271\ : LocalMux
    port map (
            O => \N__59625\,
            I => \N__59482\
        );

    \I__14270\ : LocalMux
    port map (
            O => \N__59608\,
            I => \N__59482\
        );

    \I__14269\ : InMux
    port map (
            O => \N__59607\,
            I => \N__59465\
        );

    \I__14268\ : InMux
    port map (
            O => \N__59606\,
            I => \N__59465\
        );

    \I__14267\ : InMux
    port map (
            O => \N__59605\,
            I => \N__59465\
        );

    \I__14266\ : InMux
    port map (
            O => \N__59604\,
            I => \N__59465\
        );

    \I__14265\ : InMux
    port map (
            O => \N__59603\,
            I => \N__59465\
        );

    \I__14264\ : InMux
    port map (
            O => \N__59602\,
            I => \N__59465\
        );

    \I__14263\ : InMux
    port map (
            O => \N__59601\,
            I => \N__59465\
        );

    \I__14262\ : InMux
    port map (
            O => \N__59600\,
            I => \N__59465\
        );

    \I__14261\ : InMux
    port map (
            O => \N__59599\,
            I => \N__59460\
        );

    \I__14260\ : InMux
    port map (
            O => \N__59598\,
            I => \N__59460\
        );

    \I__14259\ : InMux
    port map (
            O => \N__59597\,
            I => \N__59449\
        );

    \I__14258\ : InMux
    port map (
            O => \N__59596\,
            I => \N__59449\
        );

    \I__14257\ : InMux
    port map (
            O => \N__59595\,
            I => \N__59449\
        );

    \I__14256\ : InMux
    port map (
            O => \N__59594\,
            I => \N__59449\
        );

    \I__14255\ : InMux
    port map (
            O => \N__59593\,
            I => \N__59449\
        );

    \I__14254\ : InMux
    port map (
            O => \N__59592\,
            I => \N__59399\
        );

    \I__14253\ : InMux
    port map (
            O => \N__59591\,
            I => \N__59399\
        );

    \I__14252\ : InMux
    port map (
            O => \N__59590\,
            I => \N__59399\
        );

    \I__14251\ : InMux
    port map (
            O => \N__59589\,
            I => \N__59399\
        );

    \I__14250\ : InMux
    port map (
            O => \N__59588\,
            I => \N__59399\
        );

    \I__14249\ : InMux
    port map (
            O => \N__59587\,
            I => \N__59399\
        );

    \I__14248\ : Span4Mux_v
    port map (
            O => \N__59582\,
            I => \N__59394\
        );

    \I__14247\ : LocalMux
    port map (
            O => \N__59569\,
            I => \N__59394\
        );

    \I__14246\ : Span4Mux_h
    port map (
            O => \N__59566\,
            I => \N__59389\
        );

    \I__14245\ : LocalMux
    port map (
            O => \N__59559\,
            I => \N__59389\
        );

    \I__14244\ : InMux
    port map (
            O => \N__59558\,
            I => \N__59374\
        );

    \I__14243\ : InMux
    port map (
            O => \N__59557\,
            I => \N__59374\
        );

    \I__14242\ : InMux
    port map (
            O => \N__59556\,
            I => \N__59374\
        );

    \I__14241\ : InMux
    port map (
            O => \N__59555\,
            I => \N__59371\
        );

    \I__14240\ : InMux
    port map (
            O => \N__59554\,
            I => \N__59368\
        );

    \I__14239\ : InMux
    port map (
            O => \N__59553\,
            I => \N__59365\
        );

    \I__14238\ : InMux
    port map (
            O => \N__59552\,
            I => \N__59348\
        );

    \I__14237\ : InMux
    port map (
            O => \N__59551\,
            I => \N__59348\
        );

    \I__14236\ : InMux
    port map (
            O => \N__59550\,
            I => \N__59348\
        );

    \I__14235\ : InMux
    port map (
            O => \N__59549\,
            I => \N__59348\
        );

    \I__14234\ : InMux
    port map (
            O => \N__59548\,
            I => \N__59348\
        );

    \I__14233\ : InMux
    port map (
            O => \N__59547\,
            I => \N__59348\
        );

    \I__14232\ : InMux
    port map (
            O => \N__59546\,
            I => \N__59348\
        );

    \I__14231\ : InMux
    port map (
            O => \N__59545\,
            I => \N__59348\
        );

    \I__14230\ : CascadeMux
    port map (
            O => \N__59544\,
            I => \N__59345\
        );

    \I__14229\ : CascadeMux
    port map (
            O => \N__59543\,
            I => \N__59342\
        );

    \I__14228\ : CascadeMux
    port map (
            O => \N__59542\,
            I => \N__59339\
        );

    \I__14227\ : CascadeMux
    port map (
            O => \N__59541\,
            I => \N__59336\
        );

    \I__14226\ : LocalMux
    port map (
            O => \N__59524\,
            I => \N__59328\
        );

    \I__14225\ : LocalMux
    port map (
            O => \N__59517\,
            I => \N__59328\
        );

    \I__14224\ : InMux
    port map (
            O => \N__59516\,
            I => \N__59311\
        );

    \I__14223\ : InMux
    port map (
            O => \N__59515\,
            I => \N__59311\
        );

    \I__14222\ : InMux
    port map (
            O => \N__59514\,
            I => \N__59311\
        );

    \I__14221\ : InMux
    port map (
            O => \N__59513\,
            I => \N__59311\
        );

    \I__14220\ : InMux
    port map (
            O => \N__59512\,
            I => \N__59311\
        );

    \I__14219\ : InMux
    port map (
            O => \N__59511\,
            I => \N__59311\
        );

    \I__14218\ : InMux
    port map (
            O => \N__59510\,
            I => \N__59311\
        );

    \I__14217\ : InMux
    port map (
            O => \N__59509\,
            I => \N__59311\
        );

    \I__14216\ : InMux
    port map (
            O => \N__59508\,
            I => \N__59308\
        );

    \I__14215\ : InMux
    port map (
            O => \N__59507\,
            I => \N__59299\
        );

    \I__14214\ : InMux
    port map (
            O => \N__59506\,
            I => \N__59299\
        );

    \I__14213\ : InMux
    port map (
            O => \N__59505\,
            I => \N__59299\
        );

    \I__14212\ : InMux
    port map (
            O => \N__59504\,
            I => \N__59299\
        );

    \I__14211\ : LocalMux
    port map (
            O => \N__59487\,
            I => \N__59294\
        );

    \I__14210\ : Span4Mux_v
    port map (
            O => \N__59482\,
            I => \N__59294\
        );

    \I__14209\ : LocalMux
    port map (
            O => \N__59465\,
            I => \N__59287\
        );

    \I__14208\ : LocalMux
    port map (
            O => \N__59460\,
            I => \N__59287\
        );

    \I__14207\ : LocalMux
    port map (
            O => \N__59449\,
            I => \N__59287\
        );

    \I__14206\ : CascadeMux
    port map (
            O => \N__59448\,
            I => \N__59284\
        );

    \I__14205\ : CascadeMux
    port map (
            O => \N__59447\,
            I => \N__59281\
        );

    \I__14204\ : CascadeMux
    port map (
            O => \N__59446\,
            I => \N__59278\
        );

    \I__14203\ : CascadeMux
    port map (
            O => \N__59445\,
            I => \N__59272\
        );

    \I__14202\ : InMux
    port map (
            O => \N__59444\,
            I => \N__59269\
        );

    \I__14201\ : InMux
    port map (
            O => \N__59443\,
            I => \N__59262\
        );

    \I__14200\ : InMux
    port map (
            O => \N__59442\,
            I => \N__59262\
        );

    \I__14199\ : InMux
    port map (
            O => \N__59441\,
            I => \N__59262\
        );

    \I__14198\ : InMux
    port map (
            O => \N__59440\,
            I => \N__59245\
        );

    \I__14197\ : InMux
    port map (
            O => \N__59439\,
            I => \N__59245\
        );

    \I__14196\ : InMux
    port map (
            O => \N__59438\,
            I => \N__59245\
        );

    \I__14195\ : InMux
    port map (
            O => \N__59437\,
            I => \N__59245\
        );

    \I__14194\ : InMux
    port map (
            O => \N__59436\,
            I => \N__59245\
        );

    \I__14193\ : InMux
    port map (
            O => \N__59435\,
            I => \N__59245\
        );

    \I__14192\ : InMux
    port map (
            O => \N__59434\,
            I => \N__59245\
        );

    \I__14191\ : InMux
    port map (
            O => \N__59433\,
            I => \N__59245\
        );

    \I__14190\ : InMux
    port map (
            O => \N__59432\,
            I => \N__59240\
        );

    \I__14189\ : InMux
    port map (
            O => \N__59431\,
            I => \N__59240\
        );

    \I__14188\ : InMux
    port map (
            O => \N__59430\,
            I => \N__59223\
        );

    \I__14187\ : InMux
    port map (
            O => \N__59429\,
            I => \N__59223\
        );

    \I__14186\ : InMux
    port map (
            O => \N__59428\,
            I => \N__59223\
        );

    \I__14185\ : InMux
    port map (
            O => \N__59427\,
            I => \N__59223\
        );

    \I__14184\ : InMux
    port map (
            O => \N__59426\,
            I => \N__59223\
        );

    \I__14183\ : InMux
    port map (
            O => \N__59425\,
            I => \N__59223\
        );

    \I__14182\ : InMux
    port map (
            O => \N__59424\,
            I => \N__59223\
        );

    \I__14181\ : InMux
    port map (
            O => \N__59423\,
            I => \N__59223\
        );

    \I__14180\ : InMux
    port map (
            O => \N__59422\,
            I => \N__59216\
        );

    \I__14179\ : InMux
    port map (
            O => \N__59421\,
            I => \N__59216\
        );

    \I__14178\ : InMux
    port map (
            O => \N__59420\,
            I => \N__59216\
        );

    \I__14177\ : InMux
    port map (
            O => \N__59419\,
            I => \N__59199\
        );

    \I__14176\ : InMux
    port map (
            O => \N__59418\,
            I => \N__59199\
        );

    \I__14175\ : InMux
    port map (
            O => \N__59417\,
            I => \N__59199\
        );

    \I__14174\ : InMux
    port map (
            O => \N__59416\,
            I => \N__59199\
        );

    \I__14173\ : InMux
    port map (
            O => \N__59415\,
            I => \N__59199\
        );

    \I__14172\ : InMux
    port map (
            O => \N__59414\,
            I => \N__59199\
        );

    \I__14171\ : InMux
    port map (
            O => \N__59413\,
            I => \N__59199\
        );

    \I__14170\ : InMux
    port map (
            O => \N__59412\,
            I => \N__59199\
        );

    \I__14169\ : LocalMux
    port map (
            O => \N__59399\,
            I => \N__59194\
        );

    \I__14168\ : Span4Mux_h
    port map (
            O => \N__59394\,
            I => \N__59194\
        );

    \I__14167\ : Span4Mux_v
    port map (
            O => \N__59389\,
            I => \N__59191\
        );

    \I__14166\ : InMux
    port map (
            O => \N__59388\,
            I => \N__59180\
        );

    \I__14165\ : InMux
    port map (
            O => \N__59387\,
            I => \N__59171\
        );

    \I__14164\ : InMux
    port map (
            O => \N__59386\,
            I => \N__59171\
        );

    \I__14163\ : InMux
    port map (
            O => \N__59385\,
            I => \N__59171\
        );

    \I__14162\ : InMux
    port map (
            O => \N__59384\,
            I => \N__59171\
        );

    \I__14161\ : InMux
    port map (
            O => \N__59383\,
            I => \N__59166\
        );

    \I__14160\ : InMux
    port map (
            O => \N__59382\,
            I => \N__59166\
        );

    \I__14159\ : InMux
    port map (
            O => \N__59381\,
            I => \N__59157\
        );

    \I__14158\ : LocalMux
    port map (
            O => \N__59374\,
            I => \N__59150\
        );

    \I__14157\ : LocalMux
    port map (
            O => \N__59371\,
            I => \N__59150\
        );

    \I__14156\ : LocalMux
    port map (
            O => \N__59368\,
            I => \N__59150\
        );

    \I__14155\ : LocalMux
    port map (
            O => \N__59365\,
            I => \N__59134\
        );

    \I__14154\ : LocalMux
    port map (
            O => \N__59348\,
            I => \N__59134\
        );

    \I__14153\ : InMux
    port map (
            O => \N__59345\,
            I => \N__59119\
        );

    \I__14152\ : InMux
    port map (
            O => \N__59342\,
            I => \N__59119\
        );

    \I__14151\ : InMux
    port map (
            O => \N__59339\,
            I => \N__59119\
        );

    \I__14150\ : InMux
    port map (
            O => \N__59336\,
            I => \N__59119\
        );

    \I__14149\ : InMux
    port map (
            O => \N__59335\,
            I => \N__59119\
        );

    \I__14148\ : InMux
    port map (
            O => \N__59334\,
            I => \N__59119\
        );

    \I__14147\ : InMux
    port map (
            O => \N__59333\,
            I => \N__59119\
        );

    \I__14146\ : Span4Mux_v
    port map (
            O => \N__59328\,
            I => \N__59106\
        );

    \I__14145\ : LocalMux
    port map (
            O => \N__59311\,
            I => \N__59106\
        );

    \I__14144\ : LocalMux
    port map (
            O => \N__59308\,
            I => \N__59106\
        );

    \I__14143\ : LocalMux
    port map (
            O => \N__59299\,
            I => \N__59106\
        );

    \I__14142\ : Span4Mux_h
    port map (
            O => \N__59294\,
            I => \N__59106\
        );

    \I__14141\ : Span4Mux_v
    port map (
            O => \N__59287\,
            I => \N__59106\
        );

    \I__14140\ : InMux
    port map (
            O => \N__59284\,
            I => \N__59093\
        );

    \I__14139\ : InMux
    port map (
            O => \N__59281\,
            I => \N__59093\
        );

    \I__14138\ : InMux
    port map (
            O => \N__59278\,
            I => \N__59093\
        );

    \I__14137\ : InMux
    port map (
            O => \N__59277\,
            I => \N__59093\
        );

    \I__14136\ : InMux
    port map (
            O => \N__59276\,
            I => \N__59093\
        );

    \I__14135\ : InMux
    port map (
            O => \N__59275\,
            I => \N__59093\
        );

    \I__14134\ : InMux
    port map (
            O => \N__59272\,
            I => \N__59090\
        );

    \I__14133\ : LocalMux
    port map (
            O => \N__59269\,
            I => \N__59085\
        );

    \I__14132\ : LocalMux
    port map (
            O => \N__59262\,
            I => \N__59085\
        );

    \I__14131\ : LocalMux
    port map (
            O => \N__59245\,
            I => \N__59082\
        );

    \I__14130\ : LocalMux
    port map (
            O => \N__59240\,
            I => \N__59071\
        );

    \I__14129\ : LocalMux
    port map (
            O => \N__59223\,
            I => \N__59071\
        );

    \I__14128\ : LocalMux
    port map (
            O => \N__59216\,
            I => \N__59071\
        );

    \I__14127\ : LocalMux
    port map (
            O => \N__59199\,
            I => \N__59071\
        );

    \I__14126\ : Span4Mux_v
    port map (
            O => \N__59194\,
            I => \N__59071\
        );

    \I__14125\ : Span4Mux_v
    port map (
            O => \N__59191\,
            I => \N__59068\
        );

    \I__14124\ : InMux
    port map (
            O => \N__59190\,
            I => \N__59051\
        );

    \I__14123\ : InMux
    port map (
            O => \N__59189\,
            I => \N__59051\
        );

    \I__14122\ : InMux
    port map (
            O => \N__59188\,
            I => \N__59051\
        );

    \I__14121\ : InMux
    port map (
            O => \N__59187\,
            I => \N__59051\
        );

    \I__14120\ : InMux
    port map (
            O => \N__59186\,
            I => \N__59051\
        );

    \I__14119\ : InMux
    port map (
            O => \N__59185\,
            I => \N__59051\
        );

    \I__14118\ : InMux
    port map (
            O => \N__59184\,
            I => \N__59051\
        );

    \I__14117\ : InMux
    port map (
            O => \N__59183\,
            I => \N__59051\
        );

    \I__14116\ : LocalMux
    port map (
            O => \N__59180\,
            I => \N__59046\
        );

    \I__14115\ : LocalMux
    port map (
            O => \N__59171\,
            I => \N__59046\
        );

    \I__14114\ : LocalMux
    port map (
            O => \N__59166\,
            I => \N__59043\
        );

    \I__14113\ : InMux
    port map (
            O => \N__59165\,
            I => \N__59038\
        );

    \I__14112\ : InMux
    port map (
            O => \N__59164\,
            I => \N__59038\
        );

    \I__14111\ : CascadeMux
    port map (
            O => \N__59163\,
            I => \N__59035\
        );

    \I__14110\ : CascadeMux
    port map (
            O => \N__59162\,
            I => \N__59032\
        );

    \I__14109\ : CascadeMux
    port map (
            O => \N__59161\,
            I => \N__59029\
        );

    \I__14108\ : CascadeMux
    port map (
            O => \N__59160\,
            I => \N__59026\
        );

    \I__14107\ : LocalMux
    port map (
            O => \N__59157\,
            I => \N__59020\
        );

    \I__14106\ : Span4Mux_v
    port map (
            O => \N__59150\,
            I => \N__59017\
        );

    \I__14105\ : InMux
    port map (
            O => \N__59149\,
            I => \N__58993\
        );

    \I__14104\ : InMux
    port map (
            O => \N__59148\,
            I => \N__58993\
        );

    \I__14103\ : InMux
    port map (
            O => \N__59147\,
            I => \N__58993\
        );

    \I__14102\ : InMux
    port map (
            O => \N__59146\,
            I => \N__58993\
        );

    \I__14101\ : InMux
    port map (
            O => \N__59145\,
            I => \N__58993\
        );

    \I__14100\ : InMux
    port map (
            O => \N__59144\,
            I => \N__58993\
        );

    \I__14099\ : InMux
    port map (
            O => \N__59143\,
            I => \N__58993\
        );

    \I__14098\ : InMux
    port map (
            O => \N__59142\,
            I => \N__58993\
        );

    \I__14097\ : InMux
    port map (
            O => \N__59141\,
            I => \N__58988\
        );

    \I__14096\ : InMux
    port map (
            O => \N__59140\,
            I => \N__58988\
        );

    \I__14095\ : InMux
    port map (
            O => \N__59139\,
            I => \N__58985\
        );

    \I__14094\ : Span4Mux_v
    port map (
            O => \N__59134\,
            I => \N__58978\
        );

    \I__14093\ : LocalMux
    port map (
            O => \N__59119\,
            I => \N__58978\
        );

    \I__14092\ : Span4Mux_h
    port map (
            O => \N__59106\,
            I => \N__58978\
        );

    \I__14091\ : LocalMux
    port map (
            O => \N__59093\,
            I => \N__58971\
        );

    \I__14090\ : LocalMux
    port map (
            O => \N__59090\,
            I => \N__58971\
        );

    \I__14089\ : Span4Mux_v
    port map (
            O => \N__59085\,
            I => \N__58971\
        );

    \I__14088\ : Span4Mux_v
    port map (
            O => \N__59082\,
            I => \N__58964\
        );

    \I__14087\ : Span4Mux_v
    port map (
            O => \N__59071\,
            I => \N__58964\
        );

    \I__14086\ : Span4Mux_h
    port map (
            O => \N__59068\,
            I => \N__58964\
        );

    \I__14085\ : LocalMux
    port map (
            O => \N__59051\,
            I => \N__58955\
        );

    \I__14084\ : Span4Mux_v
    port map (
            O => \N__59046\,
            I => \N__58955\
        );

    \I__14083\ : Span4Mux_h
    port map (
            O => \N__59043\,
            I => \N__58955\
        );

    \I__14082\ : LocalMux
    port map (
            O => \N__59038\,
            I => \N__58955\
        );

    \I__14081\ : InMux
    port map (
            O => \N__59035\,
            I => \N__58940\
        );

    \I__14080\ : InMux
    port map (
            O => \N__59032\,
            I => \N__58940\
        );

    \I__14079\ : InMux
    port map (
            O => \N__59029\,
            I => \N__58940\
        );

    \I__14078\ : InMux
    port map (
            O => \N__59026\,
            I => \N__58940\
        );

    \I__14077\ : InMux
    port map (
            O => \N__59025\,
            I => \N__58940\
        );

    \I__14076\ : InMux
    port map (
            O => \N__59024\,
            I => \N__58940\
        );

    \I__14075\ : InMux
    port map (
            O => \N__59023\,
            I => \N__58940\
        );

    \I__14074\ : Span4Mux_v
    port map (
            O => \N__59020\,
            I => \N__58935\
        );

    \I__14073\ : Span4Mux_v
    port map (
            O => \N__59017\,
            I => \N__58935\
        );

    \I__14072\ : InMux
    port map (
            O => \N__59016\,
            I => \N__58926\
        );

    \I__14071\ : InMux
    port map (
            O => \N__59015\,
            I => \N__58926\
        );

    \I__14070\ : InMux
    port map (
            O => \N__59014\,
            I => \N__58926\
        );

    \I__14069\ : InMux
    port map (
            O => \N__59013\,
            I => \N__58926\
        );

    \I__14068\ : InMux
    port map (
            O => \N__59012\,
            I => \N__58919\
        );

    \I__14067\ : InMux
    port map (
            O => \N__59011\,
            I => \N__58919\
        );

    \I__14066\ : InMux
    port map (
            O => \N__59010\,
            I => \N__58919\
        );

    \I__14065\ : LocalMux
    port map (
            O => \N__58993\,
            I => \N__58916\
        );

    \I__14064\ : LocalMux
    port map (
            O => \N__58988\,
            I => \N__58909\
        );

    \I__14063\ : LocalMux
    port map (
            O => \N__58985\,
            I => \N__58909\
        );

    \I__14062\ : Span4Mux_h
    port map (
            O => \N__58978\,
            I => \N__58909\
        );

    \I__14061\ : Span4Mux_v
    port map (
            O => \N__58971\,
            I => \N__58902\
        );

    \I__14060\ : Span4Mux_h
    port map (
            O => \N__58964\,
            I => \N__58902\
        );

    \I__14059\ : Span4Mux_v
    port map (
            O => \N__58955\,
            I => \N__58902\
        );

    \I__14058\ : LocalMux
    port map (
            O => \N__58940\,
            I => \N__58897\
        );

    \I__14057\ : Span4Mux_h
    port map (
            O => \N__58935\,
            I => \N__58897\
        );

    \I__14056\ : LocalMux
    port map (
            O => \N__58926\,
            I => \N_1592_0\
        );

    \I__14055\ : LocalMux
    port map (
            O => \N__58919\,
            I => \N_1592_0\
        );

    \I__14054\ : Odrv12
    port map (
            O => \N__58916\,
            I => \N_1592_0\
        );

    \I__14053\ : Odrv4
    port map (
            O => \N__58909\,
            I => \N_1592_0\
        );

    \I__14052\ : Odrv4
    port map (
            O => \N__58902\,
            I => \N_1592_0\
        );

    \I__14051\ : Odrv4
    port map (
            O => \N__58897\,
            I => \N_1592_0\
        );

    \I__14050\ : CEMux
    port map (
            O => \N__58884\,
            I => \N__58881\
        );

    \I__14049\ : LocalMux
    port map (
            O => \N__58881\,
            I => \N__58876\
        );

    \I__14048\ : CEMux
    port map (
            O => \N__58880\,
            I => \N__58873\
        );

    \I__14047\ : CEMux
    port map (
            O => \N__58879\,
            I => \N__58870\
        );

    \I__14046\ : Span4Mux_h
    port map (
            O => \N__58876\,
            I => \N__58862\
        );

    \I__14045\ : LocalMux
    port map (
            O => \N__58873\,
            I => \N__58862\
        );

    \I__14044\ : LocalMux
    port map (
            O => \N__58870\,
            I => \N__58859\
        );

    \I__14043\ : CEMux
    port map (
            O => \N__58869\,
            I => \N__58856\
        );

    \I__14042\ : CEMux
    port map (
            O => \N__58868\,
            I => \N__58853\
        );

    \I__14041\ : CEMux
    port map (
            O => \N__58867\,
            I => \N__58850\
        );

    \I__14040\ : Span4Mux_h
    port map (
            O => \N__58862\,
            I => \N__58843\
        );

    \I__14039\ : Span4Mux_h
    port map (
            O => \N__58859\,
            I => \N__58843\
        );

    \I__14038\ : LocalMux
    port map (
            O => \N__58856\,
            I => \N__58843\
        );

    \I__14037\ : LocalMux
    port map (
            O => \N__58853\,
            I => \N__58840\
        );

    \I__14036\ : LocalMux
    port map (
            O => \N__58850\,
            I => \N__58837\
        );

    \I__14035\ : Span4Mux_v
    port map (
            O => \N__58843\,
            I => \N__58834\
        );

    \I__14034\ : Span12Mux_v
    port map (
            O => \N__58840\,
            I => \N__58831\
        );

    \I__14033\ : Span4Mux_v
    port map (
            O => \N__58837\,
            I => \N__58828\
        );

    \I__14032\ : Span4Mux_h
    port map (
            O => \N__58834\,
            I => \N__58825\
        );

    \I__14031\ : Odrv12
    port map (
            O => \N__58831\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0\
        );

    \I__14030\ : Odrv4
    port map (
            O => \N__58828\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0\
        );

    \I__14029\ : Odrv4
    port map (
            O => \N__58825\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0\
        );

    \I__14028\ : InMux
    port map (
            O => \N__58818\,
            I => \N__58815\
        );

    \I__14027\ : LocalMux
    port map (
            O => \N__58815\,
            I => \N__58812\
        );

    \I__14026\ : Span4Mux_v
    port map (
            O => \N__58812\,
            I => \N__58809\
        );

    \I__14025\ : Span4Mux_h
    port map (
            O => \N__58809\,
            I => \N__58806\
        );

    \I__14024\ : Sp12to4
    port map (
            O => \N__58806\,
            I => \N__58803\
        );

    \I__14023\ : Span12Mux_h
    port map (
            O => \N__58803\,
            I => \N__58800\
        );

    \I__14022\ : Odrv12
    port map (
            O => \N__58800\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_9\
        );

    \I__14021\ : InMux
    port map (
            O => \N__58797\,
            I => \N__58792\
        );

    \I__14020\ : InMux
    port map (
            O => \N__58796\,
            I => \N__58789\
        );

    \I__14019\ : InMux
    port map (
            O => \N__58795\,
            I => \N__58784\
        );

    \I__14018\ : LocalMux
    port map (
            O => \N__58792\,
            I => \N__58780\
        );

    \I__14017\ : LocalMux
    port map (
            O => \N__58789\,
            I => \N__58776\
        );

    \I__14016\ : InMux
    port map (
            O => \N__58788\,
            I => \N__58773\
        );

    \I__14015\ : InMux
    port map (
            O => \N__58787\,
            I => \N__58770\
        );

    \I__14014\ : LocalMux
    port map (
            O => \N__58784\,
            I => \N__58767\
        );

    \I__14013\ : InMux
    port map (
            O => \N__58783\,
            I => \N__58763\
        );

    \I__14012\ : Span4Mux_h
    port map (
            O => \N__58780\,
            I => \N__58760\
        );

    \I__14011\ : InMux
    port map (
            O => \N__58779\,
            I => \N__58757\
        );

    \I__14010\ : Span4Mux_h
    port map (
            O => \N__58776\,
            I => \N__58750\
        );

    \I__14009\ : LocalMux
    port map (
            O => \N__58773\,
            I => \N__58750\
        );

    \I__14008\ : LocalMux
    port map (
            O => \N__58770\,
            I => \N__58750\
        );

    \I__14007\ : Span4Mux_v
    port map (
            O => \N__58767\,
            I => \N__58746\
        );

    \I__14006\ : CascadeMux
    port map (
            O => \N__58766\,
            I => \N__58743\
        );

    \I__14005\ : LocalMux
    port map (
            O => \N__58763\,
            I => \N__58738\
        );

    \I__14004\ : Span4Mux_h
    port map (
            O => \N__58760\,
            I => \N__58738\
        );

    \I__14003\ : LocalMux
    port map (
            O => \N__58757\,
            I => \N__58733\
        );

    \I__14002\ : Sp12to4
    port map (
            O => \N__58750\,
            I => \N__58733\
        );

    \I__14001\ : InMux
    port map (
            O => \N__58749\,
            I => \N__58730\
        );

    \I__14000\ : Sp12to4
    port map (
            O => \N__58746\,
            I => \N__58727\
        );

    \I__13999\ : InMux
    port map (
            O => \N__58743\,
            I => \N__58724\
        );

    \I__13998\ : Span4Mux_v
    port map (
            O => \N__58738\,
            I => \N__58721\
        );

    \I__13997\ : Span12Mux_v
    port map (
            O => \N__58733\,
            I => \N__58716\
        );

    \I__13996\ : LocalMux
    port map (
            O => \N__58730\,
            I => \N__58716\
        );

    \I__13995\ : Odrv12
    port map (
            O => \N__58727\,
            I => \I2C_top_level_inst1_s_data_oreg_10\
        );

    \I__13994\ : LocalMux
    port map (
            O => \N__58724\,
            I => \I2C_top_level_inst1_s_data_oreg_10\
        );

    \I__13993\ : Odrv4
    port map (
            O => \N__58721\,
            I => \I2C_top_level_inst1_s_data_oreg_10\
        );

    \I__13992\ : Odrv12
    port map (
            O => \N__58716\,
            I => \I2C_top_level_inst1_s_data_oreg_10\
        );

    \I__13991\ : InMux
    port map (
            O => \N__58707\,
            I => \N__58704\
        );

    \I__13990\ : LocalMux
    port map (
            O => \N__58704\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_10\
        );

    \I__13989\ : InMux
    port map (
            O => \N__58701\,
            I => \N__58697\
        );

    \I__13988\ : InMux
    port map (
            O => \N__58700\,
            I => \N__58693\
        );

    \I__13987\ : LocalMux
    port map (
            O => \N__58697\,
            I => \N__58688\
        );

    \I__13986\ : InMux
    port map (
            O => \N__58696\,
            I => \N__58685\
        );

    \I__13985\ : LocalMux
    port map (
            O => \N__58693\,
            I => \N__58681\
        );

    \I__13984\ : InMux
    port map (
            O => \N__58692\,
            I => \N__58678\
        );

    \I__13983\ : InMux
    port map (
            O => \N__58691\,
            I => \N__58675\
        );

    \I__13982\ : Span4Mux_v
    port map (
            O => \N__58688\,
            I => \N__58670\
        );

    \I__13981\ : LocalMux
    port map (
            O => \N__58685\,
            I => \N__58670\
        );

    \I__13980\ : InMux
    port map (
            O => \N__58684\,
            I => \N__58667\
        );

    \I__13979\ : Span4Mux_h
    port map (
            O => \N__58681\,
            I => \N__58661\
        );

    \I__13978\ : LocalMux
    port map (
            O => \N__58678\,
            I => \N__58661\
        );

    \I__13977\ : LocalMux
    port map (
            O => \N__58675\,
            I => \N__58657\
        );

    \I__13976\ : Span4Mux_h
    port map (
            O => \N__58670\,
            I => \N__58652\
        );

    \I__13975\ : LocalMux
    port map (
            O => \N__58667\,
            I => \N__58652\
        );

    \I__13974\ : InMux
    port map (
            O => \N__58666\,
            I => \N__58649\
        );

    \I__13973\ : Span4Mux_v
    port map (
            O => \N__58661\,
            I => \N__58646\
        );

    \I__13972\ : InMux
    port map (
            O => \N__58660\,
            I => \N__58643\
        );

    \I__13971\ : Span4Mux_v
    port map (
            O => \N__58657\,
            I => \N__58638\
        );

    \I__13970\ : Span4Mux_v
    port map (
            O => \N__58652\,
            I => \N__58638\
        );

    \I__13969\ : LocalMux
    port map (
            O => \N__58649\,
            I => \N__58635\
        );

    \I__13968\ : Span4Mux_h
    port map (
            O => \N__58646\,
            I => \N__58629\
        );

    \I__13967\ : LocalMux
    port map (
            O => \N__58643\,
            I => \N__58629\
        );

    \I__13966\ : Sp12to4
    port map (
            O => \N__58638\,
            I => \N__58626\
        );

    \I__13965\ : Span4Mux_v
    port map (
            O => \N__58635\,
            I => \N__58623\
        );

    \I__13964\ : CascadeMux
    port map (
            O => \N__58634\,
            I => \N__58620\
        );

    \I__13963\ : Span4Mux_v
    port map (
            O => \N__58629\,
            I => \N__58617\
        );

    \I__13962\ : Span12Mux_h
    port map (
            O => \N__58626\,
            I => \N__58612\
        );

    \I__13961\ : Sp12to4
    port map (
            O => \N__58623\,
            I => \N__58612\
        );

    \I__13960\ : InMux
    port map (
            O => \N__58620\,
            I => \N__58609\
        );

    \I__13959\ : Odrv4
    port map (
            O => \N__58617\,
            I => \I2C_top_level_inst1_s_data_oreg_11\
        );

    \I__13958\ : Odrv12
    port map (
            O => \N__58612\,
            I => \I2C_top_level_inst1_s_data_oreg_11\
        );

    \I__13957\ : LocalMux
    port map (
            O => \N__58609\,
            I => \I2C_top_level_inst1_s_data_oreg_11\
        );

    \I__13956\ : InMux
    port map (
            O => \N__58602\,
            I => \N__58599\
        );

    \I__13955\ : LocalMux
    port map (
            O => \N__58599\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_11\
        );

    \I__13954\ : InMux
    port map (
            O => \N__58596\,
            I => \N__58586\
        );

    \I__13953\ : InMux
    port map (
            O => \N__58595\,
            I => \N__58583\
        );

    \I__13952\ : InMux
    port map (
            O => \N__58594\,
            I => \N__58580\
        );

    \I__13951\ : CascadeMux
    port map (
            O => \N__58593\,
            I => \N__58577\
        );

    \I__13950\ : InMux
    port map (
            O => \N__58592\,
            I => \N__58574\
        );

    \I__13949\ : InMux
    port map (
            O => \N__58591\,
            I => \N__58571\
        );

    \I__13948\ : InMux
    port map (
            O => \N__58590\,
            I => \N__58568\
        );

    \I__13947\ : InMux
    port map (
            O => \N__58589\,
            I => \N__58565\
        );

    \I__13946\ : LocalMux
    port map (
            O => \N__58586\,
            I => \N__58562\
        );

    \I__13945\ : LocalMux
    port map (
            O => \N__58583\,
            I => \N__58556\
        );

    \I__13944\ : LocalMux
    port map (
            O => \N__58580\,
            I => \N__58556\
        );

    \I__13943\ : InMux
    port map (
            O => \N__58577\,
            I => \N__58553\
        );

    \I__13942\ : LocalMux
    port map (
            O => \N__58574\,
            I => \N__58550\
        );

    \I__13941\ : LocalMux
    port map (
            O => \N__58571\,
            I => \N__58545\
        );

    \I__13940\ : LocalMux
    port map (
            O => \N__58568\,
            I => \N__58545\
        );

    \I__13939\ : LocalMux
    port map (
            O => \N__58565\,
            I => \N__58540\
        );

    \I__13938\ : Span4Mux_h
    port map (
            O => \N__58562\,
            I => \N__58540\
        );

    \I__13937\ : InMux
    port map (
            O => \N__58561\,
            I => \N__58537\
        );

    \I__13936\ : Span4Mux_v
    port map (
            O => \N__58556\,
            I => \N__58534\
        );

    \I__13935\ : LocalMux
    port map (
            O => \N__58553\,
            I => \N__58531\
        );

    \I__13934\ : Span4Mux_h
    port map (
            O => \N__58550\,
            I => \N__58524\
        );

    \I__13933\ : Span4Mux_v
    port map (
            O => \N__58545\,
            I => \N__58524\
        );

    \I__13932\ : Span4Mux_v
    port map (
            O => \N__58540\,
            I => \N__58524\
        );

    \I__13931\ : LocalMux
    port map (
            O => \N__58537\,
            I => \N__58521\
        );

    \I__13930\ : Span4Mux_h
    port map (
            O => \N__58534\,
            I => \N__58518\
        );

    \I__13929\ : Span4Mux_v
    port map (
            O => \N__58531\,
            I => \N__58515\
        );

    \I__13928\ : Span4Mux_h
    port map (
            O => \N__58524\,
            I => \N__58512\
        );

    \I__13927\ : Span12Mux_s8_v
    port map (
            O => \N__58521\,
            I => \N__58509\
        );

    \I__13926\ : Odrv4
    port map (
            O => \N__58518\,
            I => \I2C_top_level_inst1_s_data_oreg_12\
        );

    \I__13925\ : Odrv4
    port map (
            O => \N__58515\,
            I => \I2C_top_level_inst1_s_data_oreg_12\
        );

    \I__13924\ : Odrv4
    port map (
            O => \N__58512\,
            I => \I2C_top_level_inst1_s_data_oreg_12\
        );

    \I__13923\ : Odrv12
    port map (
            O => \N__58509\,
            I => \I2C_top_level_inst1_s_data_oreg_12\
        );

    \I__13922\ : InMux
    port map (
            O => \N__58500\,
            I => \N__58493\
        );

    \I__13921\ : InMux
    port map (
            O => \N__58499\,
            I => \N__58490\
        );

    \I__13920\ : InMux
    port map (
            O => \N__58498\,
            I => \N__58486\
        );

    \I__13919\ : InMux
    port map (
            O => \N__58497\,
            I => \N__58483\
        );

    \I__13918\ : InMux
    port map (
            O => \N__58496\,
            I => \N__58480\
        );

    \I__13917\ : LocalMux
    port map (
            O => \N__58493\,
            I => \N__58477\
        );

    \I__13916\ : LocalMux
    port map (
            O => \N__58490\,
            I => \N__58474\
        );

    \I__13915\ : InMux
    port map (
            O => \N__58489\,
            I => \N__58470\
        );

    \I__13914\ : LocalMux
    port map (
            O => \N__58486\,
            I => \N__58465\
        );

    \I__13913\ : LocalMux
    port map (
            O => \N__58483\,
            I => \N__58465\
        );

    \I__13912\ : LocalMux
    port map (
            O => \N__58480\,
            I => \N__58462\
        );

    \I__13911\ : Span4Mux_v
    port map (
            O => \N__58477\,
            I => \N__58459\
        );

    \I__13910\ : Span4Mux_v
    port map (
            O => \N__58474\,
            I => \N__58456\
        );

    \I__13909\ : InMux
    port map (
            O => \N__58473\,
            I => \N__58452\
        );

    \I__13908\ : LocalMux
    port map (
            O => \N__58470\,
            I => \N__58449\
        );

    \I__13907\ : Span4Mux_h
    port map (
            O => \N__58465\,
            I => \N__58444\
        );

    \I__13906\ : Span4Mux_v
    port map (
            O => \N__58462\,
            I => \N__58444\
        );

    \I__13905\ : Span4Mux_h
    port map (
            O => \N__58459\,
            I => \N__58441\
        );

    \I__13904\ : Span4Mux_h
    port map (
            O => \N__58456\,
            I => \N__58437\
        );

    \I__13903\ : InMux
    port map (
            O => \N__58455\,
            I => \N__58434\
        );

    \I__13902\ : LocalMux
    port map (
            O => \N__58452\,
            I => \N__58431\
        );

    \I__13901\ : Span4Mux_v
    port map (
            O => \N__58449\,
            I => \N__58428\
        );

    \I__13900\ : Span4Mux_v
    port map (
            O => \N__58444\,
            I => \N__58425\
        );

    \I__13899\ : Span4Mux_h
    port map (
            O => \N__58441\,
            I => \N__58422\
        );

    \I__13898\ : CascadeMux
    port map (
            O => \N__58440\,
            I => \N__58419\
        );

    \I__13897\ : Span4Mux_v
    port map (
            O => \N__58437\,
            I => \N__58416\
        );

    \I__13896\ : LocalMux
    port map (
            O => \N__58434\,
            I => \N__58413\
        );

    \I__13895\ : Span12Mux_v
    port map (
            O => \N__58431\,
            I => \N__58406\
        );

    \I__13894\ : Sp12to4
    port map (
            O => \N__58428\,
            I => \N__58406\
        );

    \I__13893\ : Sp12to4
    port map (
            O => \N__58425\,
            I => \N__58406\
        );

    \I__13892\ : Span4Mux_v
    port map (
            O => \N__58422\,
            I => \N__58403\
        );

    \I__13891\ : InMux
    port map (
            O => \N__58419\,
            I => \N__58400\
        );

    \I__13890\ : Span4Mux_h
    port map (
            O => \N__58416\,
            I => \N__58395\
        );

    \I__13889\ : Span4Mux_h
    port map (
            O => \N__58413\,
            I => \N__58395\
        );

    \I__13888\ : Odrv12
    port map (
            O => \N__58406\,
            I => \I2C_top_level_inst1_s_data_oreg_14\
        );

    \I__13887\ : Odrv4
    port map (
            O => \N__58403\,
            I => \I2C_top_level_inst1_s_data_oreg_14\
        );

    \I__13886\ : LocalMux
    port map (
            O => \N__58400\,
            I => \I2C_top_level_inst1_s_data_oreg_14\
        );

    \I__13885\ : Odrv4
    port map (
            O => \N__58395\,
            I => \I2C_top_level_inst1_s_data_oreg_14\
        );

    \I__13884\ : InMux
    port map (
            O => \N__58386\,
            I => \N__58383\
        );

    \I__13883\ : LocalMux
    port map (
            O => \N__58383\,
            I => \N__58380\
        );

    \I__13882\ : Odrv4
    port map (
            O => \N__58380\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_14\
        );

    \I__13881\ : InMux
    port map (
            O => \N__58377\,
            I => \N__58373\
        );

    \I__13880\ : InMux
    port map (
            O => \N__58376\,
            I => \N__58370\
        );

    \I__13879\ : LocalMux
    port map (
            O => \N__58373\,
            I => \N__58365\
        );

    \I__13878\ : LocalMux
    port map (
            O => \N__58370\,
            I => \N__58365\
        );

    \I__13877\ : Span4Mux_h
    port map (
            O => \N__58365\,
            I => \N__58361\
        );

    \I__13876\ : InMux
    port map (
            O => \N__58364\,
            I => \N__58358\
        );

    \I__13875\ : Span4Mux_v
    port map (
            O => \N__58361\,
            I => \N__58352\
        );

    \I__13874\ : LocalMux
    port map (
            O => \N__58358\,
            I => \N__58352\
        );

    \I__13873\ : CascadeMux
    port map (
            O => \N__58357\,
            I => \N__58345\
        );

    \I__13872\ : Span4Mux_v
    port map (
            O => \N__58352\,
            I => \N__58342\
        );

    \I__13871\ : InMux
    port map (
            O => \N__58351\,
            I => \N__58339\
        );

    \I__13870\ : InMux
    port map (
            O => \N__58350\,
            I => \N__58336\
        );

    \I__13869\ : InMux
    port map (
            O => \N__58349\,
            I => \N__58333\
        );

    \I__13868\ : InMux
    port map (
            O => \N__58348\,
            I => \N__58329\
        );

    \I__13867\ : InMux
    port map (
            O => \N__58345\,
            I => \N__58326\
        );

    \I__13866\ : Span4Mux_v
    port map (
            O => \N__58342\,
            I => \N__58323\
        );

    \I__13865\ : LocalMux
    port map (
            O => \N__58339\,
            I => \N__58316\
        );

    \I__13864\ : LocalMux
    port map (
            O => \N__58336\,
            I => \N__58316\
        );

    \I__13863\ : LocalMux
    port map (
            O => \N__58333\,
            I => \N__58316\
        );

    \I__13862\ : InMux
    port map (
            O => \N__58332\,
            I => \N__58313\
        );

    \I__13861\ : LocalMux
    port map (
            O => \N__58329\,
            I => \N__58310\
        );

    \I__13860\ : LocalMux
    port map (
            O => \N__58326\,
            I => \N__58307\
        );

    \I__13859\ : Span4Mux_h
    port map (
            O => \N__58323\,
            I => \N__58302\
        );

    \I__13858\ : Span4Mux_v
    port map (
            O => \N__58316\,
            I => \N__58302\
        );

    \I__13857\ : LocalMux
    port map (
            O => \N__58313\,
            I => \N__58299\
        );

    \I__13856\ : Span4Mux_v
    port map (
            O => \N__58310\,
            I => \N__58296\
        );

    \I__13855\ : Span4Mux_v
    port map (
            O => \N__58307\,
            I => \N__58293\
        );

    \I__13854\ : Span4Mux_v
    port map (
            O => \N__58302\,
            I => \N__58290\
        );

    \I__13853\ : Span4Mux_h
    port map (
            O => \N__58299\,
            I => \N__58287\
        );

    \I__13852\ : Sp12to4
    port map (
            O => \N__58296\,
            I => \N__58284\
        );

    \I__13851\ : Span4Mux_v
    port map (
            O => \N__58293\,
            I => \N__58281\
        );

    \I__13850\ : Span4Mux_h
    port map (
            O => \N__58290\,
            I => \N__58276\
        );

    \I__13849\ : Span4Mux_h
    port map (
            O => \N__58287\,
            I => \N__58276\
        );

    \I__13848\ : Odrv12
    port map (
            O => \N__58284\,
            I => \I2C_top_level_inst1_s_data_oreg_13\
        );

    \I__13847\ : Odrv4
    port map (
            O => \N__58281\,
            I => \I2C_top_level_inst1_s_data_oreg_13\
        );

    \I__13846\ : Odrv4
    port map (
            O => \N__58276\,
            I => \I2C_top_level_inst1_s_data_oreg_13\
        );

    \I__13845\ : InMux
    port map (
            O => \N__58269\,
            I => \N__58266\
        );

    \I__13844\ : LocalMux
    port map (
            O => \N__58266\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_12\
        );

    \I__13843\ : InMux
    port map (
            O => \N__58263\,
            I => \N__58260\
        );

    \I__13842\ : LocalMux
    port map (
            O => \N__58260\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_13\
        );

    \I__13841\ : CascadeMux
    port map (
            O => \N__58257\,
            I => \N__58253\
        );

    \I__13840\ : InMux
    port map (
            O => \N__58256\,
            I => \N__58250\
        );

    \I__13839\ : InMux
    port map (
            O => \N__58253\,
            I => \N__58247\
        );

    \I__13838\ : LocalMux
    port map (
            O => \N__58250\,
            I => \N__58243\
        );

    \I__13837\ : LocalMux
    port map (
            O => \N__58247\,
            I => \N__58240\
        );

    \I__13836\ : InMux
    port map (
            O => \N__58246\,
            I => \N__58237\
        );

    \I__13835\ : Span4Mux_v
    port map (
            O => \N__58243\,
            I => \N__58232\
        );

    \I__13834\ : Span4Mux_v
    port map (
            O => \N__58240\,
            I => \N__58232\
        );

    \I__13833\ : LocalMux
    port map (
            O => \N__58237\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_0
        );

    \I__13832\ : Odrv4
    port map (
            O => \N__58232\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_0
        );

    \I__13831\ : InMux
    port map (
            O => \N__58227\,
            I => \N__58224\
        );

    \I__13830\ : LocalMux
    port map (
            O => \N__58224\,
            I => \N__58220\
        );

    \I__13829\ : InMux
    port map (
            O => \N__58223\,
            I => \N__58217\
        );

    \I__13828\ : Span4Mux_v
    port map (
            O => \N__58220\,
            I => \N__58212\
        );

    \I__13827\ : LocalMux
    port map (
            O => \N__58217\,
            I => \N__58212\
        );

    \I__13826\ : Span4Mux_v
    port map (
            O => \N__58212\,
            I => \N__58208\
        );

    \I__13825\ : InMux
    port map (
            O => \N__58211\,
            I => \N__58205\
        );

    \I__13824\ : Odrv4
    port map (
            O => \N__58208\,
            I => cemf_module_64ch_ctrl_inst1_data_config_0
        );

    \I__13823\ : LocalMux
    port map (
            O => \N__58205\,
            I => cemf_module_64ch_ctrl_inst1_data_config_0
        );

    \I__13822\ : InMux
    port map (
            O => \N__58200\,
            I => \N__58191\
        );

    \I__13821\ : InMux
    port map (
            O => \N__58199\,
            I => \N__58191\
        );

    \I__13820\ : CascadeMux
    port map (
            O => \N__58198\,
            I => \N__58187\
        );

    \I__13819\ : InMux
    port map (
            O => \N__58197\,
            I => \N__58174\
        );

    \I__13818\ : InMux
    port map (
            O => \N__58196\,
            I => \N__58174\
        );

    \I__13817\ : LocalMux
    port map (
            O => \N__58191\,
            I => \N__58171\
        );

    \I__13816\ : InMux
    port map (
            O => \N__58190\,
            I => \N__58166\
        );

    \I__13815\ : InMux
    port map (
            O => \N__58187\,
            I => \N__58166\
        );

    \I__13814\ : InMux
    port map (
            O => \N__58186\,
            I => \N__58160\
        );

    \I__13813\ : InMux
    port map (
            O => \N__58185\,
            I => \N__58160\
        );

    \I__13812\ : InMux
    port map (
            O => \N__58184\,
            I => \N__58153\
        );

    \I__13811\ : InMux
    port map (
            O => \N__58183\,
            I => \N__58148\
        );

    \I__13810\ : InMux
    port map (
            O => \N__58182\,
            I => \N__58148\
        );

    \I__13809\ : InMux
    port map (
            O => \N__58181\,
            I => \N__58143\
        );

    \I__13808\ : InMux
    port map (
            O => \N__58180\,
            I => \N__58143\
        );

    \I__13807\ : InMux
    port map (
            O => \N__58179\,
            I => \N__58140\
        );

    \I__13806\ : LocalMux
    port map (
            O => \N__58174\,
            I => \N__58135\
        );

    \I__13805\ : Span4Mux_v
    port map (
            O => \N__58171\,
            I => \N__58135\
        );

    \I__13804\ : LocalMux
    port map (
            O => \N__58166\,
            I => \N__58132\
        );

    \I__13803\ : InMux
    port map (
            O => \N__58165\,
            I => \N__58129\
        );

    \I__13802\ : LocalMux
    port map (
            O => \N__58160\,
            I => \N__58126\
        );

    \I__13801\ : InMux
    port map (
            O => \N__58159\,
            I => \N__58121\
        );

    \I__13800\ : InMux
    port map (
            O => \N__58158\,
            I => \N__58121\
        );

    \I__13799\ : InMux
    port map (
            O => \N__58157\,
            I => \N__58117\
        );

    \I__13798\ : InMux
    port map (
            O => \N__58156\,
            I => \N__58114\
        );

    \I__13797\ : LocalMux
    port map (
            O => \N__58153\,
            I => \N__58105\
        );

    \I__13796\ : LocalMux
    port map (
            O => \N__58148\,
            I => \N__58105\
        );

    \I__13795\ : LocalMux
    port map (
            O => \N__58143\,
            I => \N__58102\
        );

    \I__13794\ : LocalMux
    port map (
            O => \N__58140\,
            I => \N__58099\
        );

    \I__13793\ : Span4Mux_h
    port map (
            O => \N__58135\,
            I => \N__58094\
        );

    \I__13792\ : Span4Mux_h
    port map (
            O => \N__58132\,
            I => \N__58094\
        );

    \I__13791\ : LocalMux
    port map (
            O => \N__58129\,
            I => \N__58089\
        );

    \I__13790\ : Span4Mux_h
    port map (
            O => \N__58126\,
            I => \N__58089\
        );

    \I__13789\ : LocalMux
    port map (
            O => \N__58121\,
            I => \N__58086\
        );

    \I__13788\ : InMux
    port map (
            O => \N__58120\,
            I => \N__58083\
        );

    \I__13787\ : LocalMux
    port map (
            O => \N__58117\,
            I => \N__58078\
        );

    \I__13786\ : LocalMux
    port map (
            O => \N__58114\,
            I => \N__58078\
        );

    \I__13785\ : InMux
    port map (
            O => \N__58113\,
            I => \N__58073\
        );

    \I__13784\ : InMux
    port map (
            O => \N__58112\,
            I => \N__58073\
        );

    \I__13783\ : InMux
    port map (
            O => \N__58111\,
            I => \N__58068\
        );

    \I__13782\ : InMux
    port map (
            O => \N__58110\,
            I => \N__58068\
        );

    \I__13781\ : Span4Mux_v
    port map (
            O => \N__58105\,
            I => \N__58065\
        );

    \I__13780\ : Span4Mux_v
    port map (
            O => \N__58102\,
            I => \N__58060\
        );

    \I__13779\ : Span4Mux_v
    port map (
            O => \N__58099\,
            I => \N__58060\
        );

    \I__13778\ : Span4Mux_v
    port map (
            O => \N__58094\,
            I => \N__58057\
        );

    \I__13777\ : Span4Mux_v
    port map (
            O => \N__58089\,
            I => \N__58050\
        );

    \I__13776\ : Span4Mux_v
    port map (
            O => \N__58086\,
            I => \N__58050\
        );

    \I__13775\ : LocalMux
    port map (
            O => \N__58083\,
            I => \N__58050\
        );

    \I__13774\ : Span4Mux_v
    port map (
            O => \N__58078\,
            I => \N__58045\
        );

    \I__13773\ : LocalMux
    port map (
            O => \N__58073\,
            I => \N__58045\
        );

    \I__13772\ : LocalMux
    port map (
            O => \N__58068\,
            I => \N__58038\
        );

    \I__13771\ : Sp12to4
    port map (
            O => \N__58065\,
            I => \N__58038\
        );

    \I__13770\ : Sp12to4
    port map (
            O => \N__58060\,
            I => \N__58038\
        );

    \I__13769\ : Sp12to4
    port map (
            O => \N__58057\,
            I => \N__58035\
        );

    \I__13768\ : Span4Mux_h
    port map (
            O => \N__58050\,
            I => \N__58032\
        );

    \I__13767\ : Sp12to4
    port map (
            O => \N__58045\,
            I => \N__58027\
        );

    \I__13766\ : Span12Mux_h
    port map (
            O => \N__58038\,
            I => \N__58027\
        );

    \I__13765\ : Span12Mux_v
    port map (
            O => \N__58035\,
            I => \N__58024\
        );

    \I__13764\ : Odrv4
    port map (
            O => \N__58032\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0\
        );

    \I__13763\ : Odrv12
    port map (
            O => \N__58027\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0\
        );

    \I__13762\ : Odrv12
    port map (
            O => \N__58024\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0\
        );

    \I__13761\ : InMux
    port map (
            O => \N__58017\,
            I => \N__58008\
        );

    \I__13760\ : InMux
    port map (
            O => \N__58016\,
            I => \N__58008\
        );

    \I__13759\ : InMux
    port map (
            O => \N__58015\,
            I => \N__58001\
        );

    \I__13758\ : InMux
    port map (
            O => \N__58014\,
            I => \N__57996\
        );

    \I__13757\ : InMux
    port map (
            O => \N__58013\,
            I => \N__57996\
        );

    \I__13756\ : LocalMux
    port map (
            O => \N__58008\,
            I => \N__57993\
        );

    \I__13755\ : InMux
    port map (
            O => \N__58007\,
            I => \N__57982\
        );

    \I__13754\ : InMux
    port map (
            O => \N__58006\,
            I => \N__57982\
        );

    \I__13753\ : InMux
    port map (
            O => \N__58005\,
            I => \N__57973\
        );

    \I__13752\ : InMux
    port map (
            O => \N__58004\,
            I => \N__57973\
        );

    \I__13751\ : LocalMux
    port map (
            O => \N__58001\,
            I => \N__57970\
        );

    \I__13750\ : LocalMux
    port map (
            O => \N__57996\,
            I => \N__57967\
        );

    \I__13749\ : Span4Mux_v
    port map (
            O => \N__57993\,
            I => \N__57964\
        );

    \I__13748\ : InMux
    port map (
            O => \N__57992\,
            I => \N__57959\
        );

    \I__13747\ : InMux
    port map (
            O => \N__57991\,
            I => \N__57959\
        );

    \I__13746\ : InMux
    port map (
            O => \N__57990\,
            I => \N__57954\
        );

    \I__13745\ : InMux
    port map (
            O => \N__57989\,
            I => \N__57954\
        );

    \I__13744\ : InMux
    port map (
            O => \N__57988\,
            I => \N__57949\
        );

    \I__13743\ : InMux
    port map (
            O => \N__57987\,
            I => \N__57949\
        );

    \I__13742\ : LocalMux
    port map (
            O => \N__57982\,
            I => \N__57946\
        );

    \I__13741\ : InMux
    port map (
            O => \N__57981\,
            I => \N__57943\
        );

    \I__13740\ : InMux
    port map (
            O => \N__57980\,
            I => \N__57936\
        );

    \I__13739\ : InMux
    port map (
            O => \N__57979\,
            I => \N__57936\
        );

    \I__13738\ : InMux
    port map (
            O => \N__57978\,
            I => \N__57932\
        );

    \I__13737\ : LocalMux
    port map (
            O => \N__57973\,
            I => \N__57927\
        );

    \I__13736\ : Span4Mux_v
    port map (
            O => \N__57970\,
            I => \N__57927\
        );

    \I__13735\ : Span4Mux_v
    port map (
            O => \N__57967\,
            I => \N__57923\
        );

    \I__13734\ : Span4Mux_h
    port map (
            O => \N__57964\,
            I => \N__57918\
        );

    \I__13733\ : LocalMux
    port map (
            O => \N__57959\,
            I => \N__57918\
        );

    \I__13732\ : LocalMux
    port map (
            O => \N__57954\,
            I => \N__57915\
        );

    \I__13731\ : LocalMux
    port map (
            O => \N__57949\,
            I => \N__57911\
        );

    \I__13730\ : Span4Mux_h
    port map (
            O => \N__57946\,
            I => \N__57906\
        );

    \I__13729\ : LocalMux
    port map (
            O => \N__57943\,
            I => \N__57906\
        );

    \I__13728\ : InMux
    port map (
            O => \N__57942\,
            I => \N__57901\
        );

    \I__13727\ : InMux
    port map (
            O => \N__57941\,
            I => \N__57901\
        );

    \I__13726\ : LocalMux
    port map (
            O => \N__57936\,
            I => \N__57898\
        );

    \I__13725\ : InMux
    port map (
            O => \N__57935\,
            I => \N__57895\
        );

    \I__13724\ : LocalMux
    port map (
            O => \N__57932\,
            I => \N__57890\
        );

    \I__13723\ : Span4Mux_h
    port map (
            O => \N__57927\,
            I => \N__57890\
        );

    \I__13722\ : InMux
    port map (
            O => \N__57926\,
            I => \N__57887\
        );

    \I__13721\ : Span4Mux_h
    port map (
            O => \N__57923\,
            I => \N__57880\
        );

    \I__13720\ : Span4Mux_v
    port map (
            O => \N__57918\,
            I => \N__57880\
        );

    \I__13719\ : Span4Mux_v
    port map (
            O => \N__57915\,
            I => \N__57880\
        );

    \I__13718\ : InMux
    port map (
            O => \N__57914\,
            I => \N__57877\
        );

    \I__13717\ : Span4Mux_v
    port map (
            O => \N__57911\,
            I => \N__57872\
        );

    \I__13716\ : Span4Mux_v
    port map (
            O => \N__57906\,
            I => \N__57872\
        );

    \I__13715\ : LocalMux
    port map (
            O => \N__57901\,
            I => \N__57869\
        );

    \I__13714\ : Span4Mux_h
    port map (
            O => \N__57898\,
            I => \N__57866\
        );

    \I__13713\ : LocalMux
    port map (
            O => \N__57895\,
            I => \N__57861\
        );

    \I__13712\ : Span4Mux_h
    port map (
            O => \N__57890\,
            I => \N__57861\
        );

    \I__13711\ : LocalMux
    port map (
            O => \N__57887\,
            I => \N__57852\
        );

    \I__13710\ : Sp12to4
    port map (
            O => \N__57880\,
            I => \N__57852\
        );

    \I__13709\ : LocalMux
    port map (
            O => \N__57877\,
            I => \N__57852\
        );

    \I__13708\ : Sp12to4
    port map (
            O => \N__57872\,
            I => \N__57852\
        );

    \I__13707\ : Span4Mux_v
    port map (
            O => \N__57869\,
            I => \N__57849\
        );

    \I__13706\ : Span4Mux_h
    port map (
            O => \N__57866\,
            I => \N__57846\
        );

    \I__13705\ : Sp12to4
    port map (
            O => \N__57861\,
            I => \N__57841\
        );

    \I__13704\ : Span12Mux_h
    port map (
            O => \N__57852\,
            I => \N__57841\
        );

    \I__13703\ : Odrv4
    port map (
            O => \N__57849\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273\
        );

    \I__13702\ : Odrv4
    port map (
            O => \N__57846\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273\
        );

    \I__13701\ : Odrv12
    port map (
            O => \N__57841\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273\
        );

    \I__13700\ : InMux
    port map (
            O => \N__57834\,
            I => \N__57830\
        );

    \I__13699\ : CascadeMux
    port map (
            O => \N__57833\,
            I => \N__57827\
        );

    \I__13698\ : LocalMux
    port map (
            O => \N__57830\,
            I => \N__57823\
        );

    \I__13697\ : InMux
    port map (
            O => \N__57827\,
            I => \N__57820\
        );

    \I__13696\ : InMux
    port map (
            O => \N__57826\,
            I => \N__57817\
        );

    \I__13695\ : Span12Mux_h
    port map (
            O => \N__57823\,
            I => \N__57814\
        );

    \I__13694\ : LocalMux
    port map (
            O => \N__57820\,
            I => \N__57811\
        );

    \I__13693\ : LocalMux
    port map (
            O => \N__57817\,
            I => \N__57808\
        );

    \I__13692\ : Odrv12
    port map (
            O => \N__57814\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_1
        );

    \I__13691\ : Odrv12
    port map (
            O => \N__57811\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_1
        );

    \I__13690\ : Odrv4
    port map (
            O => \N__57808\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_1
        );

    \I__13689\ : InMux
    port map (
            O => \N__57801\,
            I => \N__57796\
        );

    \I__13688\ : InMux
    port map (
            O => \N__57800\,
            I => \N__57793\
        );

    \I__13687\ : InMux
    port map (
            O => \N__57799\,
            I => \N__57790\
        );

    \I__13686\ : LocalMux
    port map (
            O => \N__57796\,
            I => \N__57787\
        );

    \I__13685\ : LocalMux
    port map (
            O => \N__57793\,
            I => \N__57784\
        );

    \I__13684\ : LocalMux
    port map (
            O => \N__57790\,
            I => \N__57781\
        );

    \I__13683\ : Span4Mux_v
    port map (
            O => \N__57787\,
            I => \N__57778\
        );

    \I__13682\ : Span4Mux_v
    port map (
            O => \N__57784\,
            I => \N__57775\
        );

    \I__13681\ : Span4Mux_h
    port map (
            O => \N__57781\,
            I => \N__57772\
        );

    \I__13680\ : Span4Mux_h
    port map (
            O => \N__57778\,
            I => \N__57769\
        );

    \I__13679\ : Span4Mux_h
    port map (
            O => \N__57775\,
            I => \N__57764\
        );

    \I__13678\ : Span4Mux_h
    port map (
            O => \N__57772\,
            I => \N__57764\
        );

    \I__13677\ : Span4Mux_h
    port map (
            O => \N__57769\,
            I => \N__57761\
        );

    \I__13676\ : Span4Mux_h
    port map (
            O => \N__57764\,
            I => \N__57758\
        );

    \I__13675\ : Odrv4
    port map (
            O => \N__57761\,
            I => cemf_module_64ch_ctrl_inst1_data_config_1
        );

    \I__13674\ : Odrv4
    port map (
            O => \N__57758\,
            I => cemf_module_64ch_ctrl_inst1_data_config_1
        );

    \I__13673\ : InMux
    port map (
            O => \N__57753\,
            I => \N__57750\
        );

    \I__13672\ : LocalMux
    port map (
            O => \N__57750\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1776\
        );

    \I__13671\ : CascadeMux
    port map (
            O => \N__57747\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0_cascade_\
        );

    \I__13670\ : InMux
    port map (
            O => \N__57744\,
            I => \N__57740\
        );

    \I__13669\ : InMux
    port map (
            O => \N__57743\,
            I => \N__57737\
        );

    \I__13668\ : LocalMux
    port map (
            O => \N__57740\,
            I => \N__57731\
        );

    \I__13667\ : LocalMux
    port map (
            O => \N__57737\,
            I => \N__57731\
        );

    \I__13666\ : InMux
    port map (
            O => \N__57736\,
            I => \N__57728\
        );

    \I__13665\ : Span4Mux_v
    port map (
            O => \N__57731\,
            I => \N__57723\
        );

    \I__13664\ : LocalMux
    port map (
            O => \N__57728\,
            I => \N__57723\
        );

    \I__13663\ : Span4Mux_v
    port map (
            O => \N__57723\,
            I => \N__57720\
        );

    \I__13662\ : Sp12to4
    port map (
            O => \N__57720\,
            I => \N__57715\
        );

    \I__13661\ : InMux
    port map (
            O => \N__57719\,
            I => \N__57710\
        );

    \I__13660\ : InMux
    port map (
            O => \N__57718\,
            I => \N__57710\
        );

    \I__13659\ : Odrv12
    port map (
            O => \N__57715\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11\
        );

    \I__13658\ : LocalMux
    port map (
            O => \N__57710\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11\
        );

    \I__13657\ : InMux
    port map (
            O => \N__57705\,
            I => \N__57702\
        );

    \I__13656\ : LocalMux
    port map (
            O => \N__57702\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_209\
        );

    \I__13655\ : IoInMux
    port map (
            O => \N__57699\,
            I => \N__57696\
        );

    \I__13654\ : LocalMux
    port map (
            O => \N__57696\,
            I => \N__57693\
        );

    \I__13653\ : IoSpan4Mux
    port map (
            O => \N__57693\,
            I => \N__57690\
        );

    \I__13652\ : Span4Mux_s1_h
    port map (
            O => \N__57690\,
            I => \N__57687\
        );

    \I__13651\ : Span4Mux_h
    port map (
            O => \N__57687\,
            I => \N__57682\
        );

    \I__13650\ : InMux
    port map (
            O => \N__57686\,
            I => \N__57679\
        );

    \I__13649\ : InMux
    port map (
            O => \N__57685\,
            I => \N__57676\
        );

    \I__13648\ : Span4Mux_h
    port map (
            O => \N__57682\,
            I => \N__57671\
        );

    \I__13647\ : LocalMux
    port map (
            O => \N__57679\,
            I => \N__57671\
        );

    \I__13646\ : LocalMux
    port map (
            O => \N__57676\,
            I => \N__57668\
        );

    \I__13645\ : Span4Mux_v
    port map (
            O => \N__57671\,
            I => \N__57665\
        );

    \I__13644\ : Span4Mux_v
    port map (
            O => \N__57668\,
            I => \N__57662\
        );

    \I__13643\ : Span4Mux_v
    port map (
            O => \N__57665\,
            I => \N__57659\
        );

    \I__13642\ : Span4Mux_h
    port map (
            O => \N__57662\,
            I => \N__57656\
        );

    \I__13641\ : Sp12to4
    port map (
            O => \N__57659\,
            I => \N__57653\
        );

    \I__13640\ : Sp12to4
    port map (
            O => \N__57656\,
            I => \N__57650\
        );

    \I__13639\ : Span12Mux_h
    port map (
            O => \N__57653\,
            I => \N__57645\
        );

    \I__13638\ : Span12Mux_v
    port map (
            O => \N__57650\,
            I => \N__57645\
        );

    \I__13637\ : Odrv12
    port map (
            O => \N__57645\,
            I => s_sda_i
        );

    \I__13636\ : InMux
    port map (
            O => \N__57642\,
            I => \N__57639\
        );

    \I__13635\ : LocalMux
    port map (
            O => \N__57639\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_0\
        );

    \I__13634\ : InMux
    port map (
            O => \N__57636\,
            I => \N__57633\
        );

    \I__13633\ : LocalMux
    port map (
            O => \N__57633\,
            I => \N__57629\
        );

    \I__13632\ : InMux
    port map (
            O => \N__57632\,
            I => \N__57624\
        );

    \I__13631\ : Span4Mux_v
    port map (
            O => \N__57629\,
            I => \N__57621\
        );

    \I__13630\ : InMux
    port map (
            O => \N__57628\,
            I => \N__57615\
        );

    \I__13629\ : InMux
    port map (
            O => \N__57627\,
            I => \N__57612\
        );

    \I__13628\ : LocalMux
    port map (
            O => \N__57624\,
            I => \N__57609\
        );

    \I__13627\ : Span4Mux_h
    port map (
            O => \N__57621\,
            I => \N__57605\
        );

    \I__13626\ : InMux
    port map (
            O => \N__57620\,
            I => \N__57602\
        );

    \I__13625\ : InMux
    port map (
            O => \N__57619\,
            I => \N__57598\
        );

    \I__13624\ : InMux
    port map (
            O => \N__57618\,
            I => \N__57595\
        );

    \I__13623\ : LocalMux
    port map (
            O => \N__57615\,
            I => \N__57592\
        );

    \I__13622\ : LocalMux
    port map (
            O => \N__57612\,
            I => \N__57589\
        );

    \I__13621\ : Span4Mux_h
    port map (
            O => \N__57609\,
            I => \N__57586\
        );

    \I__13620\ : CascadeMux
    port map (
            O => \N__57608\,
            I => \N__57583\
        );

    \I__13619\ : Span4Mux_h
    port map (
            O => \N__57605\,
            I => \N__57580\
        );

    \I__13618\ : LocalMux
    port map (
            O => \N__57602\,
            I => \N__57577\
        );

    \I__13617\ : InMux
    port map (
            O => \N__57601\,
            I => \N__57574\
        );

    \I__13616\ : LocalMux
    port map (
            O => \N__57598\,
            I => \N__57571\
        );

    \I__13615\ : LocalMux
    port map (
            O => \N__57595\,
            I => \N__57568\
        );

    \I__13614\ : Span4Mux_h
    port map (
            O => \N__57592\,
            I => \N__57561\
        );

    \I__13613\ : Span4Mux_h
    port map (
            O => \N__57589\,
            I => \N__57561\
        );

    \I__13612\ : Span4Mux_h
    port map (
            O => \N__57586\,
            I => \N__57561\
        );

    \I__13611\ : InMux
    port map (
            O => \N__57583\,
            I => \N__57558\
        );

    \I__13610\ : Span4Mux_h
    port map (
            O => \N__57580\,
            I => \N__57555\
        );

    \I__13609\ : Odrv12
    port map (
            O => \N__57577\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13608\ : LocalMux
    port map (
            O => \N__57574\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13607\ : Odrv4
    port map (
            O => \N__57571\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13606\ : Odrv12
    port map (
            O => \N__57568\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13605\ : Odrv4
    port map (
            O => \N__57561\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13604\ : LocalMux
    port map (
            O => \N__57558\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13603\ : Odrv4
    port map (
            O => \N__57555\,
            I => \I2C_top_level_inst1_s_data_oreg_16\
        );

    \I__13602\ : InMux
    port map (
            O => \N__57540\,
            I => \N__57537\
        );

    \I__13601\ : LocalMux
    port map (
            O => \N__57537\,
            I => \N__57531\
        );

    \I__13600\ : InMux
    port map (
            O => \N__57536\,
            I => \N__57528\
        );

    \I__13599\ : InMux
    port map (
            O => \N__57535\,
            I => \N__57525\
        );

    \I__13598\ : InMux
    port map (
            O => \N__57534\,
            I => \N__57521\
        );

    \I__13597\ : Span4Mux_v
    port map (
            O => \N__57531\,
            I => \N__57513\
        );

    \I__13596\ : LocalMux
    port map (
            O => \N__57528\,
            I => \N__57513\
        );

    \I__13595\ : LocalMux
    port map (
            O => \N__57525\,
            I => \N__57513\
        );

    \I__13594\ : InMux
    port map (
            O => \N__57524\,
            I => \N__57510\
        );

    \I__13593\ : LocalMux
    port map (
            O => \N__57521\,
            I => \N__57506\
        );

    \I__13592\ : InMux
    port map (
            O => \N__57520\,
            I => \N__57503\
        );

    \I__13591\ : Span4Mux_h
    port map (
            O => \N__57513\,
            I => \N__57500\
        );

    \I__13590\ : LocalMux
    port map (
            O => \N__57510\,
            I => \N__57497\
        );

    \I__13589\ : InMux
    port map (
            O => \N__57509\,
            I => \N__57493\
        );

    \I__13588\ : Span4Mux_v
    port map (
            O => \N__57506\,
            I => \N__57490\
        );

    \I__13587\ : LocalMux
    port map (
            O => \N__57503\,
            I => \N__57487\
        );

    \I__13586\ : Span4Mux_v
    port map (
            O => \N__57500\,
            I => \N__57482\
        );

    \I__13585\ : Span4Mux_v
    port map (
            O => \N__57497\,
            I => \N__57482\
        );

    \I__13584\ : InMux
    port map (
            O => \N__57496\,
            I => \N__57479\
        );

    \I__13583\ : LocalMux
    port map (
            O => \N__57493\,
            I => \N__57476\
        );

    \I__13582\ : Span4Mux_h
    port map (
            O => \N__57490\,
            I => \N__57472\
        );

    \I__13581\ : Span4Mux_v
    port map (
            O => \N__57487\,
            I => \N__57469\
        );

    \I__13580\ : Sp12to4
    port map (
            O => \N__57482\,
            I => \N__57464\
        );

    \I__13579\ : LocalMux
    port map (
            O => \N__57479\,
            I => \N__57464\
        );

    \I__13578\ : Span4Mux_v
    port map (
            O => \N__57476\,
            I => \N__57461\
        );

    \I__13577\ : CascadeMux
    port map (
            O => \N__57475\,
            I => \N__57458\
        );

    \I__13576\ : Span4Mux_h
    port map (
            O => \N__57472\,
            I => \N__57453\
        );

    \I__13575\ : Span4Mux_v
    port map (
            O => \N__57469\,
            I => \N__57453\
        );

    \I__13574\ : Span12Mux_h
    port map (
            O => \N__57464\,
            I => \N__57450\
        );

    \I__13573\ : Span4Mux_h
    port map (
            O => \N__57461\,
            I => \N__57447\
        );

    \I__13572\ : InMux
    port map (
            O => \N__57458\,
            I => \N__57444\
        );

    \I__13571\ : Odrv4
    port map (
            O => \N__57453\,
            I => \I2C_top_level_inst1_s_data_oreg_15\
        );

    \I__13570\ : Odrv12
    port map (
            O => \N__57450\,
            I => \I2C_top_level_inst1_s_data_oreg_15\
        );

    \I__13569\ : Odrv4
    port map (
            O => \N__57447\,
            I => \I2C_top_level_inst1_s_data_oreg_15\
        );

    \I__13568\ : LocalMux
    port map (
            O => \N__57444\,
            I => \I2C_top_level_inst1_s_data_oreg_15\
        );

    \I__13567\ : InMux
    port map (
            O => \N__57435\,
            I => \N__57432\
        );

    \I__13566\ : LocalMux
    port map (
            O => \N__57432\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_15\
        );

    \I__13565\ : InMux
    port map (
            O => \N__57429\,
            I => \N__57426\
        );

    \I__13564\ : LocalMux
    port map (
            O => \N__57426\,
            I => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_16\
        );

    \I__13563\ : InMux
    port map (
            O => \N__57423\,
            I => \N__57420\
        );

    \I__13562\ : LocalMux
    port map (
            O => \N__57420\,
            I => \N__57415\
        );

    \I__13561\ : InMux
    port map (
            O => \N__57419\,
            I => \N__57409\
        );

    \I__13560\ : InMux
    port map (
            O => \N__57418\,
            I => \N__57406\
        );

    \I__13559\ : Span4Mux_v
    port map (
            O => \N__57415\,
            I => \N__57403\
        );

    \I__13558\ : InMux
    port map (
            O => \N__57414\,
            I => \N__57400\
        );

    \I__13557\ : InMux
    port map (
            O => \N__57413\,
            I => \N__57397\
        );

    \I__13556\ : InMux
    port map (
            O => \N__57412\,
            I => \N__57394\
        );

    \I__13555\ : LocalMux
    port map (
            O => \N__57409\,
            I => \N__57389\
        );

    \I__13554\ : LocalMux
    port map (
            O => \N__57406\,
            I => \N__57386\
        );

    \I__13553\ : Span4Mux_h
    port map (
            O => \N__57403\,
            I => \N__57383\
        );

    \I__13552\ : LocalMux
    port map (
            O => \N__57400\,
            I => \N__57380\
        );

    \I__13551\ : LocalMux
    port map (
            O => \N__57397\,
            I => \N__57375\
        );

    \I__13550\ : LocalMux
    port map (
            O => \N__57394\,
            I => \N__57375\
        );

    \I__13549\ : InMux
    port map (
            O => \N__57393\,
            I => \N__57371\
        );

    \I__13548\ : InMux
    port map (
            O => \N__57392\,
            I => \N__57368\
        );

    \I__13547\ : Span4Mux_v
    port map (
            O => \N__57389\,
            I => \N__57361\
        );

    \I__13546\ : Span4Mux_v
    port map (
            O => \N__57386\,
            I => \N__57361\
        );

    \I__13545\ : Span4Mux_v
    port map (
            O => \N__57383\,
            I => \N__57361\
        );

    \I__13544\ : Span4Mux_v
    port map (
            O => \N__57380\,
            I => \N__57356\
        );

    \I__13543\ : Span4Mux_v
    port map (
            O => \N__57375\,
            I => \N__57356\
        );

    \I__13542\ : CascadeMux
    port map (
            O => \N__57374\,
            I => \N__57353\
        );

    \I__13541\ : LocalMux
    port map (
            O => \N__57371\,
            I => \N__57350\
        );

    \I__13540\ : LocalMux
    port map (
            O => \N__57368\,
            I => \N__57343\
        );

    \I__13539\ : Sp12to4
    port map (
            O => \N__57361\,
            I => \N__57343\
        );

    \I__13538\ : Sp12to4
    port map (
            O => \N__57356\,
            I => \N__57343\
        );

    \I__13537\ : InMux
    port map (
            O => \N__57353\,
            I => \N__57340\
        );

    \I__13536\ : Span4Mux_h
    port map (
            O => \N__57350\,
            I => \N__57337\
        );

    \I__13535\ : Odrv12
    port map (
            O => \N__57343\,
            I => \I2C_top_level_inst1_s_data_oreg_17\
        );

    \I__13534\ : LocalMux
    port map (
            O => \N__57340\,
            I => \I2C_top_level_inst1_s_data_oreg_17\
        );

    \I__13533\ : Odrv4
    port map (
            O => \N__57337\,
            I => \I2C_top_level_inst1_s_data_oreg_17\
        );

    \I__13532\ : InMux
    port map (
            O => \N__57330\,
            I => \N__57327\
        );

    \I__13531\ : LocalMux
    port map (
            O => \N__57327\,
            I => \N__57324\
        );

    \I__13530\ : Span4Mux_h
    port map (
            O => \N__57324\,
            I => \N__57320\
        );

    \I__13529\ : InMux
    port map (
            O => \N__57323\,
            I => \N__57316\
        );

    \I__13528\ : Span4Mux_h
    port map (
            O => \N__57320\,
            I => \N__57313\
        );

    \I__13527\ : InMux
    port map (
            O => \N__57319\,
            I => \N__57310\
        );

    \I__13526\ : LocalMux
    port map (
            O => \N__57316\,
            I => \N__57307\
        );

    \I__13525\ : Odrv4
    port map (
            O => \N__57313\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_19
        );

    \I__13524\ : LocalMux
    port map (
            O => \N__57310\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_19
        );

    \I__13523\ : Odrv12
    port map (
            O => \N__57307\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_19
        );

    \I__13522\ : InMux
    port map (
            O => \N__57300\,
            I => \N__57297\
        );

    \I__13521\ : LocalMux
    port map (
            O => \N__57297\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_211\
        );

    \I__13520\ : CascadeMux
    port map (
            O => \N__57294\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1653_cascade_\
        );

    \I__13519\ : CascadeMux
    port map (
            O => \N__57291\,
            I => \N__57288\
        );

    \I__13518\ : InMux
    port map (
            O => \N__57288\,
            I => \N__57284\
        );

    \I__13517\ : InMux
    port map (
            O => \N__57287\,
            I => \N__57281\
        );

    \I__13516\ : LocalMux
    port map (
            O => \N__57284\,
            I => \N__57278\
        );

    \I__13515\ : LocalMux
    port map (
            O => \N__57281\,
            I => \N__57275\
        );

    \I__13514\ : Span4Mux_v
    port map (
            O => \N__57278\,
            I => \N__57272\
        );

    \I__13513\ : Odrv4
    port map (
            O => \N__57275\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0\
        );

    \I__13512\ : Odrv4
    port map (
            O => \N__57272\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0\
        );

    \I__13511\ : CascadeMux
    port map (
            O => \N__57267\,
            I => \N__57264\
        );

    \I__13510\ : InMux
    port map (
            O => \N__57264\,
            I => \N__57261\
        );

    \I__13509\ : LocalMux
    port map (
            O => \N__57261\,
            I => \N__57258\
        );

    \I__13508\ : Odrv4
    port map (
            O => \N__57258\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_122_0\
        );

    \I__13507\ : InMux
    port map (
            O => \N__57255\,
            I => \N__57252\
        );

    \I__13506\ : LocalMux
    port map (
            O => \N__57252\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_208\
        );

    \I__13505\ : InMux
    port map (
            O => \N__57249\,
            I => \N__57243\
        );

    \I__13504\ : InMux
    port map (
            O => \N__57248\,
            I => \N__57243\
        );

    \I__13503\ : LocalMux
    port map (
            O => \N__57243\,
            I => \N__57239\
        );

    \I__13502\ : InMux
    port map (
            O => \N__57242\,
            I => \N__57234\
        );

    \I__13501\ : Span4Mux_h
    port map (
            O => \N__57239\,
            I => \N__57231\
        );

    \I__13500\ : InMux
    port map (
            O => \N__57238\,
            I => \N__57228\
        );

    \I__13499\ : InMux
    port map (
            O => \N__57237\,
            I => \N__57224\
        );

    \I__13498\ : LocalMux
    port map (
            O => \N__57234\,
            I => \N__57220\
        );

    \I__13497\ : Span4Mux_h
    port map (
            O => \N__57231\,
            I => \N__57217\
        );

    \I__13496\ : LocalMux
    port map (
            O => \N__57228\,
            I => \N__57213\
        );

    \I__13495\ : CascadeMux
    port map (
            O => \N__57227\,
            I => \N__57210\
        );

    \I__13494\ : LocalMux
    port map (
            O => \N__57224\,
            I => \N__57205\
        );

    \I__13493\ : InMux
    port map (
            O => \N__57223\,
            I => \N__57202\
        );

    \I__13492\ : Span4Mux_h
    port map (
            O => \N__57220\,
            I => \N__57197\
        );

    \I__13491\ : Span4Mux_v
    port map (
            O => \N__57217\,
            I => \N__57197\
        );

    \I__13490\ : CascadeMux
    port map (
            O => \N__57216\,
            I => \N__57194\
        );

    \I__13489\ : Span4Mux_h
    port map (
            O => \N__57213\,
            I => \N__57191\
        );

    \I__13488\ : InMux
    port map (
            O => \N__57210\,
            I => \N__57188\
        );

    \I__13487\ : InMux
    port map (
            O => \N__57209\,
            I => \N__57185\
        );

    \I__13486\ : InMux
    port map (
            O => \N__57208\,
            I => \N__57182\
        );

    \I__13485\ : Span4Mux_v
    port map (
            O => \N__57205\,
            I => \N__57179\
        );

    \I__13484\ : LocalMux
    port map (
            O => \N__57202\,
            I => \N__57176\
        );

    \I__13483\ : Span4Mux_h
    port map (
            O => \N__57197\,
            I => \N__57173\
        );

    \I__13482\ : InMux
    port map (
            O => \N__57194\,
            I => \N__57170\
        );

    \I__13481\ : Span4Mux_h
    port map (
            O => \N__57191\,
            I => \N__57167\
        );

    \I__13480\ : LocalMux
    port map (
            O => \N__57188\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13479\ : LocalMux
    port map (
            O => \N__57185\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13478\ : LocalMux
    port map (
            O => \N__57182\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13477\ : Odrv4
    port map (
            O => \N__57179\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13476\ : Odrv12
    port map (
            O => \N__57176\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13475\ : Odrv4
    port map (
            O => \N__57173\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13474\ : LocalMux
    port map (
            O => \N__57170\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13473\ : Odrv4
    port map (
            O => \N__57167\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\
        );

    \I__13472\ : CascadeMux
    port map (
            O => \N__57150\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0_cascade_\
        );

    \I__13471\ : CascadeMux
    port map (
            O => \N__57147\,
            I => \N__57143\
        );

    \I__13470\ : InMux
    port map (
            O => \N__57146\,
            I => \N__57138\
        );

    \I__13469\ : InMux
    port map (
            O => \N__57143\,
            I => \N__57138\
        );

    \I__13468\ : LocalMux
    port map (
            O => \N__57138\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_239\
        );

    \I__13467\ : CascadeMux
    port map (
            O => \N__57135\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_239_cascade_\
        );

    \I__13466\ : InMux
    port map (
            O => \N__57132\,
            I => \N__57128\
        );

    \I__13465\ : InMux
    port map (
            O => \N__57131\,
            I => \N__57125\
        );

    \I__13464\ : LocalMux
    port map (
            O => \N__57128\,
            I => \N__57120\
        );

    \I__13463\ : LocalMux
    port map (
            O => \N__57125\,
            I => \N__57117\
        );

    \I__13462\ : InMux
    port map (
            O => \N__57124\,
            I => \N__57114\
        );

    \I__13461\ : InMux
    port map (
            O => \N__57123\,
            I => \N__57111\
        );

    \I__13460\ : Span4Mux_h
    port map (
            O => \N__57120\,
            I => \N__57104\
        );

    \I__13459\ : Span4Mux_h
    port map (
            O => \N__57117\,
            I => \N__57104\
        );

    \I__13458\ : LocalMux
    port map (
            O => \N__57114\,
            I => \N__57104\
        );

    \I__13457\ : LocalMux
    port map (
            O => \N__57111\,
            I => \N__57101\
        );

    \I__13456\ : Span4Mux_v
    port map (
            O => \N__57104\,
            I => \N__57098\
        );

    \I__13455\ : Odrv4
    port map (
            O => \N__57101\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_294\
        );

    \I__13454\ : Odrv4
    port map (
            O => \N__57098\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_294\
        );

    \I__13453\ : CascadeMux
    port map (
            O => \N__57093\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_1_0_0_cascade_\
        );

    \I__13452\ : InMux
    port map (
            O => \N__57090\,
            I => \N__57086\
        );

    \I__13451\ : InMux
    port map (
            O => \N__57089\,
            I => \N__57083\
        );

    \I__13450\ : LocalMux
    port map (
            O => \N__57086\,
            I => \N__57079\
        );

    \I__13449\ : LocalMux
    port map (
            O => \N__57083\,
            I => \N__57076\
        );

    \I__13448\ : InMux
    port map (
            O => \N__57082\,
            I => \N__57073\
        );

    \I__13447\ : Odrv4
    port map (
            O => \N__57079\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2\
        );

    \I__13446\ : Odrv12
    port map (
            O => \N__57076\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2\
        );

    \I__13445\ : LocalMux
    port map (
            O => \N__57073\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2\
        );

    \I__13444\ : InMux
    port map (
            O => \N__57066\,
            I => \N__57063\
        );

    \I__13443\ : LocalMux
    port map (
            O => \N__57063\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_0_0\
        );

    \I__13442\ : CascadeMux
    port map (
            O => \N__57060\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446_cascade_\
        );

    \I__13441\ : CascadeMux
    port map (
            O => \N__57057\,
            I => \N__57053\
        );

    \I__13440\ : InMux
    port map (
            O => \N__57056\,
            I => \N__57050\
        );

    \I__13439\ : InMux
    port map (
            O => \N__57053\,
            I => \N__57047\
        );

    \I__13438\ : LocalMux
    port map (
            O => \N__57050\,
            I => \N__57044\
        );

    \I__13437\ : LocalMux
    port map (
            O => \N__57047\,
            I => \N__57041\
        );

    \I__13436\ : Span4Mux_v
    port map (
            O => \N__57044\,
            I => \N__57036\
        );

    \I__13435\ : Span4Mux_v
    port map (
            O => \N__57041\,
            I => \N__57036\
        );

    \I__13434\ : Span4Mux_h
    port map (
            O => \N__57036\,
            I => \N__57033\
        );

    \I__13433\ : Odrv4
    port map (
            O => \N__57033\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_291\
        );

    \I__13432\ : InMux
    port map (
            O => \N__57030\,
            I => \N__57023\
        );

    \I__13431\ : InMux
    port map (
            O => \N__57029\,
            I => \N__57023\
        );

    \I__13430\ : InMux
    port map (
            O => \N__57028\,
            I => \N__57020\
        );

    \I__13429\ : LocalMux
    port map (
            O => \N__57023\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24\
        );

    \I__13428\ : LocalMux
    port map (
            O => \N__57020\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24\
        );

    \I__13427\ : CascadeMux
    port map (
            O => \N__57015\,
            I => \N__57009\
        );

    \I__13426\ : CascadeMux
    port map (
            O => \N__57014\,
            I => \N__57006\
        );

    \I__13425\ : CascadeMux
    port map (
            O => \N__57013\,
            I => \N__57003\
        );

    \I__13424\ : InMux
    port map (
            O => \N__57012\,
            I => \N__56999\
        );

    \I__13423\ : InMux
    port map (
            O => \N__57009\,
            I => \N__56996\
        );

    \I__13422\ : InMux
    port map (
            O => \N__57006\,
            I => \N__56990\
        );

    \I__13421\ : InMux
    port map (
            O => \N__57003\,
            I => \N__56985\
        );

    \I__13420\ : InMux
    port map (
            O => \N__57002\,
            I => \N__56985\
        );

    \I__13419\ : LocalMux
    port map (
            O => \N__56999\,
            I => \N__56980\
        );

    \I__13418\ : LocalMux
    port map (
            O => \N__56996\,
            I => \N__56980\
        );

    \I__13417\ : InMux
    port map (
            O => \N__56995\,
            I => \N__56973\
        );

    \I__13416\ : InMux
    port map (
            O => \N__56994\,
            I => \N__56973\
        );

    \I__13415\ : InMux
    port map (
            O => \N__56993\,
            I => \N__56973\
        );

    \I__13414\ : LocalMux
    port map (
            O => \N__56990\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25\
        );

    \I__13413\ : LocalMux
    port map (
            O => \N__56985\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25\
        );

    \I__13412\ : Odrv4
    port map (
            O => \N__56980\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25\
        );

    \I__13411\ : LocalMux
    port map (
            O => \N__56973\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25\
        );

    \I__13410\ : InMux
    port map (
            O => \N__56964\,
            I => \N__56961\
        );

    \I__13409\ : LocalMux
    port map (
            O => \N__56961\,
            I => \N__56958\
        );

    \I__13408\ : Odrv4
    port map (
            O => \N__56958\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_0_1\
        );

    \I__13407\ : CascadeMux
    port map (
            O => \N__56955\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_232_cascade_\
        );

    \I__13406\ : CascadeMux
    port map (
            O => \N__56952\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_2_1_cascade_\
        );

    \I__13405\ : InMux
    port map (
            O => \N__56949\,
            I => \N__56943\
        );

    \I__13404\ : InMux
    port map (
            O => \N__56948\,
            I => \N__56940\
        );

    \I__13403\ : InMux
    port map (
            O => \N__56947\,
            I => \N__56935\
        );

    \I__13402\ : InMux
    port map (
            O => \N__56946\,
            I => \N__56935\
        );

    \I__13401\ : LocalMux
    port map (
            O => \N__56943\,
            I => \N__56932\
        );

    \I__13400\ : LocalMux
    port map (
            O => \N__56940\,
            I => \N__56929\
        );

    \I__13399\ : LocalMux
    port map (
            O => \N__56935\,
            I => \N__56926\
        );

    \I__13398\ : Span4Mux_h
    port map (
            O => \N__56932\,
            I => \N__56921\
        );

    \I__13397\ : Span4Mux_h
    port map (
            O => \N__56929\,
            I => \N__56921\
        );

    \I__13396\ : Odrv12
    port map (
            O => \N__56926\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4\
        );

    \I__13395\ : Odrv4
    port map (
            O => \N__56921\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4\
        );

    \I__13394\ : InMux
    port map (
            O => \N__56916\,
            I => \N__56910\
        );

    \I__13393\ : InMux
    port map (
            O => \N__56915\,
            I => \N__56910\
        );

    \I__13392\ : LocalMux
    port map (
            O => \N__56910\,
            I => \N__56905\
        );

    \I__13391\ : InMux
    port map (
            O => \N__56909\,
            I => \N__56902\
        );

    \I__13390\ : InMux
    port map (
            O => \N__56908\,
            I => \N__56899\
        );

    \I__13389\ : Span4Mux_h
    port map (
            O => \N__56905\,
            I => \N__56896\
        );

    \I__13388\ : LocalMux
    port map (
            O => \N__56902\,
            I => \N__56889\
        );

    \I__13387\ : LocalMux
    port map (
            O => \N__56899\,
            I => \N__56889\
        );

    \I__13386\ : Span4Mux_v
    port map (
            O => \N__56896\,
            I => \N__56889\
        );

    \I__13385\ : Odrv4
    port map (
            O => \N__56889\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_20\
        );

    \I__13384\ : InMux
    port map (
            O => \N__56886\,
            I => \N__56882\
        );

    \I__13383\ : InMux
    port map (
            O => \N__56885\,
            I => \N__56879\
        );

    \I__13382\ : LocalMux
    port map (
            O => \N__56882\,
            I => \N__56873\
        );

    \I__13381\ : LocalMux
    port map (
            O => \N__56879\,
            I => \N__56873\
        );

    \I__13380\ : InMux
    port map (
            O => \N__56878\,
            I => \N__56870\
        );

    \I__13379\ : Span12Mux_h
    port map (
            O => \N__56873\,
            I => \N__56863\
        );

    \I__13378\ : LocalMux
    port map (
            O => \N__56870\,
            I => \N__56863\
        );

    \I__13377\ : InMux
    port map (
            O => \N__56869\,
            I => \N__56858\
        );

    \I__13376\ : InMux
    port map (
            O => \N__56868\,
            I => \N__56858\
        );

    \I__13375\ : Odrv12
    port map (
            O => \N__56863\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12\
        );

    \I__13374\ : LocalMux
    port map (
            O => \N__56858\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12\
        );

    \I__13373\ : InMux
    port map (
            O => \N__56853\,
            I => \N__56850\
        );

    \I__13372\ : LocalMux
    port map (
            O => \N__56850\,
            I => \N__56847\
        );

    \I__13371\ : Odrv4
    port map (
            O => \N__56847\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_4_0\
        );

    \I__13370\ : CascadeMux
    port map (
            O => \N__56844\,
            I => \N__56840\
        );

    \I__13369\ : InMux
    port map (
            O => \N__56843\,
            I => \N__56837\
        );

    \I__13368\ : InMux
    port map (
            O => \N__56840\,
            I => \N__56834\
        );

    \I__13367\ : LocalMux
    port map (
            O => \N__56837\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_232\
        );

    \I__13366\ : LocalMux
    port map (
            O => \N__56834\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_232\
        );

    \I__13365\ : InMux
    port map (
            O => \N__56829\,
            I => \N__56825\
        );

    \I__13364\ : InMux
    port map (
            O => \N__56828\,
            I => \N__56822\
        );

    \I__13363\ : LocalMux
    port map (
            O => \N__56825\,
            I => \N__56819\
        );

    \I__13362\ : LocalMux
    port map (
            O => \N__56822\,
            I => \N__56812\
        );

    \I__13361\ : Span4Mux_h
    port map (
            O => \N__56819\,
            I => \N__56809\
        );

    \I__13360\ : InMux
    port map (
            O => \N__56818\,
            I => \N__56806\
        );

    \I__13359\ : InMux
    port map (
            O => \N__56817\,
            I => \N__56799\
        );

    \I__13358\ : InMux
    port map (
            O => \N__56816\,
            I => \N__56799\
        );

    \I__13357\ : InMux
    port map (
            O => \N__56815\,
            I => \N__56799\
        );

    \I__13356\ : Span4Mux_h
    port map (
            O => \N__56812\,
            I => \N__56796\
        );

    \I__13355\ : Odrv4
    port map (
            O => \N__56809\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22\
        );

    \I__13354\ : LocalMux
    port map (
            O => \N__56806\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22\
        );

    \I__13353\ : LocalMux
    port map (
            O => \N__56799\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22\
        );

    \I__13352\ : Odrv4
    port map (
            O => \N__56796\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22\
        );

    \I__13351\ : InMux
    port map (
            O => \N__56787\,
            I => \N__56784\
        );

    \I__13350\ : LocalMux
    port map (
            O => \N__56784\,
            I => \N__56781\
        );

    \I__13349\ : Odrv12
    port map (
            O => \N__56781\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_1_0\
        );

    \I__13348\ : CascadeMux
    port map (
            O => \N__56778\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_2_0_cascade_\
        );

    \I__13347\ : InMux
    port map (
            O => \N__56775\,
            I => \N__56772\
        );

    \I__13346\ : LocalMux
    port map (
            O => \N__56772\,
            I => \N__56767\
        );

    \I__13345\ : InMux
    port map (
            O => \N__56771\,
            I => \N__56762\
        );

    \I__13344\ : InMux
    port map (
            O => \N__56770\,
            I => \N__56762\
        );

    \I__13343\ : Odrv4
    port map (
            O => \N__56767\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_231\
        );

    \I__13342\ : LocalMux
    port map (
            O => \N__56762\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_231\
        );

    \I__13341\ : CascadeMux
    port map (
            O => \N__56757\,
            I => \N__56754\
        );

    \I__13340\ : InMux
    port map (
            O => \N__56754\,
            I => \N__56751\
        );

    \I__13339\ : LocalMux
    port map (
            O => \N__56751\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_212\
        );

    \I__13338\ : InMux
    port map (
            O => \N__56748\,
            I => \N__56745\
        );

    \I__13337\ : LocalMux
    port map (
            O => \N__56745\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_288\
        );

    \I__13336\ : CascadeMux
    port map (
            O => \N__56742\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_288_cascade_\
        );

    \I__13335\ : InMux
    port map (
            O => \N__56739\,
            I => \N__56736\
        );

    \I__13334\ : LocalMux
    port map (
            O => \N__56736\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_23\
        );

    \I__13333\ : InMux
    port map (
            O => \N__56733\,
            I => \N__56730\
        );

    \I__13332\ : LocalMux
    port map (
            O => \N__56730\,
            I => \N__56722\
        );

    \I__13331\ : InMux
    port map (
            O => \N__56729\,
            I => \N__56719\
        );

    \I__13330\ : InMux
    port map (
            O => \N__56728\,
            I => \N__56713\
        );

    \I__13329\ : InMux
    port map (
            O => \N__56727\,
            I => \N__56713\
        );

    \I__13328\ : InMux
    port map (
            O => \N__56726\,
            I => \N__56708\
        );

    \I__13327\ : InMux
    port map (
            O => \N__56725\,
            I => \N__56708\
        );

    \I__13326\ : Span4Mux_v
    port map (
            O => \N__56722\,
            I => \N__56705\
        );

    \I__13325\ : LocalMux
    port map (
            O => \N__56719\,
            I => \N__56702\
        );

    \I__13324\ : InMux
    port map (
            O => \N__56718\,
            I => \N__56697\
        );

    \I__13323\ : LocalMux
    port map (
            O => \N__56713\,
            I => \N__56692\
        );

    \I__13322\ : LocalMux
    port map (
            O => \N__56708\,
            I => \N__56692\
        );

    \I__13321\ : Span4Mux_h
    port map (
            O => \N__56705\,
            I => \N__56687\
        );

    \I__13320\ : Span4Mux_h
    port map (
            O => \N__56702\,
            I => \N__56687\
        );

    \I__13319\ : InMux
    port map (
            O => \N__56701\,
            I => \N__56684\
        );

    \I__13318\ : InMux
    port map (
            O => \N__56700\,
            I => \N__56681\
        );

    \I__13317\ : LocalMux
    port map (
            O => \N__56697\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\
        );

    \I__13316\ : Odrv4
    port map (
            O => \N__56692\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\
        );

    \I__13315\ : Odrv4
    port map (
            O => \N__56687\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\
        );

    \I__13314\ : LocalMux
    port map (
            O => \N__56684\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\
        );

    \I__13313\ : LocalMux
    port map (
            O => \N__56681\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\
        );

    \I__13312\ : InMux
    port map (
            O => \N__56670\,
            I => \N__56667\
        );

    \I__13311\ : LocalMux
    port map (
            O => \N__56667\,
            I => \N__56664\
        );

    \I__13310\ : Odrv4
    port map (
            O => \N__56664\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_115\
        );

    \I__13309\ : InMux
    port map (
            O => \N__56661\,
            I => \N__56657\
        );

    \I__13308\ : InMux
    port map (
            O => \N__56660\,
            I => \N__56654\
        );

    \I__13307\ : LocalMux
    port map (
            O => \N__56657\,
            I => \N__56651\
        );

    \I__13306\ : LocalMux
    port map (
            O => \N__56654\,
            I => \N__56646\
        );

    \I__13305\ : Span4Mux_h
    port map (
            O => \N__56651\,
            I => \N__56643\
        );

    \I__13304\ : InMux
    port map (
            O => \N__56650\,
            I => \N__56638\
        );

    \I__13303\ : InMux
    port map (
            O => \N__56649\,
            I => \N__56638\
        );

    \I__13302\ : Odrv4
    port map (
            O => \N__56646\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16\
        );

    \I__13301\ : Odrv4
    port map (
            O => \N__56643\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16\
        );

    \I__13300\ : LocalMux
    port map (
            O => \N__56638\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16\
        );

    \I__13299\ : CascadeMux
    port map (
            O => \N__56631\,
            I => \N__56628\
        );

    \I__13298\ : InMux
    port map (
            O => \N__56628\,
            I => \N__56622\
        );

    \I__13297\ : InMux
    port map (
            O => \N__56627\,
            I => \N__56622\
        );

    \I__13296\ : LocalMux
    port map (
            O => \N__56622\,
            I => \N__56617\
        );

    \I__13295\ : InMux
    port map (
            O => \N__56621\,
            I => \N__56612\
        );

    \I__13294\ : InMux
    port map (
            O => \N__56620\,
            I => \N__56612\
        );

    \I__13293\ : Odrv4
    port map (
            O => \N__56617\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2\
        );

    \I__13292\ : LocalMux
    port map (
            O => \N__56612\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2\
        );

    \I__13291\ : InMux
    port map (
            O => \N__56607\,
            I => \N__56601\
        );

    \I__13290\ : InMux
    port map (
            O => \N__56606\,
            I => \N__56601\
        );

    \I__13289\ : LocalMux
    port map (
            O => \N__56601\,
            I => \N__56598\
        );

    \I__13288\ : Span4Mux_h
    port map (
            O => \N__56598\,
            I => \N__56595\
        );

    \I__13287\ : Span4Mux_v
    port map (
            O => \N__56595\,
            I => \N__56588\
        );

    \I__13286\ : InMux
    port map (
            O => \N__56594\,
            I => \N__56585\
        );

    \I__13285\ : InMux
    port map (
            O => \N__56593\,
            I => \N__56578\
        );

    \I__13284\ : InMux
    port map (
            O => \N__56592\,
            I => \N__56578\
        );

    \I__13283\ : CascadeMux
    port map (
            O => \N__56591\,
            I => \N__56575\
        );

    \I__13282\ : Span4Mux_v
    port map (
            O => \N__56588\,
            I => \N__56569\
        );

    \I__13281\ : LocalMux
    port map (
            O => \N__56585\,
            I => \N__56569\
        );

    \I__13280\ : InMux
    port map (
            O => \N__56584\,
            I => \N__56564\
        );

    \I__13279\ : InMux
    port map (
            O => \N__56583\,
            I => \N__56564\
        );

    \I__13278\ : LocalMux
    port map (
            O => \N__56578\,
            I => \N__56561\
        );

    \I__13277\ : InMux
    port map (
            O => \N__56575\,
            I => \N__56554\
        );

    \I__13276\ : InMux
    port map (
            O => \N__56574\,
            I => \N__56554\
        );

    \I__13275\ : Span4Mux_v
    port map (
            O => \N__56569\,
            I => \N__56549\
        );

    \I__13274\ : LocalMux
    port map (
            O => \N__56564\,
            I => \N__56549\
        );

    \I__13273\ : Span4Mux_h
    port map (
            O => \N__56561\,
            I => \N__56546\
        );

    \I__13272\ : InMux
    port map (
            O => \N__56560\,
            I => \N__56543\
        );

    \I__13271\ : InMux
    port map (
            O => \N__56559\,
            I => \N__56540\
        );

    \I__13270\ : LocalMux
    port map (
            O => \N__56554\,
            I => \N__56537\
        );

    \I__13269\ : Span4Mux_h
    port map (
            O => \N__56549\,
            I => \N__56534\
        );

    \I__13268\ : Span4Mux_h
    port map (
            O => \N__56546\,
            I => \N__56529\
        );

    \I__13267\ : LocalMux
    port map (
            O => \N__56543\,
            I => \N__56529\
        );

    \I__13266\ : LocalMux
    port map (
            O => \N__56540\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1\
        );

    \I__13265\ : Odrv4
    port map (
            O => \N__56537\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1\
        );

    \I__13264\ : Odrv4
    port map (
            O => \N__56534\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1\
        );

    \I__13263\ : Odrv4
    port map (
            O => \N__56529\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1\
        );

    \I__13262\ : CascadeMux
    port map (
            O => \N__56520\,
            I => \N__56517\
        );

    \I__13261\ : InMux
    port map (
            O => \N__56517\,
            I => \N__56513\
        );

    \I__13260\ : InMux
    port map (
            O => \N__56516\,
            I => \N__56508\
        );

    \I__13259\ : LocalMux
    port map (
            O => \N__56513\,
            I => \N__56505\
        );

    \I__13258\ : InMux
    port map (
            O => \N__56512\,
            I => \N__56500\
        );

    \I__13257\ : InMux
    port map (
            O => \N__56511\,
            I => \N__56500\
        );

    \I__13256\ : LocalMux
    port map (
            O => \N__56508\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_904\
        );

    \I__13255\ : Odrv4
    port map (
            O => \N__56505\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_904\
        );

    \I__13254\ : LocalMux
    port map (
            O => \N__56500\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_904\
        );

    \I__13253\ : CascadeMux
    port map (
            O => \N__56493\,
            I => \N__56490\
        );

    \I__13252\ : InMux
    port map (
            O => \N__56490\,
            I => \N__56486\
        );

    \I__13251\ : InMux
    port map (
            O => \N__56489\,
            I => \N__56483\
        );

    \I__13250\ : LocalMux
    port map (
            O => \N__56486\,
            I => \N__56480\
        );

    \I__13249\ : LocalMux
    port map (
            O => \N__56483\,
            I => \N__56477\
        );

    \I__13248\ : Span4Mux_h
    port map (
            O => \N__56480\,
            I => \N__56472\
        );

    \I__13247\ : Span4Mux_h
    port map (
            O => \N__56477\,
            I => \N__56472\
        );

    \I__13246\ : Odrv4
    port map (
            O => \N__56472\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_2\
        );

    \I__13245\ : InMux
    port map (
            O => \N__56469\,
            I => \N__56465\
        );

    \I__13244\ : InMux
    port map (
            O => \N__56468\,
            I => \N__56462\
        );

    \I__13243\ : LocalMux
    port map (
            O => \N__56465\,
            I => \N__56459\
        );

    \I__13242\ : LocalMux
    port map (
            O => \N__56462\,
            I => \N__56456\
        );

    \I__13241\ : Span4Mux_v
    port map (
            O => \N__56459\,
            I => \N__56453\
        );

    \I__13240\ : Odrv4
    port map (
            O => \N__56456\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1\
        );

    \I__13239\ : Odrv4
    port map (
            O => \N__56453\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1\
        );

    \I__13238\ : InMux
    port map (
            O => \N__56448\,
            I => \N__56443\
        );

    \I__13237\ : InMux
    port map (
            O => \N__56447\,
            I => \N__56434\
        );

    \I__13236\ : InMux
    port map (
            O => \N__56446\,
            I => \N__56434\
        );

    \I__13235\ : LocalMux
    port map (
            O => \N__56443\,
            I => \N__56431\
        );

    \I__13234\ : InMux
    port map (
            O => \N__56442\,
            I => \N__56428\
        );

    \I__13233\ : InMux
    port map (
            O => \N__56441\,
            I => \N__56425\
        );

    \I__13232\ : CascadeMux
    port map (
            O => \N__56440\,
            I => \N__56422\
        );

    \I__13231\ : InMux
    port map (
            O => \N__56439\,
            I => \N__56419\
        );

    \I__13230\ : LocalMux
    port map (
            O => \N__56434\,
            I => \N__56416\
        );

    \I__13229\ : Span4Mux_v
    port map (
            O => \N__56431\,
            I => \N__56411\
        );

    \I__13228\ : LocalMux
    port map (
            O => \N__56428\,
            I => \N__56411\
        );

    \I__13227\ : LocalMux
    port map (
            O => \N__56425\,
            I => \N__56408\
        );

    \I__13226\ : InMux
    port map (
            O => \N__56422\,
            I => \N__56403\
        );

    \I__13225\ : LocalMux
    port map (
            O => \N__56419\,
            I => \N__56394\
        );

    \I__13224\ : Span4Mux_v
    port map (
            O => \N__56416\,
            I => \N__56394\
        );

    \I__13223\ : Span4Mux_v
    port map (
            O => \N__56411\,
            I => \N__56394\
        );

    \I__13222\ : Span4Mux_h
    port map (
            O => \N__56408\,
            I => \N__56394\
        );

    \I__13221\ : InMux
    port map (
            O => \N__56407\,
            I => \N__56389\
        );

    \I__13220\ : InMux
    port map (
            O => \N__56406\,
            I => \N__56389\
        );

    \I__13219\ : LocalMux
    port map (
            O => \N__56403\,
            I => \N__56384\
        );

    \I__13218\ : Span4Mux_h
    port map (
            O => \N__56394\,
            I => \N__56384\
        );

    \I__13217\ : LocalMux
    port map (
            O => \N__56389\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26\
        );

    \I__13216\ : Odrv4
    port map (
            O => \N__56384\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26\
        );

    \I__13215\ : CascadeMux
    port map (
            O => \N__56379\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un30_i_a2_9_a2_4_a2_0_1_2_cascade_\
        );

    \I__13214\ : InMux
    port map (
            O => \N__56376\,
            I => \N__56373\
        );

    \I__13213\ : LocalMux
    port map (
            O => \N__56373\,
            I => \N__56370\
        );

    \I__13212\ : Span12Mux_h
    port map (
            O => \N__56370\,
            I => \N__56367\
        );

    \I__13211\ : Odrv12
    port map (
            O => \N__56367\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446\
        );

    \I__13210\ : CascadeMux
    port map (
            O => \N__56364\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0_cascade_\
        );

    \I__13209\ : InMux
    port map (
            O => \N__56361\,
            I => \N__56354\
        );

    \I__13208\ : InMux
    port map (
            O => \N__56360\,
            I => \N__56347\
        );

    \I__13207\ : InMux
    port map (
            O => \N__56359\,
            I => \N__56340\
        );

    \I__13206\ : InMux
    port map (
            O => \N__56358\,
            I => \N__56340\
        );

    \I__13205\ : InMux
    port map (
            O => \N__56357\,
            I => \N__56340\
        );

    \I__13204\ : LocalMux
    port map (
            O => \N__56354\,
            I => \N__56337\
        );

    \I__13203\ : CascadeMux
    port map (
            O => \N__56353\,
            I => \N__56333\
        );

    \I__13202\ : InMux
    port map (
            O => \N__56352\,
            I => \N__56330\
        );

    \I__13201\ : InMux
    port map (
            O => \N__56351\,
            I => \N__56327\
        );

    \I__13200\ : InMux
    port map (
            O => \N__56350\,
            I => \N__56324\
        );

    \I__13199\ : LocalMux
    port map (
            O => \N__56347\,
            I => \N__56317\
        );

    \I__13198\ : LocalMux
    port map (
            O => \N__56340\,
            I => \N__56317\
        );

    \I__13197\ : Span4Mux_h
    port map (
            O => \N__56337\,
            I => \N__56317\
        );

    \I__13196\ : InMux
    port map (
            O => \N__56336\,
            I => \N__56312\
        );

    \I__13195\ : InMux
    port map (
            O => \N__56333\,
            I => \N__56312\
        );

    \I__13194\ : LocalMux
    port map (
            O => \N__56330\,
            I => \N__56309\
        );

    \I__13193\ : LocalMux
    port map (
            O => \N__56327\,
            I => \N__56299\
        );

    \I__13192\ : LocalMux
    port map (
            O => \N__56324\,
            I => \N__56299\
        );

    \I__13191\ : Sp12to4
    port map (
            O => \N__56317\,
            I => \N__56299\
        );

    \I__13190\ : LocalMux
    port map (
            O => \N__56312\,
            I => \N__56299\
        );

    \I__13189\ : Span4Mux_v
    port map (
            O => \N__56309\,
            I => \N__56296\
        );

    \I__13188\ : InMux
    port map (
            O => \N__56308\,
            I => \N__56293\
        );

    \I__13187\ : Span12Mux_v
    port map (
            O => \N__56299\,
            I => \N__56290\
        );

    \I__13186\ : Odrv4
    port map (
            O => \N__56296\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15\
        );

    \I__13185\ : LocalMux
    port map (
            O => \N__56293\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15\
        );

    \I__13184\ : Odrv12
    port map (
            O => \N__56290\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15\
        );

    \I__13183\ : CascadeMux
    port map (
            O => \N__56283\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_5_0_cascade_\
        );

    \I__13182\ : InMux
    port map (
            O => \N__56280\,
            I => \N__56277\
        );

    \I__13181\ : LocalMux
    port map (
            O => \N__56277\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_6_0\
        );

    \I__13180\ : InMux
    port map (
            O => \N__56274\,
            I => \N__56271\
        );

    \I__13179\ : LocalMux
    port map (
            O => \N__56271\,
            I => \N__56268\
        );

    \I__13178\ : Span4Mux_h
    port map (
            O => \N__56268\,
            I => \N__56265\
        );

    \I__13177\ : Odrv4
    port map (
            O => \N__56265\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_7_0\
        );

    \I__13176\ : InMux
    port map (
            O => \N__56262\,
            I => \N__56259\
        );

    \I__13175\ : LocalMux
    port map (
            O => \N__56259\,
            I => \N__56256\
        );

    \I__13174\ : Odrv4
    port map (
            O => \N__56256\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_0\
        );

    \I__13173\ : CascadeMux
    port map (
            O => \N__56253\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_11_0_cascade_\
        );

    \I__13172\ : CascadeMux
    port map (
            O => \N__56250\,
            I => \N__56242\
        );

    \I__13171\ : InMux
    port map (
            O => \N__56249\,
            I => \N__56239\
        );

    \I__13170\ : InMux
    port map (
            O => \N__56248\,
            I => \N__56236\
        );

    \I__13169\ : InMux
    port map (
            O => \N__56247\,
            I => \N__56233\
        );

    \I__13168\ : InMux
    port map (
            O => \N__56246\,
            I => \N__56229\
        );

    \I__13167\ : CascadeMux
    port map (
            O => \N__56245\,
            I => \N__56226\
        );

    \I__13166\ : InMux
    port map (
            O => \N__56242\,
            I => \N__56223\
        );

    \I__13165\ : LocalMux
    port map (
            O => \N__56239\,
            I => \N__56216\
        );

    \I__13164\ : LocalMux
    port map (
            O => \N__56236\,
            I => \N__56216\
        );

    \I__13163\ : LocalMux
    port map (
            O => \N__56233\,
            I => \N__56216\
        );

    \I__13162\ : InMux
    port map (
            O => \N__56232\,
            I => \N__56213\
        );

    \I__13161\ : LocalMux
    port map (
            O => \N__56229\,
            I => \N__56210\
        );

    \I__13160\ : InMux
    port map (
            O => \N__56226\,
            I => \N__56207\
        );

    \I__13159\ : LocalMux
    port map (
            O => \N__56223\,
            I => \N__56204\
        );

    \I__13158\ : Span4Mux_v
    port map (
            O => \N__56216\,
            I => \N__56201\
        );

    \I__13157\ : LocalMux
    port map (
            O => \N__56213\,
            I => \N__56198\
        );

    \I__13156\ : Span4Mux_h
    port map (
            O => \N__56210\,
            I => \N__56195\
        );

    \I__13155\ : LocalMux
    port map (
            O => \N__56207\,
            I => \N__56186\
        );

    \I__13154\ : Span4Mux_v
    port map (
            O => \N__56204\,
            I => \N__56186\
        );

    \I__13153\ : Span4Mux_h
    port map (
            O => \N__56201\,
            I => \N__56186\
        );

    \I__13152\ : Span4Mux_v
    port map (
            O => \N__56198\,
            I => \N__56186\
        );

    \I__13151\ : Odrv4
    port map (
            O => \N__56195\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13\
        );

    \I__13150\ : Odrv4
    port map (
            O => \N__56186\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13\
        );

    \I__13149\ : InMux
    port map (
            O => \N__56181\,
            I => \N__56177\
        );

    \I__13148\ : InMux
    port map (
            O => \N__56180\,
            I => \N__56174\
        );

    \I__13147\ : LocalMux
    port map (
            O => \N__56177\,
            I => \N__56170\
        );

    \I__13146\ : LocalMux
    port map (
            O => \N__56174\,
            I => \N__56167\
        );

    \I__13145\ : InMux
    port map (
            O => \N__56173\,
            I => \N__56164\
        );

    \I__13144\ : Span4Mux_v
    port map (
            O => \N__56170\,
            I => \N__56159\
        );

    \I__13143\ : Span4Mux_v
    port map (
            O => \N__56167\,
            I => \N__56159\
        );

    \I__13142\ : LocalMux
    port map (
            O => \N__56164\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6\
        );

    \I__13141\ : Odrv4
    port map (
            O => \N__56159\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6\
        );

    \I__13140\ : CascadeMux
    port map (
            O => \N__56154\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_23_cascade_\
        );

    \I__13139\ : CascadeMux
    port map (
            O => \N__56151\,
            I => \N__56148\
        );

    \I__13138\ : InMux
    port map (
            O => \N__56148\,
            I => \N__56141\
        );

    \I__13137\ : InMux
    port map (
            O => \N__56147\,
            I => \N__56138\
        );

    \I__13136\ : InMux
    port map (
            O => \N__56146\,
            I => \N__56131\
        );

    \I__13135\ : InMux
    port map (
            O => \N__56145\,
            I => \N__56131\
        );

    \I__13134\ : InMux
    port map (
            O => \N__56144\,
            I => \N__56131\
        );

    \I__13133\ : LocalMux
    port map (
            O => \N__56141\,
            I => \N__56124\
        );

    \I__13132\ : LocalMux
    port map (
            O => \N__56138\,
            I => \N__56119\
        );

    \I__13131\ : LocalMux
    port map (
            O => \N__56131\,
            I => \N__56116\
        );

    \I__13130\ : InMux
    port map (
            O => \N__56130\,
            I => \N__56113\
        );

    \I__13129\ : InMux
    port map (
            O => \N__56129\,
            I => \N__56110\
        );

    \I__13128\ : InMux
    port map (
            O => \N__56128\,
            I => \N__56105\
        );

    \I__13127\ : InMux
    port map (
            O => \N__56127\,
            I => \N__56105\
        );

    \I__13126\ : Span4Mux_h
    port map (
            O => \N__56124\,
            I => \N__56102\
        );

    \I__13125\ : InMux
    port map (
            O => \N__56123\,
            I => \N__56099\
        );

    \I__13124\ : InMux
    port map (
            O => \N__56122\,
            I => \N__56096\
        );

    \I__13123\ : Span4Mux_h
    port map (
            O => \N__56119\,
            I => \N__56093\
        );

    \I__13122\ : Span4Mux_h
    port map (
            O => \N__56116\,
            I => \N__56088\
        );

    \I__13121\ : LocalMux
    port map (
            O => \N__56113\,
            I => \N__56088\
        );

    \I__13120\ : LocalMux
    port map (
            O => \N__56110\,
            I => \N__56081\
        );

    \I__13119\ : LocalMux
    port map (
            O => \N__56105\,
            I => \N__56081\
        );

    \I__13118\ : Span4Mux_h
    port map (
            O => \N__56102\,
            I => \N__56081\
        );

    \I__13117\ : LocalMux
    port map (
            O => \N__56099\,
            I => \s_paddr_I2C_8\
        );

    \I__13116\ : LocalMux
    port map (
            O => \N__56096\,
            I => \s_paddr_I2C_8\
        );

    \I__13115\ : Odrv4
    port map (
            O => \N__56093\,
            I => \s_paddr_I2C_8\
        );

    \I__13114\ : Odrv4
    port map (
            O => \N__56088\,
            I => \s_paddr_I2C_8\
        );

    \I__13113\ : Odrv4
    port map (
            O => \N__56081\,
            I => \s_paddr_I2C_8\
        );

    \I__13112\ : InMux
    port map (
            O => \N__56070\,
            I => \N__56066\
        );

    \I__13111\ : InMux
    port map (
            O => \N__56069\,
            I => \N__56063\
        );

    \I__13110\ : LocalMux
    port map (
            O => \N__56066\,
            I => \N__56058\
        );

    \I__13109\ : LocalMux
    port map (
            O => \N__56063\,
            I => \N__56058\
        );

    \I__13108\ : Span4Mux_h
    port map (
            O => \N__56058\,
            I => \N__56053\
        );

    \I__13107\ : InMux
    port map (
            O => \N__56057\,
            I => \N__56050\
        );

    \I__13106\ : InMux
    port map (
            O => \N__56056\,
            I => \N__56047\
        );

    \I__13105\ : Odrv4
    port map (
            O => \N__56053\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0\
        );

    \I__13104\ : LocalMux
    port map (
            O => \N__56050\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0\
        );

    \I__13103\ : LocalMux
    port map (
            O => \N__56047\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0\
        );

    \I__13102\ : CascadeMux
    port map (
            O => \N__56040\,
            I => \N__56037\
        );

    \I__13101\ : InMux
    port map (
            O => \N__56037\,
            I => \N__56031\
        );

    \I__13100\ : InMux
    port map (
            O => \N__56036\,
            I => \N__56031\
        );

    \I__13099\ : LocalMux
    port map (
            O => \N__56031\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_230\
        );

    \I__13098\ : InMux
    port map (
            O => \N__56028\,
            I => \N__56022\
        );

    \I__13097\ : InMux
    port map (
            O => \N__56027\,
            I => \N__56022\
        );

    \I__13096\ : LocalMux
    port map (
            O => \N__56022\,
            I => \N__56019\
        );

    \I__13095\ : Span4Mux_v
    port map (
            O => \N__56019\,
            I => \N__56016\
        );

    \I__13094\ : Odrv4
    port map (
            O => \N__56016\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0\
        );

    \I__13093\ : CascadeMux
    port map (
            O => \N__56013\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0_cascade_\
        );

    \I__13092\ : InMux
    port map (
            O => \N__56010\,
            I => \N__56007\
        );

    \I__13091\ : LocalMux
    port map (
            O => \N__56007\,
            I => \N__56004\
        );

    \I__13090\ : Span4Mux_h
    port map (
            O => \N__56004\,
            I => \N__56001\
        );

    \I__13089\ : Odrv4
    port map (
            O => \N__56001\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_4\
        );

    \I__13088\ : CascadeMux
    port map (
            O => \N__55998\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_365_0_cascade_\
        );

    \I__13087\ : CascadeMux
    port map (
            O => \N__55995\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_4_0_a2_2_cascade_\
        );

    \I__13086\ : CascadeMux
    port map (
            O => \N__55992\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_676_0_cascade_\
        );

    \I__13085\ : InMux
    port map (
            O => \N__55989\,
            I => \N__55983\
        );

    \I__13084\ : InMux
    port map (
            O => \N__55988\,
            I => \N__55983\
        );

    \I__13083\ : LocalMux
    port map (
            O => \N__55983\,
            I => \N__55979\
        );

    \I__13082\ : InMux
    port map (
            O => \N__55982\,
            I => \N__55976\
        );

    \I__13081\ : Span4Mux_v
    port map (
            O => \N__55979\,
            I => \N__55971\
        );

    \I__13080\ : LocalMux
    port map (
            O => \N__55976\,
            I => \N__55971\
        );

    \I__13079\ : Odrv4
    port map (
            O => \N__55971\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address\
        );

    \I__13078\ : InMux
    port map (
            O => \N__55968\,
            I => \N__55965\
        );

    \I__13077\ : LocalMux
    port map (
            O => \N__55965\,
            I => \N__55961\
        );

    \I__13076\ : InMux
    port map (
            O => \N__55964\,
            I => \N__55957\
        );

    \I__13075\ : Span4Mux_v
    port map (
            O => \N__55961\,
            I => \N__55954\
        );

    \I__13074\ : InMux
    port map (
            O => \N__55960\,
            I => \N__55951\
        );

    \I__13073\ : LocalMux
    port map (
            O => \N__55957\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1\
        );

    \I__13072\ : Odrv4
    port map (
            O => \N__55954\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1\
        );

    \I__13071\ : LocalMux
    port map (
            O => \N__55951\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1\
        );

    \I__13070\ : CascadeMux
    port map (
            O => \N__55944\,
            I => \N__55940\
        );

    \I__13069\ : InMux
    port map (
            O => \N__55943\,
            I => \N__55937\
        );

    \I__13068\ : InMux
    port map (
            O => \N__55940\,
            I => \N__55934\
        );

    \I__13067\ : LocalMux
    port map (
            O => \N__55937\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3\
        );

    \I__13066\ : LocalMux
    port map (
            O => \N__55934\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3\
        );

    \I__13065\ : InMux
    port map (
            O => \N__55929\,
            I => \N__55924\
        );

    \I__13064\ : InMux
    port map (
            O => \N__55928\,
            I => \N__55921\
        );

    \I__13063\ : InMux
    port map (
            O => \N__55927\,
            I => \N__55917\
        );

    \I__13062\ : LocalMux
    port map (
            O => \N__55924\,
            I => \N__55913\
        );

    \I__13061\ : LocalMux
    port map (
            O => \N__55921\,
            I => \N__55910\
        );

    \I__13060\ : InMux
    port map (
            O => \N__55920\,
            I => \N__55907\
        );

    \I__13059\ : LocalMux
    port map (
            O => \N__55917\,
            I => \N__55904\
        );

    \I__13058\ : InMux
    port map (
            O => \N__55916\,
            I => \N__55901\
        );

    \I__13057\ : Span4Mux_h
    port map (
            O => \N__55913\,
            I => \N__55896\
        );

    \I__13056\ : Span4Mux_v
    port map (
            O => \N__55910\,
            I => \N__55896\
        );

    \I__13055\ : LocalMux
    port map (
            O => \N__55907\,
            I => \N__55893\
        );

    \I__13054\ : Span12Mux_v
    port map (
            O => \N__55904\,
            I => \N__55890\
        );

    \I__13053\ : LocalMux
    port map (
            O => \N__55901\,
            I => \N__55887\
        );

    \I__13052\ : Span4Mux_v
    port map (
            O => \N__55896\,
            I => \N__55884\
        );

    \I__13051\ : Odrv4
    port map (
            O => \N__55893\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16\
        );

    \I__13050\ : Odrv12
    port map (
            O => \N__55890\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16\
        );

    \I__13049\ : Odrv12
    port map (
            O => \N__55887\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16\
        );

    \I__13048\ : Odrv4
    port map (
            O => \N__55884\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16\
        );

    \I__13047\ : InMux
    port map (
            O => \N__55875\,
            I => \N__55872\
        );

    \I__13046\ : LocalMux
    port map (
            O => \N__55872\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_1\
        );

    \I__13045\ : InMux
    port map (
            O => \N__55869\,
            I => \N__55865\
        );

    \I__13044\ : InMux
    port map (
            O => \N__55868\,
            I => \N__55858\
        );

    \I__13043\ : LocalMux
    port map (
            O => \N__55865\,
            I => \N__55850\
        );

    \I__13042\ : InMux
    port map (
            O => \N__55864\,
            I => \N__55847\
        );

    \I__13041\ : InMux
    port map (
            O => \N__55863\,
            I => \N__55844\
        );

    \I__13040\ : InMux
    port map (
            O => \N__55862\,
            I => \N__55841\
        );

    \I__13039\ : InMux
    port map (
            O => \N__55861\,
            I => \N__55838\
        );

    \I__13038\ : LocalMux
    port map (
            O => \N__55858\,
            I => \N__55835\
        );

    \I__13037\ : InMux
    port map (
            O => \N__55857\,
            I => \N__55824\
        );

    \I__13036\ : InMux
    port map (
            O => \N__55856\,
            I => \N__55824\
        );

    \I__13035\ : InMux
    port map (
            O => \N__55855\,
            I => \N__55824\
        );

    \I__13034\ : InMux
    port map (
            O => \N__55854\,
            I => \N__55824\
        );

    \I__13033\ : InMux
    port map (
            O => \N__55853\,
            I => \N__55824\
        );

    \I__13032\ : Span4Mux_h
    port map (
            O => \N__55850\,
            I => \N__55817\
        );

    \I__13031\ : LocalMux
    port map (
            O => \N__55847\,
            I => \N__55817\
        );

    \I__13030\ : LocalMux
    port map (
            O => \N__55844\,
            I => \N__55817\
        );

    \I__13029\ : LocalMux
    port map (
            O => \N__55841\,
            I => \N__55808\
        );

    \I__13028\ : LocalMux
    port map (
            O => \N__55838\,
            I => \N__55808\
        );

    \I__13027\ : Span4Mux_v
    port map (
            O => \N__55835\,
            I => \N__55808\
        );

    \I__13026\ : LocalMux
    port map (
            O => \N__55824\,
            I => \N__55808\
        );

    \I__13025\ : Span4Mux_v
    port map (
            O => \N__55817\,
            I => \N__55805\
        );

    \I__13024\ : Odrv4
    port map (
            O => \N__55808\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0\
        );

    \I__13023\ : Odrv4
    port map (
            O => \N__55805\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0\
        );

    \I__13022\ : InMux
    port map (
            O => \N__55800\,
            I => \N__55797\
        );

    \I__13021\ : LocalMux
    port map (
            O => \N__55797\,
            I => \N__55791\
        );

    \I__13020\ : InMux
    port map (
            O => \N__55796\,
            I => \N__55788\
        );

    \I__13019\ : InMux
    port map (
            O => \N__55795\,
            I => \N__55785\
        );

    \I__13018\ : InMux
    port map (
            O => \N__55794\,
            I => \N__55782\
        );

    \I__13017\ : Span4Mux_v
    port map (
            O => \N__55791\,
            I => \N__55775\
        );

    \I__13016\ : LocalMux
    port map (
            O => \N__55788\,
            I => \N__55775\
        );

    \I__13015\ : LocalMux
    port map (
            O => \N__55785\,
            I => \N__55775\
        );

    \I__13014\ : LocalMux
    port map (
            O => \N__55782\,
            I => \N__55770\
        );

    \I__13013\ : Span4Mux_h
    port map (
            O => \N__55775\,
            I => \N__55770\
        );

    \I__13012\ : Odrv4
    port map (
            O => \N__55770\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1606_0\
        );

    \I__13011\ : InMux
    port map (
            O => \N__55767\,
            I => \N__55764\
        );

    \I__13010\ : LocalMux
    port map (
            O => \N__55764\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1565_0\
        );

    \I__13009\ : InMux
    port map (
            O => \N__55761\,
            I => \N__55758\
        );

    \I__13008\ : LocalMux
    port map (
            O => \N__55758\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0\
        );

    \I__13007\ : CascadeMux
    port map (
            O => \N__55755\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RLZ0Z7_cascade_\
        );

    \I__13006\ : InMux
    port map (
            O => \N__55752\,
            I => \N__55749\
        );

    \I__13005\ : LocalMux
    port map (
            O => \N__55749\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2\
        );

    \I__13004\ : InMux
    port map (
            O => \N__55746\,
            I => \N__55735\
        );

    \I__13003\ : InMux
    port map (
            O => \N__55745\,
            I => \N__55735\
        );

    \I__13002\ : InMux
    port map (
            O => \N__55744\,
            I => \N__55728\
        );

    \I__13001\ : InMux
    port map (
            O => \N__55743\,
            I => \N__55728\
        );

    \I__13000\ : InMux
    port map (
            O => \N__55742\,
            I => \N__55728\
        );

    \I__12999\ : InMux
    port map (
            O => \N__55741\,
            I => \N__55717\
        );

    \I__12998\ : InMux
    port map (
            O => \N__55740\,
            I => \N__55717\
        );

    \I__12997\ : LocalMux
    port map (
            O => \N__55735\,
            I => \N__55712\
        );

    \I__12996\ : LocalMux
    port map (
            O => \N__55728\,
            I => \N__55712\
        );

    \I__12995\ : InMux
    port map (
            O => \N__55727\,
            I => \N__55707\
        );

    \I__12994\ : InMux
    port map (
            O => \N__55726\,
            I => \N__55707\
        );

    \I__12993\ : InMux
    port map (
            O => \N__55725\,
            I => \N__55702\
        );

    \I__12992\ : InMux
    port map (
            O => \N__55724\,
            I => \N__55702\
        );

    \I__12991\ : InMux
    port map (
            O => \N__55723\,
            I => \N__55697\
        );

    \I__12990\ : InMux
    port map (
            O => \N__55722\,
            I => \N__55697\
        );

    \I__12989\ : LocalMux
    port map (
            O => \N__55717\,
            I => \N__55690\
        );

    \I__12988\ : Span4Mux_v
    port map (
            O => \N__55712\,
            I => \N__55683\
        );

    \I__12987\ : LocalMux
    port map (
            O => \N__55707\,
            I => \N__55680\
        );

    \I__12986\ : LocalMux
    port map (
            O => \N__55702\,
            I => \N__55675\
        );

    \I__12985\ : LocalMux
    port map (
            O => \N__55697\,
            I => \N__55675\
        );

    \I__12984\ : InMux
    port map (
            O => \N__55696\,
            I => \N__55670\
        );

    \I__12983\ : InMux
    port map (
            O => \N__55695\,
            I => \N__55670\
        );

    \I__12982\ : InMux
    port map (
            O => \N__55694\,
            I => \N__55665\
        );

    \I__12981\ : InMux
    port map (
            O => \N__55693\,
            I => \N__55665\
        );

    \I__12980\ : Span4Mux_h
    port map (
            O => \N__55690\,
            I => \N__55662\
        );

    \I__12979\ : InMux
    port map (
            O => \N__55689\,
            I => \N__55653\
        );

    \I__12978\ : InMux
    port map (
            O => \N__55688\,
            I => \N__55653\
        );

    \I__12977\ : InMux
    port map (
            O => \N__55687\,
            I => \N__55653\
        );

    \I__12976\ : InMux
    port map (
            O => \N__55686\,
            I => \N__55653\
        );

    \I__12975\ : Span4Mux_v
    port map (
            O => \N__55683\,
            I => \N__55645\
        );

    \I__12974\ : Span4Mux_v
    port map (
            O => \N__55680\,
            I => \N__55645\
        );

    \I__12973\ : Span4Mux_v
    port map (
            O => \N__55675\,
            I => \N__55640\
        );

    \I__12972\ : LocalMux
    port map (
            O => \N__55670\,
            I => \N__55640\
        );

    \I__12971\ : LocalMux
    port map (
            O => \N__55665\,
            I => \N__55637\
        );

    \I__12970\ : Span4Mux_h
    port map (
            O => \N__55662\,
            I => \N__55632\
        );

    \I__12969\ : LocalMux
    port map (
            O => \N__55653\,
            I => \N__55632\
        );

    \I__12968\ : InMux
    port map (
            O => \N__55652\,
            I => \N__55625\
        );

    \I__12967\ : InMux
    port map (
            O => \N__55651\,
            I => \N__55625\
        );

    \I__12966\ : InMux
    port map (
            O => \N__55650\,
            I => \N__55625\
        );

    \I__12965\ : Span4Mux_h
    port map (
            O => \N__55645\,
            I => \N__55622\
        );

    \I__12964\ : Span4Mux_h
    port map (
            O => \N__55640\,
            I => \N__55619\
        );

    \I__12963\ : Span4Mux_v
    port map (
            O => \N__55637\,
            I => \N__55612\
        );

    \I__12962\ : Span4Mux_h
    port map (
            O => \N__55632\,
            I => \N__55612\
        );

    \I__12961\ : LocalMux
    port map (
            O => \N__55625\,
            I => \N__55612\
        );

    \I__12960\ : Span4Mux_h
    port map (
            O => \N__55622\,
            I => \N__55609\
        );

    \I__12959\ : Span4Mux_h
    port map (
            O => \N__55619\,
            I => \N__55606\
        );

    \I__12958\ : Span4Mux_h
    port map (
            O => \N__55612\,
            I => \N__55603\
        );

    \I__12957\ : Odrv4
    port map (
            O => \N__55609\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3\
        );

    \I__12956\ : Odrv4
    port map (
            O => \N__55606\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3\
        );

    \I__12955\ : Odrv4
    port map (
            O => \N__55603\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3\
        );

    \I__12954\ : CascadeMux
    port map (
            O => \N__55596\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2_cascade_\
        );

    \I__12953\ : InMux
    port map (
            O => \N__55593\,
            I => \N__55590\
        );

    \I__12952\ : LocalMux
    port map (
            O => \N__55590\,
            I => \N__55587\
        );

    \I__12951\ : Odrv4
    port map (
            O => \N__55587\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_1\
        );

    \I__12950\ : InMux
    port map (
            O => \N__55584\,
            I => \N__55581\
        );

    \I__12949\ : LocalMux
    port map (
            O => \N__55581\,
            I => \N__55578\
        );

    \I__12948\ : Span12Mux_h
    port map (
            O => \N__55578\,
            I => \N__55575\
        );

    \I__12947\ : Odrv12
    port map (
            O => \N__55575\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_2\
        );

    \I__12946\ : CEMux
    port map (
            O => \N__55572\,
            I => \N__55567\
        );

    \I__12945\ : CEMux
    port map (
            O => \N__55571\,
            I => \N__55564\
        );

    \I__12944\ : CEMux
    port map (
            O => \N__55570\,
            I => \N__55560\
        );

    \I__12943\ : LocalMux
    port map (
            O => \N__55567\,
            I => \N__55555\
        );

    \I__12942\ : LocalMux
    port map (
            O => \N__55564\,
            I => \N__55552\
        );

    \I__12941\ : CEMux
    port map (
            O => \N__55563\,
            I => \N__55549\
        );

    \I__12940\ : LocalMux
    port map (
            O => \N__55560\,
            I => \N__55546\
        );

    \I__12939\ : CEMux
    port map (
            O => \N__55559\,
            I => \N__55543\
        );

    \I__12938\ : CEMux
    port map (
            O => \N__55558\,
            I => \N__55540\
        );

    \I__12937\ : Span4Mux_h
    port map (
            O => \N__55555\,
            I => \N__55531\
        );

    \I__12936\ : Span4Mux_v
    port map (
            O => \N__55552\,
            I => \N__55531\
        );

    \I__12935\ : LocalMux
    port map (
            O => \N__55549\,
            I => \N__55531\
        );

    \I__12934\ : Span4Mux_h
    port map (
            O => \N__55546\,
            I => \N__55526\
        );

    \I__12933\ : LocalMux
    port map (
            O => \N__55543\,
            I => \N__55526\
        );

    \I__12932\ : LocalMux
    port map (
            O => \N__55540\,
            I => \N__55523\
        );

    \I__12931\ : CEMux
    port map (
            O => \N__55539\,
            I => \N__55518\
        );

    \I__12930\ : CEMux
    port map (
            O => \N__55538\,
            I => \N__55515\
        );

    \I__12929\ : Span4Mux_h
    port map (
            O => \N__55531\,
            I => \N__55512\
        );

    \I__12928\ : Span4Mux_h
    port map (
            O => \N__55526\,
            I => \N__55507\
        );

    \I__12927\ : Span4Mux_h
    port map (
            O => \N__55523\,
            I => \N__55507\
        );

    \I__12926\ : CEMux
    port map (
            O => \N__55522\,
            I => \N__55504\
        );

    \I__12925\ : CEMux
    port map (
            O => \N__55521\,
            I => \N__55501\
        );

    \I__12924\ : LocalMux
    port map (
            O => \N__55518\,
            I => \N__55498\
        );

    \I__12923\ : LocalMux
    port map (
            O => \N__55515\,
            I => \N__55495\
        );

    \I__12922\ : Span4Mux_h
    port map (
            O => \N__55512\,
            I => \N__55492\
        );

    \I__12921\ : Span4Mux_h
    port map (
            O => \N__55507\,
            I => \N__55489\
        );

    \I__12920\ : LocalMux
    port map (
            O => \N__55504\,
            I => \N__55484\
        );

    \I__12919\ : LocalMux
    port map (
            O => \N__55501\,
            I => \N__55484\
        );

    \I__12918\ : Span4Mux_v
    port map (
            O => \N__55498\,
            I => \N__55481\
        );

    \I__12917\ : Span4Mux_v
    port map (
            O => \N__55495\,
            I => \N__55478\
        );

    \I__12916\ : Sp12to4
    port map (
            O => \N__55492\,
            I => \N__55475\
        );

    \I__12915\ : Sp12to4
    port map (
            O => \N__55489\,
            I => \N__55472\
        );

    \I__12914\ : Span4Mux_v
    port map (
            O => \N__55484\,
            I => \N__55467\
        );

    \I__12913\ : Span4Mux_h
    port map (
            O => \N__55481\,
            I => \N__55467\
        );

    \I__12912\ : Sp12to4
    port map (
            O => \N__55478\,
            I => \N__55460\
        );

    \I__12911\ : Span12Mux_v
    port map (
            O => \N__55475\,
            I => \N__55460\
        );

    \I__12910\ : Span12Mux_v
    port map (
            O => \N__55472\,
            I => \N__55460\
        );

    \I__12909\ : Odrv4
    port map (
            O => \N__55467\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i\
        );

    \I__12908\ : Odrv12
    port map (
            O => \N__55460\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i\
        );

    \I__12907\ : InMux
    port map (
            O => \N__55455\,
            I => \N__55439\
        );

    \I__12906\ : InMux
    port map (
            O => \N__55454\,
            I => \N__55439\
        );

    \I__12905\ : InMux
    port map (
            O => \N__55453\,
            I => \N__55435\
        );

    \I__12904\ : InMux
    port map (
            O => \N__55452\,
            I => \N__55432\
        );

    \I__12903\ : CascadeMux
    port map (
            O => \N__55451\,
            I => \N__55424\
        );

    \I__12902\ : InMux
    port map (
            O => \N__55450\,
            I => \N__55420\
        );

    \I__12901\ : InMux
    port map (
            O => \N__55449\,
            I => \N__55417\
        );

    \I__12900\ : InMux
    port map (
            O => \N__55448\,
            I => \N__55410\
        );

    \I__12899\ : InMux
    port map (
            O => \N__55447\,
            I => \N__55410\
        );

    \I__12898\ : InMux
    port map (
            O => \N__55446\,
            I => \N__55410\
        );

    \I__12897\ : InMux
    port map (
            O => \N__55445\,
            I => \N__55406\
        );

    \I__12896\ : InMux
    port map (
            O => \N__55444\,
            I => \N__55403\
        );

    \I__12895\ : LocalMux
    port map (
            O => \N__55439\,
            I => \N__55400\
        );

    \I__12894\ : InMux
    port map (
            O => \N__55438\,
            I => \N__55396\
        );

    \I__12893\ : LocalMux
    port map (
            O => \N__55435\,
            I => \N__55391\
        );

    \I__12892\ : LocalMux
    port map (
            O => \N__55432\,
            I => \N__55391\
        );

    \I__12891\ : InMux
    port map (
            O => \N__55431\,
            I => \N__55388\
        );

    \I__12890\ : InMux
    port map (
            O => \N__55430\,
            I => \N__55383\
        );

    \I__12889\ : InMux
    port map (
            O => \N__55429\,
            I => \N__55376\
        );

    \I__12888\ : InMux
    port map (
            O => \N__55428\,
            I => \N__55376\
        );

    \I__12887\ : InMux
    port map (
            O => \N__55427\,
            I => \N__55376\
        );

    \I__12886\ : InMux
    port map (
            O => \N__55424\,
            I => \N__55373\
        );

    \I__12885\ : InMux
    port map (
            O => \N__55423\,
            I => \N__55370\
        );

    \I__12884\ : LocalMux
    port map (
            O => \N__55420\,
            I => \N__55367\
        );

    \I__12883\ : LocalMux
    port map (
            O => \N__55417\,
            I => \N__55362\
        );

    \I__12882\ : LocalMux
    port map (
            O => \N__55410\,
            I => \N__55362\
        );

    \I__12881\ : InMux
    port map (
            O => \N__55409\,
            I => \N__55359\
        );

    \I__12880\ : LocalMux
    port map (
            O => \N__55406\,
            I => \N__55352\
        );

    \I__12879\ : LocalMux
    port map (
            O => \N__55403\,
            I => \N__55352\
        );

    \I__12878\ : Span4Mux_h
    port map (
            O => \N__55400\,
            I => \N__55352\
        );

    \I__12877\ : InMux
    port map (
            O => \N__55399\,
            I => \N__55348\
        );

    \I__12876\ : LocalMux
    port map (
            O => \N__55396\,
            I => \N__55345\
        );

    \I__12875\ : Span4Mux_v
    port map (
            O => \N__55391\,
            I => \N__55342\
        );

    \I__12874\ : LocalMux
    port map (
            O => \N__55388\,
            I => \N__55339\
        );

    \I__12873\ : InMux
    port map (
            O => \N__55387\,
            I => \N__55336\
        );

    \I__12872\ : InMux
    port map (
            O => \N__55386\,
            I => \N__55333\
        );

    \I__12871\ : LocalMux
    port map (
            O => \N__55383\,
            I => \N__55328\
        );

    \I__12870\ : LocalMux
    port map (
            O => \N__55376\,
            I => \N__55328\
        );

    \I__12869\ : LocalMux
    port map (
            O => \N__55373\,
            I => \N__55319\
        );

    \I__12868\ : LocalMux
    port map (
            O => \N__55370\,
            I => \N__55319\
        );

    \I__12867\ : Span4Mux_h
    port map (
            O => \N__55367\,
            I => \N__55319\
        );

    \I__12866\ : Span4Mux_h
    port map (
            O => \N__55362\,
            I => \N__55319\
        );

    \I__12865\ : LocalMux
    port map (
            O => \N__55359\,
            I => \N__55314\
        );

    \I__12864\ : Span4Mux_v
    port map (
            O => \N__55352\,
            I => \N__55314\
        );

    \I__12863\ : InMux
    port map (
            O => \N__55351\,
            I => \N__55311\
        );

    \I__12862\ : LocalMux
    port map (
            O => \N__55348\,
            I => \N__55306\
        );

    \I__12861\ : Span4Mux_h
    port map (
            O => \N__55345\,
            I => \N__55306\
        );

    \I__12860\ : Span4Mux_h
    port map (
            O => \N__55342\,
            I => \N__55303\
        );

    \I__12859\ : Span4Mux_v
    port map (
            O => \N__55339\,
            I => \N__55296\
        );

    \I__12858\ : LocalMux
    port map (
            O => \N__55336\,
            I => \N__55296\
        );

    \I__12857\ : LocalMux
    port map (
            O => \N__55333\,
            I => \N__55296\
        );

    \I__12856\ : Span4Mux_h
    port map (
            O => \N__55328\,
            I => \N__55291\
        );

    \I__12855\ : Span4Mux_v
    port map (
            O => \N__55319\,
            I => \N__55291\
        );

    \I__12854\ : Span4Mux_h
    port map (
            O => \N__55314\,
            I => \N__55288\
        );

    \I__12853\ : LocalMux
    port map (
            O => \N__55311\,
            I => \N__55283\
        );

    \I__12852\ : Span4Mux_v
    port map (
            O => \N__55306\,
            I => \N__55283\
        );

    \I__12851\ : Span4Mux_h
    port map (
            O => \N__55303\,
            I => \N__55278\
        );

    \I__12850\ : Span4Mux_v
    port map (
            O => \N__55296\,
            I => \N__55278\
        );

    \I__12849\ : Span4Mux_h
    port map (
            O => \N__55291\,
            I => \N__55275\
        );

    \I__12848\ : Span4Mux_v
    port map (
            O => \N__55288\,
            I => \N__55272\
        );

    \I__12847\ : Odrv4
    port map (
            O => \N__55283\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270\
        );

    \I__12846\ : Odrv4
    port map (
            O => \N__55278\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270\
        );

    \I__12845\ : Odrv4
    port map (
            O => \N__55275\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270\
        );

    \I__12844\ : Odrv4
    port map (
            O => \N__55272\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270\
        );

    \I__12843\ : InMux
    port map (
            O => \N__55263\,
            I => \N__55259\
        );

    \I__12842\ : InMux
    port map (
            O => \N__55262\,
            I => \N__55251\
        );

    \I__12841\ : LocalMux
    port map (
            O => \N__55259\,
            I => \N__55246\
        );

    \I__12840\ : InMux
    port map (
            O => \N__55258\,
            I => \N__55239\
        );

    \I__12839\ : InMux
    port map (
            O => \N__55257\,
            I => \N__55239\
        );

    \I__12838\ : InMux
    port map (
            O => \N__55256\,
            I => \N__55239\
        );

    \I__12837\ : InMux
    port map (
            O => \N__55255\,
            I => \N__55236\
        );

    \I__12836\ : InMux
    port map (
            O => \N__55254\,
            I => \N__55233\
        );

    \I__12835\ : LocalMux
    port map (
            O => \N__55251\,
            I => \N__55225\
        );

    \I__12834\ : InMux
    port map (
            O => \N__55250\,
            I => \N__55222\
        );

    \I__12833\ : InMux
    port map (
            O => \N__55249\,
            I => \N__55218\
        );

    \I__12832\ : Span4Mux_h
    port map (
            O => \N__55246\,
            I => \N__55212\
        );

    \I__12831\ : LocalMux
    port map (
            O => \N__55239\,
            I => \N__55212\
        );

    \I__12830\ : LocalMux
    port map (
            O => \N__55236\,
            I => \N__55209\
        );

    \I__12829\ : LocalMux
    port map (
            O => \N__55233\,
            I => \N__55206\
        );

    \I__12828\ : InMux
    port map (
            O => \N__55232\,
            I => \N__55199\
        );

    \I__12827\ : InMux
    port map (
            O => \N__55231\,
            I => \N__55199\
        );

    \I__12826\ : InMux
    port map (
            O => \N__55230\,
            I => \N__55199\
        );

    \I__12825\ : InMux
    port map (
            O => \N__55229\,
            I => \N__55193\
        );

    \I__12824\ : InMux
    port map (
            O => \N__55228\,
            I => \N__55193\
        );

    \I__12823\ : Span4Mux_v
    port map (
            O => \N__55225\,
            I => \N__55187\
        );

    \I__12822\ : LocalMux
    port map (
            O => \N__55222\,
            I => \N__55187\
        );

    \I__12821\ : InMux
    port map (
            O => \N__55221\,
            I => \N__55184\
        );

    \I__12820\ : LocalMux
    port map (
            O => \N__55218\,
            I => \N__55180\
        );

    \I__12819\ : InMux
    port map (
            O => \N__55217\,
            I => \N__55177\
        );

    \I__12818\ : Span4Mux_h
    port map (
            O => \N__55212\,
            I => \N__55174\
        );

    \I__12817\ : Span4Mux_h
    port map (
            O => \N__55209\,
            I => \N__55167\
        );

    \I__12816\ : Span4Mux_v
    port map (
            O => \N__55206\,
            I => \N__55167\
        );

    \I__12815\ : LocalMux
    port map (
            O => \N__55199\,
            I => \N__55167\
        );

    \I__12814\ : InMux
    port map (
            O => \N__55198\,
            I => \N__55164\
        );

    \I__12813\ : LocalMux
    port map (
            O => \N__55193\,
            I => \N__55160\
        );

    \I__12812\ : CascadeMux
    port map (
            O => \N__55192\,
            I => \N__55157\
        );

    \I__12811\ : Span4Mux_h
    port map (
            O => \N__55187\,
            I => \N__55151\
        );

    \I__12810\ : LocalMux
    port map (
            O => \N__55184\,
            I => \N__55148\
        );

    \I__12809\ : InMux
    port map (
            O => \N__55183\,
            I => \N__55145\
        );

    \I__12808\ : Span4Mux_h
    port map (
            O => \N__55180\,
            I => \N__55140\
        );

    \I__12807\ : LocalMux
    port map (
            O => \N__55177\,
            I => \N__55140\
        );

    \I__12806\ : Span4Mux_v
    port map (
            O => \N__55174\,
            I => \N__55135\
        );

    \I__12805\ : Span4Mux_h
    port map (
            O => \N__55167\,
            I => \N__55135\
        );

    \I__12804\ : LocalMux
    port map (
            O => \N__55164\,
            I => \N__55132\
        );

    \I__12803\ : InMux
    port map (
            O => \N__55163\,
            I => \N__55129\
        );

    \I__12802\ : Span4Mux_v
    port map (
            O => \N__55160\,
            I => \N__55126\
        );

    \I__12801\ : InMux
    port map (
            O => \N__55157\,
            I => \N__55123\
        );

    \I__12800\ : InMux
    port map (
            O => \N__55156\,
            I => \N__55120\
        );

    \I__12799\ : InMux
    port map (
            O => \N__55155\,
            I => \N__55117\
        );

    \I__12798\ : InMux
    port map (
            O => \N__55154\,
            I => \N__55114\
        );

    \I__12797\ : Span4Mux_h
    port map (
            O => \N__55151\,
            I => \N__55110\
        );

    \I__12796\ : Span4Mux_h
    port map (
            O => \N__55148\,
            I => \N__55105\
        );

    \I__12795\ : LocalMux
    port map (
            O => \N__55145\,
            I => \N__55105\
        );

    \I__12794\ : Span4Mux_h
    port map (
            O => \N__55140\,
            I => \N__55098\
        );

    \I__12793\ : Span4Mux_h
    port map (
            O => \N__55135\,
            I => \N__55098\
        );

    \I__12792\ : Span4Mux_v
    port map (
            O => \N__55132\,
            I => \N__55098\
        );

    \I__12791\ : LocalMux
    port map (
            O => \N__55129\,
            I => \N__55085\
        );

    \I__12790\ : Sp12to4
    port map (
            O => \N__55126\,
            I => \N__55085\
        );

    \I__12789\ : LocalMux
    port map (
            O => \N__55123\,
            I => \N__55085\
        );

    \I__12788\ : LocalMux
    port map (
            O => \N__55120\,
            I => \N__55085\
        );

    \I__12787\ : LocalMux
    port map (
            O => \N__55117\,
            I => \N__55085\
        );

    \I__12786\ : LocalMux
    port map (
            O => \N__55114\,
            I => \N__55085\
        );

    \I__12785\ : InMux
    port map (
            O => \N__55113\,
            I => \N__55082\
        );

    \I__12784\ : Span4Mux_v
    port map (
            O => \N__55110\,
            I => \N__55079\
        );

    \I__12783\ : Span4Mux_v
    port map (
            O => \N__55105\,
            I => \N__55076\
        );

    \I__12782\ : Sp12to4
    port map (
            O => \N__55098\,
            I => \N__55069\
        );

    \I__12781\ : Span12Mux_h
    port map (
            O => \N__55085\,
            I => \N__55069\
        );

    \I__12780\ : LocalMux
    port map (
            O => \N__55082\,
            I => \N__55069\
        );

    \I__12779\ : Odrv4
    port map (
            O => \N__55079\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274\
        );

    \I__12778\ : Odrv4
    port map (
            O => \N__55076\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274\
        );

    \I__12777\ : Odrv12
    port map (
            O => \N__55069\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274\
        );

    \I__12776\ : CascadeMux
    port map (
            O => \N__55062\,
            I => \N__55059\
        );

    \I__12775\ : InMux
    port map (
            O => \N__55059\,
            I => \N__55049\
        );

    \I__12774\ : InMux
    port map (
            O => \N__55058\,
            I => \N__55046\
        );

    \I__12773\ : InMux
    port map (
            O => \N__55057\,
            I => \N__55043\
        );

    \I__12772\ : InMux
    port map (
            O => \N__55056\,
            I => \N__55040\
        );

    \I__12771\ : InMux
    port map (
            O => \N__55055\,
            I => \N__55037\
        );

    \I__12770\ : InMux
    port map (
            O => \N__55054\,
            I => \N__55032\
        );

    \I__12769\ : CascadeMux
    port map (
            O => \N__55053\,
            I => \N__55026\
        );

    \I__12768\ : CascadeMux
    port map (
            O => \N__55052\,
            I => \N__55023\
        );

    \I__12767\ : LocalMux
    port map (
            O => \N__55049\,
            I => \N__55014\
        );

    \I__12766\ : LocalMux
    port map (
            O => \N__55046\,
            I => \N__55014\
        );

    \I__12765\ : LocalMux
    port map (
            O => \N__55043\,
            I => \N__55011\
        );

    \I__12764\ : LocalMux
    port map (
            O => \N__55040\,
            I => \N__55005\
        );

    \I__12763\ : LocalMux
    port map (
            O => \N__55037\,
            I => \N__55005\
        );

    \I__12762\ : InMux
    port map (
            O => \N__55036\,
            I => \N__55002\
        );

    \I__12761\ : CascadeMux
    port map (
            O => \N__55035\,
            I => \N__54998\
        );

    \I__12760\ : LocalMux
    port map (
            O => \N__55032\,
            I => \N__54995\
        );

    \I__12759\ : InMux
    port map (
            O => \N__55031\,
            I => \N__54992\
        );

    \I__12758\ : InMux
    port map (
            O => \N__55030\,
            I => \N__54989\
        );

    \I__12757\ : InMux
    port map (
            O => \N__55029\,
            I => \N__54986\
        );

    \I__12756\ : InMux
    port map (
            O => \N__55026\,
            I => \N__54979\
        );

    \I__12755\ : InMux
    port map (
            O => \N__55023\,
            I => \N__54979\
        );

    \I__12754\ : InMux
    port map (
            O => \N__55022\,
            I => \N__54979\
        );

    \I__12753\ : InMux
    port map (
            O => \N__55021\,
            I => \N__54976\
        );

    \I__12752\ : InMux
    port map (
            O => \N__55020\,
            I => \N__54973\
        );

    \I__12751\ : CascadeMux
    port map (
            O => \N__55019\,
            I => \N__54970\
        );

    \I__12750\ : Span4Mux_v
    port map (
            O => \N__55014\,
            I => \N__54967\
        );

    \I__12749\ : Span4Mux_v
    port map (
            O => \N__55011\,
            I => \N__54964\
        );

    \I__12748\ : InMux
    port map (
            O => \N__55010\,
            I => \N__54960\
        );

    \I__12747\ : Span4Mux_v
    port map (
            O => \N__55005\,
            I => \N__54955\
        );

    \I__12746\ : LocalMux
    port map (
            O => \N__55002\,
            I => \N__54955\
        );

    \I__12745\ : InMux
    port map (
            O => \N__55001\,
            I => \N__54950\
        );

    \I__12744\ : InMux
    port map (
            O => \N__54998\,
            I => \N__54947\
        );

    \I__12743\ : Span4Mux_v
    port map (
            O => \N__54995\,
            I => \N__54944\
        );

    \I__12742\ : LocalMux
    port map (
            O => \N__54992\,
            I => \N__54939\
        );

    \I__12741\ : LocalMux
    port map (
            O => \N__54989\,
            I => \N__54939\
        );

    \I__12740\ : LocalMux
    port map (
            O => \N__54986\,
            I => \N__54930\
        );

    \I__12739\ : LocalMux
    port map (
            O => \N__54979\,
            I => \N__54930\
        );

    \I__12738\ : LocalMux
    port map (
            O => \N__54976\,
            I => \N__54930\
        );

    \I__12737\ : LocalMux
    port map (
            O => \N__54973\,
            I => \N__54930\
        );

    \I__12736\ : InMux
    port map (
            O => \N__54970\,
            I => \N__54925\
        );

    \I__12735\ : Span4Mux_v
    port map (
            O => \N__54967\,
            I => \N__54920\
        );

    \I__12734\ : Span4Mux_v
    port map (
            O => \N__54964\,
            I => \N__54920\
        );

    \I__12733\ : InMux
    port map (
            O => \N__54963\,
            I => \N__54917\
        );

    \I__12732\ : LocalMux
    port map (
            O => \N__54960\,
            I => \N__54914\
        );

    \I__12731\ : Span4Mux_v
    port map (
            O => \N__54955\,
            I => \N__54911\
        );

    \I__12730\ : InMux
    port map (
            O => \N__54954\,
            I => \N__54908\
        );

    \I__12729\ : InMux
    port map (
            O => \N__54953\,
            I => \N__54905\
        );

    \I__12728\ : LocalMux
    port map (
            O => \N__54950\,
            I => \N__54902\
        );

    \I__12727\ : LocalMux
    port map (
            O => \N__54947\,
            I => \N__54893\
        );

    \I__12726\ : Span4Mux_h
    port map (
            O => \N__54944\,
            I => \N__54893\
        );

    \I__12725\ : Span4Mux_v
    port map (
            O => \N__54939\,
            I => \N__54893\
        );

    \I__12724\ : Span4Mux_v
    port map (
            O => \N__54930\,
            I => \N__54893\
        );

    \I__12723\ : InMux
    port map (
            O => \N__54929\,
            I => \N__54888\
        );

    \I__12722\ : InMux
    port map (
            O => \N__54928\,
            I => \N__54888\
        );

    \I__12721\ : LocalMux
    port map (
            O => \N__54925\,
            I => \N__54885\
        );

    \I__12720\ : Span4Mux_h
    port map (
            O => \N__54920\,
            I => \N__54882\
        );

    \I__12719\ : LocalMux
    port map (
            O => \N__54917\,
            I => \N__54879\
        );

    \I__12718\ : Span4Mux_v
    port map (
            O => \N__54914\,
            I => \N__54874\
        );

    \I__12717\ : Span4Mux_h
    port map (
            O => \N__54911\,
            I => \N__54874\
        );

    \I__12716\ : LocalMux
    port map (
            O => \N__54908\,
            I => \N__54871\
        );

    \I__12715\ : LocalMux
    port map (
            O => \N__54905\,
            I => \N__54862\
        );

    \I__12714\ : Span4Mux_v
    port map (
            O => \N__54902\,
            I => \N__54862\
        );

    \I__12713\ : Span4Mux_h
    port map (
            O => \N__54893\,
            I => \N__54862\
        );

    \I__12712\ : LocalMux
    port map (
            O => \N__54888\,
            I => \N__54862\
        );

    \I__12711\ : Span12Mux_h
    port map (
            O => \N__54885\,
            I => \N__54859\
        );

    \I__12710\ : Sp12to4
    port map (
            O => \N__54882\,
            I => \N__54854\
        );

    \I__12709\ : Span12Mux_v
    port map (
            O => \N__54879\,
            I => \N__54854\
        );

    \I__12708\ : Span4Mux_h
    port map (
            O => \N__54874\,
            I => \N__54851\
        );

    \I__12707\ : Span4Mux_v
    port map (
            O => \N__54871\,
            I => \N__54846\
        );

    \I__12706\ : Span4Mux_h
    port map (
            O => \N__54862\,
            I => \N__54846\
        );

    \I__12705\ : Odrv12
    port map (
            O => \N__54859\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0\
        );

    \I__12704\ : Odrv12
    port map (
            O => \N__54854\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0\
        );

    \I__12703\ : Odrv4
    port map (
            O => \N__54851\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0\
        );

    \I__12702\ : Odrv4
    port map (
            O => \N__54846\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0\
        );

    \I__12701\ : InMux
    port map (
            O => \N__54837\,
            I => \N__54829\
        );

    \I__12700\ : CascadeMux
    port map (
            O => \N__54836\,
            I => \N__54826\
        );

    \I__12699\ : CascadeMux
    port map (
            O => \N__54835\,
            I => \N__54822\
        );

    \I__12698\ : InMux
    port map (
            O => \N__54834\,
            I => \N__54813\
        );

    \I__12697\ : InMux
    port map (
            O => \N__54833\,
            I => \N__54810\
        );

    \I__12696\ : InMux
    port map (
            O => \N__54832\,
            I => \N__54807\
        );

    \I__12695\ : LocalMux
    port map (
            O => \N__54829\,
            I => \N__54803\
        );

    \I__12694\ : InMux
    port map (
            O => \N__54826\,
            I => \N__54799\
        );

    \I__12693\ : InMux
    port map (
            O => \N__54825\,
            I => \N__54795\
        );

    \I__12692\ : InMux
    port map (
            O => \N__54822\,
            I => \N__54792\
        );

    \I__12691\ : InMux
    port map (
            O => \N__54821\,
            I => \N__54789\
        );

    \I__12690\ : InMux
    port map (
            O => \N__54820\,
            I => \N__54784\
        );

    \I__12689\ : InMux
    port map (
            O => \N__54819\,
            I => \N__54784\
        );

    \I__12688\ : InMux
    port map (
            O => \N__54818\,
            I => \N__54775\
        );

    \I__12687\ : InMux
    port map (
            O => \N__54817\,
            I => \N__54775\
        );

    \I__12686\ : InMux
    port map (
            O => \N__54816\,
            I => \N__54772\
        );

    \I__12685\ : LocalMux
    port map (
            O => \N__54813\,
            I => \N__54769\
        );

    \I__12684\ : LocalMux
    port map (
            O => \N__54810\,
            I => \N__54764\
        );

    \I__12683\ : LocalMux
    port map (
            O => \N__54807\,
            I => \N__54764\
        );

    \I__12682\ : InMux
    port map (
            O => \N__54806\,
            I => \N__54761\
        );

    \I__12681\ : Span4Mux_h
    port map (
            O => \N__54803\,
            I => \N__54758\
        );

    \I__12680\ : InMux
    port map (
            O => \N__54802\,
            I => \N__54753\
        );

    \I__12679\ : LocalMux
    port map (
            O => \N__54799\,
            I => \N__54750\
        );

    \I__12678\ : InMux
    port map (
            O => \N__54798\,
            I => \N__54747\
        );

    \I__12677\ : LocalMux
    port map (
            O => \N__54795\,
            I => \N__54744\
        );

    \I__12676\ : LocalMux
    port map (
            O => \N__54792\,
            I => \N__54737\
        );

    \I__12675\ : LocalMux
    port map (
            O => \N__54789\,
            I => \N__54737\
        );

    \I__12674\ : LocalMux
    port map (
            O => \N__54784\,
            I => \N__54737\
        );

    \I__12673\ : InMux
    port map (
            O => \N__54783\,
            I => \N__54732\
        );

    \I__12672\ : InMux
    port map (
            O => \N__54782\,
            I => \N__54729\
        );

    \I__12671\ : InMux
    port map (
            O => \N__54781\,
            I => \N__54724\
        );

    \I__12670\ : InMux
    port map (
            O => \N__54780\,
            I => \N__54724\
        );

    \I__12669\ : LocalMux
    port map (
            O => \N__54775\,
            I => \N__54721\
        );

    \I__12668\ : LocalMux
    port map (
            O => \N__54772\,
            I => \N__54712\
        );

    \I__12667\ : Span4Mux_v
    port map (
            O => \N__54769\,
            I => \N__54712\
        );

    \I__12666\ : Span4Mux_h
    port map (
            O => \N__54764\,
            I => \N__54712\
        );

    \I__12665\ : LocalMux
    port map (
            O => \N__54761\,
            I => \N__54712\
        );

    \I__12664\ : Span4Mux_v
    port map (
            O => \N__54758\,
            I => \N__54709\
        );

    \I__12663\ : InMux
    port map (
            O => \N__54757\,
            I => \N__54706\
        );

    \I__12662\ : InMux
    port map (
            O => \N__54756\,
            I => \N__54703\
        );

    \I__12661\ : LocalMux
    port map (
            O => \N__54753\,
            I => \N__54698\
        );

    \I__12660\ : Span4Mux_v
    port map (
            O => \N__54750\,
            I => \N__54698\
        );

    \I__12659\ : LocalMux
    port map (
            O => \N__54747\,
            I => \N__54691\
        );

    \I__12658\ : Span4Mux_h
    port map (
            O => \N__54744\,
            I => \N__54691\
        );

    \I__12657\ : Span4Mux_v
    port map (
            O => \N__54737\,
            I => \N__54691\
        );

    \I__12656\ : InMux
    port map (
            O => \N__54736\,
            I => \N__54686\
        );

    \I__12655\ : InMux
    port map (
            O => \N__54735\,
            I => \N__54686\
        );

    \I__12654\ : LocalMux
    port map (
            O => \N__54732\,
            I => \N__54675\
        );

    \I__12653\ : LocalMux
    port map (
            O => \N__54729\,
            I => \N__54675\
        );

    \I__12652\ : LocalMux
    port map (
            O => \N__54724\,
            I => \N__54675\
        );

    \I__12651\ : Span4Mux_v
    port map (
            O => \N__54721\,
            I => \N__54675\
        );

    \I__12650\ : Span4Mux_v
    port map (
            O => \N__54712\,
            I => \N__54675\
        );

    \I__12649\ : Span4Mux_h
    port map (
            O => \N__54709\,
            I => \N__54672\
        );

    \I__12648\ : LocalMux
    port map (
            O => \N__54706\,
            I => \N__54669\
        );

    \I__12647\ : LocalMux
    port map (
            O => \N__54703\,
            I => \N__54660\
        );

    \I__12646\ : Span4Mux_h
    port map (
            O => \N__54698\,
            I => \N__54660\
        );

    \I__12645\ : Span4Mux_h
    port map (
            O => \N__54691\,
            I => \N__54660\
        );

    \I__12644\ : LocalMux
    port map (
            O => \N__54686\,
            I => \N__54660\
        );

    \I__12643\ : Span4Mux_h
    port map (
            O => \N__54675\,
            I => \N__54657\
        );

    \I__12642\ : Span4Mux_h
    port map (
            O => \N__54672\,
            I => \N__54654\
        );

    \I__12641\ : Span4Mux_v
    port map (
            O => \N__54669\,
            I => \N__54649\
        );

    \I__12640\ : Span4Mux_h
    port map (
            O => \N__54660\,
            I => \N__54649\
        );

    \I__12639\ : Span4Mux_h
    port map (
            O => \N__54657\,
            I => \N__54646\
        );

    \I__12638\ : Odrv4
    port map (
            O => \N__54654\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270\
        );

    \I__12637\ : Odrv4
    port map (
            O => \N__54649\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270\
        );

    \I__12636\ : Odrv4
    port map (
            O => \N__54646\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270\
        );

    \I__12635\ : InMux
    port map (
            O => \N__54639\,
            I => \N__54635\
        );

    \I__12634\ : CascadeMux
    port map (
            O => \N__54638\,
            I => \N__54631\
        );

    \I__12633\ : LocalMux
    port map (
            O => \N__54635\,
            I => \N__54628\
        );

    \I__12632\ : InMux
    port map (
            O => \N__54634\,
            I => \N__54623\
        );

    \I__12631\ : InMux
    port map (
            O => \N__54631\,
            I => \N__54623\
        );

    \I__12630\ : Span4Mux_h
    port map (
            O => \N__54628\,
            I => \N__54620\
        );

    \I__12629\ : LocalMux
    port map (
            O => \N__54623\,
            I => \N__54617\
        );

    \I__12628\ : Span4Mux_v
    port map (
            O => \N__54620\,
            I => \N__54614\
        );

    \I__12627\ : Span4Mux_v
    port map (
            O => \N__54617\,
            I => \N__54611\
        );

    \I__12626\ : Span4Mux_h
    port map (
            O => \N__54614\,
            I => \N__54606\
        );

    \I__12625\ : Span4Mux_h
    port map (
            O => \N__54611\,
            I => \N__54606\
        );

    \I__12624\ : Odrv4
    port map (
            O => \N__54606\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_1
        );

    \I__12623\ : InMux
    port map (
            O => \N__54603\,
            I => \N__54600\
        );

    \I__12622\ : LocalMux
    port map (
            O => \N__54600\,
            I => \N__54595\
        );

    \I__12621\ : InMux
    port map (
            O => \N__54599\,
            I => \N__54592\
        );

    \I__12620\ : InMux
    port map (
            O => \N__54598\,
            I => \N__54589\
        );

    \I__12619\ : Span12Mux_h
    port map (
            O => \N__54595\,
            I => \N__54586\
        );

    \I__12618\ : LocalMux
    port map (
            O => \N__54592\,
            I => \N__54581\
        );

    \I__12617\ : LocalMux
    port map (
            O => \N__54589\,
            I => \N__54581\
        );

    \I__12616\ : Odrv12
    port map (
            O => \N__54586\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_1
        );

    \I__12615\ : Odrv12
    port map (
            O => \N__54581\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_1
        );

    \I__12614\ : InMux
    port map (
            O => \N__54576\,
            I => \N__54573\
        );

    \I__12613\ : LocalMux
    port map (
            O => \N__54573\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_1\
        );

    \I__12612\ : InMux
    port map (
            O => \N__54570\,
            I => \N__54567\
        );

    \I__12611\ : LocalMux
    port map (
            O => \N__54567\,
            I => \N__54564\
        );

    \I__12610\ : Span12Mux_h
    port map (
            O => \N__54564\,
            I => \N__54561\
        );

    \I__12609\ : Odrv12
    port map (
            O => \N__54561\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_3_26\
        );

    \I__12608\ : InMux
    port map (
            O => \N__54558\,
            I => \N__54555\
        );

    \I__12607\ : LocalMux
    port map (
            O => \N__54555\,
            I => \N__54552\
        );

    \I__12606\ : Span12Mux_v
    port map (
            O => \N__54552\,
            I => \N__54549\
        );

    \I__12605\ : Odrv12
    port map (
            O => \N__54549\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_4093_0\
        );

    \I__12604\ : CascadeMux
    port map (
            O => \N__54546\,
            I => \N__54543\
        );

    \I__12603\ : InMux
    port map (
            O => \N__54543\,
            I => \N__54540\
        );

    \I__12602\ : LocalMux
    port map (
            O => \N__54540\,
            I => \N__54537\
        );

    \I__12601\ : Span4Mux_h
    port map (
            O => \N__54537\,
            I => \N__54534\
        );

    \I__12600\ : Span4Mux_h
    port map (
            O => \N__54534\,
            I => \N__54531\
        );

    \I__12599\ : Span4Mux_h
    port map (
            O => \N__54531\,
            I => \N__54528\
        );

    \I__12598\ : Odrv4
    port map (
            O => \N__54528\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_26\
        );

    \I__12597\ : CEMux
    port map (
            O => \N__54525\,
            I => \N__54429\
        );

    \I__12596\ : CEMux
    port map (
            O => \N__54524\,
            I => \N__54429\
        );

    \I__12595\ : CEMux
    port map (
            O => \N__54523\,
            I => \N__54429\
        );

    \I__12594\ : CEMux
    port map (
            O => \N__54522\,
            I => \N__54429\
        );

    \I__12593\ : CEMux
    port map (
            O => \N__54521\,
            I => \N__54429\
        );

    \I__12592\ : CEMux
    port map (
            O => \N__54520\,
            I => \N__54429\
        );

    \I__12591\ : CEMux
    port map (
            O => \N__54519\,
            I => \N__54429\
        );

    \I__12590\ : CEMux
    port map (
            O => \N__54518\,
            I => \N__54429\
        );

    \I__12589\ : CEMux
    port map (
            O => \N__54517\,
            I => \N__54429\
        );

    \I__12588\ : CEMux
    port map (
            O => \N__54516\,
            I => \N__54429\
        );

    \I__12587\ : CEMux
    port map (
            O => \N__54515\,
            I => \N__54429\
        );

    \I__12586\ : CEMux
    port map (
            O => \N__54514\,
            I => \N__54429\
        );

    \I__12585\ : CEMux
    port map (
            O => \N__54513\,
            I => \N__54429\
        );

    \I__12584\ : CEMux
    port map (
            O => \N__54512\,
            I => \N__54429\
        );

    \I__12583\ : CEMux
    port map (
            O => \N__54511\,
            I => \N__54429\
        );

    \I__12582\ : CEMux
    port map (
            O => \N__54510\,
            I => \N__54429\
        );

    \I__12581\ : CEMux
    port map (
            O => \N__54509\,
            I => \N__54429\
        );

    \I__12580\ : CEMux
    port map (
            O => \N__54508\,
            I => \N__54429\
        );

    \I__12579\ : CEMux
    port map (
            O => \N__54507\,
            I => \N__54429\
        );

    \I__12578\ : CEMux
    port map (
            O => \N__54506\,
            I => \N__54429\
        );

    \I__12577\ : CEMux
    port map (
            O => \N__54505\,
            I => \N__54429\
        );

    \I__12576\ : CEMux
    port map (
            O => \N__54504\,
            I => \N__54429\
        );

    \I__12575\ : CEMux
    port map (
            O => \N__54503\,
            I => \N__54429\
        );

    \I__12574\ : CEMux
    port map (
            O => \N__54502\,
            I => \N__54429\
        );

    \I__12573\ : CEMux
    port map (
            O => \N__54501\,
            I => \N__54429\
        );

    \I__12572\ : CEMux
    port map (
            O => \N__54500\,
            I => \N__54429\
        );

    \I__12571\ : CEMux
    port map (
            O => \N__54499\,
            I => \N__54429\
        );

    \I__12570\ : CEMux
    port map (
            O => \N__54498\,
            I => \N__54429\
        );

    \I__12569\ : CEMux
    port map (
            O => \N__54497\,
            I => \N__54429\
        );

    \I__12568\ : CEMux
    port map (
            O => \N__54496\,
            I => \N__54429\
        );

    \I__12567\ : CEMux
    port map (
            O => \N__54495\,
            I => \N__54429\
        );

    \I__12566\ : CEMux
    port map (
            O => \N__54494\,
            I => \N__54429\
        );

    \I__12565\ : GlobalMux
    port map (
            O => \N__54429\,
            I => \N__54426\
        );

    \I__12564\ : gio2CtrlBuf
    port map (
            O => \N__54426\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_g\
        );

    \I__12563\ : InMux
    port map (
            O => \N__54423\,
            I => \N__54420\
        );

    \I__12562\ : LocalMux
    port map (
            O => \N__54420\,
            I => \N__54416\
        );

    \I__12561\ : InMux
    port map (
            O => \N__54419\,
            I => \N__54413\
        );

    \I__12560\ : Span4Mux_v
    port map (
            O => \N__54416\,
            I => \N__54410\
        );

    \I__12559\ : LocalMux
    port map (
            O => \N__54413\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i\
        );

    \I__12558\ : Odrv4
    port map (
            O => \N__54410\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i\
        );

    \I__12557\ : CascadeMux
    port map (
            O => \N__54405\,
            I => \N__54399\
        );

    \I__12556\ : InMux
    port map (
            O => \N__54404\,
            I => \N__54395\
        );

    \I__12555\ : InMux
    port map (
            O => \N__54403\,
            I => \N__54392\
        );

    \I__12554\ : InMux
    port map (
            O => \N__54402\,
            I => \N__54389\
        );

    \I__12553\ : InMux
    port map (
            O => \N__54399\,
            I => \N__54384\
        );

    \I__12552\ : InMux
    port map (
            O => \N__54398\,
            I => \N__54384\
        );

    \I__12551\ : LocalMux
    port map (
            O => \N__54395\,
            I => \N__54381\
        );

    \I__12550\ : LocalMux
    port map (
            O => \N__54392\,
            I => \N__54373\
        );

    \I__12549\ : LocalMux
    port map (
            O => \N__54389\,
            I => \N__54373\
        );

    \I__12548\ : LocalMux
    port map (
            O => \N__54384\,
            I => \N__54373\
        );

    \I__12547\ : Span4Mux_v
    port map (
            O => \N__54381\,
            I => \N__54370\
        );

    \I__12546\ : InMux
    port map (
            O => \N__54380\,
            I => \N__54367\
        );

    \I__12545\ : Span4Mux_h
    port map (
            O => \N__54373\,
            I => \N__54364\
        );

    \I__12544\ : Sp12to4
    port map (
            O => \N__54370\,
            I => \N__54359\
        );

    \I__12543\ : LocalMux
    port map (
            O => \N__54367\,
            I => \N__54359\
        );

    \I__12542\ : Span4Mux_h
    port map (
            O => \N__54364\,
            I => \N__54356\
        );

    \I__12541\ : Odrv12
    port map (
            O => \N__54359\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0\
        );

    \I__12540\ : Odrv4
    port map (
            O => \N__54356\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0\
        );

    \I__12539\ : CascadeMux
    port map (
            O => \N__54351\,
            I => \N__54348\
        );

    \I__12538\ : InMux
    port map (
            O => \N__54348\,
            I => \N__54345\
        );

    \I__12537\ : LocalMux
    port map (
            O => \N__54345\,
            I => \N__54339\
        );

    \I__12536\ : InMux
    port map (
            O => \N__54344\,
            I => \N__54331\
        );

    \I__12535\ : InMux
    port map (
            O => \N__54343\,
            I => \N__54326\
        );

    \I__12534\ : InMux
    port map (
            O => \N__54342\,
            I => \N__54326\
        );

    \I__12533\ : Span4Mux_v
    port map (
            O => \N__54339\,
            I => \N__54323\
        );

    \I__12532\ : InMux
    port map (
            O => \N__54338\,
            I => \N__54320\
        );

    \I__12531\ : InMux
    port map (
            O => \N__54337\,
            I => \N__54315\
        );

    \I__12530\ : InMux
    port map (
            O => \N__54336\,
            I => \N__54315\
        );

    \I__12529\ : InMux
    port map (
            O => \N__54335\,
            I => \N__54312\
        );

    \I__12528\ : InMux
    port map (
            O => \N__54334\,
            I => \N__54309\
        );

    \I__12527\ : LocalMux
    port map (
            O => \N__54331\,
            I => \N__54306\
        );

    \I__12526\ : LocalMux
    port map (
            O => \N__54326\,
            I => \N__54303\
        );

    \I__12525\ : Span4Mux_h
    port map (
            O => \N__54323\,
            I => \N__54300\
        );

    \I__12524\ : LocalMux
    port map (
            O => \N__54320\,
            I => \N__54293\
        );

    \I__12523\ : LocalMux
    port map (
            O => \N__54315\,
            I => \N__54293\
        );

    \I__12522\ : LocalMux
    port map (
            O => \N__54312\,
            I => \N__54293\
        );

    \I__12521\ : LocalMux
    port map (
            O => \N__54309\,
            I => \N__54290\
        );

    \I__12520\ : Span12Mux_v
    port map (
            O => \N__54306\,
            I => \N__54285\
        );

    \I__12519\ : Span4Mux_v
    port map (
            O => \N__54303\,
            I => \N__54282\
        );

    \I__12518\ : Span4Mux_h
    port map (
            O => \N__54300\,
            I => \N__54277\
        );

    \I__12517\ : Span4Mux_v
    port map (
            O => \N__54293\,
            I => \N__54277\
        );

    \I__12516\ : Span4Mux_h
    port map (
            O => \N__54290\,
            I => \N__54274\
        );

    \I__12515\ : InMux
    port map (
            O => \N__54289\,
            I => \N__54269\
        );

    \I__12514\ : InMux
    port map (
            O => \N__54288\,
            I => \N__54269\
        );

    \I__12513\ : Odrv12
    port map (
            O => \N__54285\,
            I => \s_paddr_I2C_3\
        );

    \I__12512\ : Odrv4
    port map (
            O => \N__54282\,
            I => \s_paddr_I2C_3\
        );

    \I__12511\ : Odrv4
    port map (
            O => \N__54277\,
            I => \s_paddr_I2C_3\
        );

    \I__12510\ : Odrv4
    port map (
            O => \N__54274\,
            I => \s_paddr_I2C_3\
        );

    \I__12509\ : LocalMux
    port map (
            O => \N__54269\,
            I => \s_paddr_I2C_3\
        );

    \I__12508\ : InMux
    port map (
            O => \N__54258\,
            I => \N__54255\
        );

    \I__12507\ : LocalMux
    port map (
            O => \N__54255\,
            I => \N__54252\
        );

    \I__12506\ : Span4Mux_v
    port map (
            O => \N__54252\,
            I => \N__54248\
        );

    \I__12505\ : InMux
    port map (
            O => \N__54251\,
            I => \N__54245\
        );

    \I__12504\ : Odrv4
    port map (
            O => \N__54248\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0\
        );

    \I__12503\ : LocalMux
    port map (
            O => \N__54245\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0\
        );

    \I__12502\ : CascadeMux
    port map (
            O => \N__54240\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_230_cascade_\
        );

    \I__12501\ : InMux
    port map (
            O => \N__54237\,
            I => \N__54234\
        );

    \I__12500\ : LocalMux
    port map (
            O => \N__54234\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_0_sqmuxa\
        );

    \I__12499\ : CascadeMux
    port map (
            O => \N__54231\,
            I => \N__54228\
        );

    \I__12498\ : InMux
    port map (
            O => \N__54228\,
            I => \N__54225\
        );

    \I__12497\ : LocalMux
    port map (
            O => \N__54225\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_2_sqmuxa\
        );

    \I__12496\ : InMux
    port map (
            O => \N__54222\,
            I => \N__54219\
        );

    \I__12495\ : LocalMux
    port map (
            O => \N__54219\,
            I => \N__54216\
        );

    \I__12494\ : Span4Mux_v
    port map (
            O => \N__54216\,
            I => \N__54213\
        );

    \I__12493\ : Span4Mux_h
    port map (
            O => \N__54213\,
            I => \N__54210\
        );

    \I__12492\ : Odrv4
    port map (
            O => \N__54210\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_24\
        );

    \I__12491\ : InMux
    port map (
            O => \N__54207\,
            I => \N__54203\
        );

    \I__12490\ : InMux
    port map (
            O => \N__54206\,
            I => \N__54200\
        );

    \I__12489\ : LocalMux
    port map (
            O => \N__54203\,
            I => \N__54197\
        );

    \I__12488\ : LocalMux
    port map (
            O => \N__54200\,
            I => \N__54194\
        );

    \I__12487\ : Span4Mux_h
    port map (
            O => \N__54197\,
            I => \N__54190\
        );

    \I__12486\ : Span4Mux_h
    port map (
            O => \N__54194\,
            I => \N__54187\
        );

    \I__12485\ : InMux
    port map (
            O => \N__54193\,
            I => \N__54184\
        );

    \I__12484\ : Odrv4
    port map (
            O => \N__54190\,
            I => cemf_module_64ch_ctrl_inst1_data_config_16
        );

    \I__12483\ : Odrv4
    port map (
            O => \N__54187\,
            I => cemf_module_64ch_ctrl_inst1_data_config_16
        );

    \I__12482\ : LocalMux
    port map (
            O => \N__54184\,
            I => cemf_module_64ch_ctrl_inst1_data_config_16
        );

    \I__12481\ : InMux
    port map (
            O => \N__54177\,
            I => \N__54174\
        );

    \I__12480\ : LocalMux
    port map (
            O => \N__54174\,
            I => \N__54171\
        );

    \I__12479\ : Span12Mux_v
    port map (
            O => \N__54171\,
            I => \N__54168\
        );

    \I__12478\ : Odrv12
    port map (
            O => \N__54168\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_28\
        );

    \I__12477\ : CascadeMux
    port map (
            O => \N__54165\,
            I => \N__54162\
        );

    \I__12476\ : InMux
    port map (
            O => \N__54162\,
            I => \N__54159\
        );

    \I__12475\ : LocalMux
    port map (
            O => \N__54159\,
            I => \N__54156\
        );

    \I__12474\ : Span4Mux_v
    port map (
            O => \N__54156\,
            I => \N__54153\
        );

    \I__12473\ : Span4Mux_h
    port map (
            O => \N__54153\,
            I => \N__54149\
        );

    \I__12472\ : InMux
    port map (
            O => \N__54152\,
            I => \N__54146\
        );

    \I__12471\ : Span4Mux_h
    port map (
            O => \N__54149\,
            I => \N__54143\
        );

    \I__12470\ : LocalMux
    port map (
            O => \N__54146\,
            I => \N__54139\
        );

    \I__12469\ : Span4Mux_h
    port map (
            O => \N__54143\,
            I => \N__54136\
        );

    \I__12468\ : InMux
    port map (
            O => \N__54142\,
            I => \N__54133\
        );

    \I__12467\ : Span4Mux_h
    port map (
            O => \N__54139\,
            I => \N__54130\
        );

    \I__12466\ : Odrv4
    port map (
            O => \N__54136\,
            I => cemf_module_64ch_ctrl_inst1_data_config_17
        );

    \I__12465\ : LocalMux
    port map (
            O => \N__54133\,
            I => cemf_module_64ch_ctrl_inst1_data_config_17
        );

    \I__12464\ : Odrv4
    port map (
            O => \N__54130\,
            I => cemf_module_64ch_ctrl_inst1_data_config_17
        );

    \I__12463\ : CEMux
    port map (
            O => \N__54123\,
            I => \N__54120\
        );

    \I__12462\ : LocalMux
    port map (
            O => \N__54120\,
            I => \N__54115\
        );

    \I__12461\ : CEMux
    port map (
            O => \N__54119\,
            I => \N__54109\
        );

    \I__12460\ : CEMux
    port map (
            O => \N__54118\,
            I => \N__54106\
        );

    \I__12459\ : Span4Mux_h
    port map (
            O => \N__54115\,
            I => \N__54103\
        );

    \I__12458\ : CEMux
    port map (
            O => \N__54114\,
            I => \N__54100\
        );

    \I__12457\ : CEMux
    port map (
            O => \N__54113\,
            I => \N__54097\
        );

    \I__12456\ : CEMux
    port map (
            O => \N__54112\,
            I => \N__54094\
        );

    \I__12455\ : LocalMux
    port map (
            O => \N__54109\,
            I => \N__54091\
        );

    \I__12454\ : LocalMux
    port map (
            O => \N__54106\,
            I => \N__54086\
        );

    \I__12453\ : Span4Mux_v
    port map (
            O => \N__54103\,
            I => \N__54086\
        );

    \I__12452\ : LocalMux
    port map (
            O => \N__54100\,
            I => \N__54083\
        );

    \I__12451\ : LocalMux
    port map (
            O => \N__54097\,
            I => \N__54080\
        );

    \I__12450\ : LocalMux
    port map (
            O => \N__54094\,
            I => \N__54077\
        );

    \I__12449\ : Span4Mux_h
    port map (
            O => \N__54091\,
            I => \N__54074\
        );

    \I__12448\ : Span4Mux_h
    port map (
            O => \N__54086\,
            I => \N__54071\
        );

    \I__12447\ : Span12Mux_h
    port map (
            O => \N__54083\,
            I => \N__54068\
        );

    \I__12446\ : Span4Mux_h
    port map (
            O => \N__54080\,
            I => \N__54065\
        );

    \I__12445\ : Span4Mux_h
    port map (
            O => \N__54077\,
            I => \N__54060\
        );

    \I__12444\ : Span4Mux_h
    port map (
            O => \N__54074\,
            I => \N__54060\
        );

    \I__12443\ : Span4Mux_h
    port map (
            O => \N__54071\,
            I => \N__54057\
        );

    \I__12442\ : Odrv12
    port map (
            O => \N__54068\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0\
        );

    \I__12441\ : Odrv4
    port map (
            O => \N__54065\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0\
        );

    \I__12440\ : Odrv4
    port map (
            O => \N__54060\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0\
        );

    \I__12439\ : Odrv4
    port map (
            O => \N__54057\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0\
        );

    \I__12438\ : CascadeMux
    port map (
            O => \N__54048\,
            I => \N__54045\
        );

    \I__12437\ : InMux
    port map (
            O => \N__54045\,
            I => \N__54042\
        );

    \I__12436\ : LocalMux
    port map (
            O => \N__54042\,
            I => \N__54039\
        );

    \I__12435\ : Span4Mux_h
    port map (
            O => \N__54039\,
            I => \N__54036\
        );

    \I__12434\ : Span4Mux_h
    port map (
            O => \N__54036\,
            I => \N__54033\
        );

    \I__12433\ : Odrv4
    port map (
            O => \N__54033\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_1\
        );

    \I__12432\ : CascadeMux
    port map (
            O => \N__54030\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RLZ0Z7_cascade_\
        );

    \I__12431\ : InMux
    port map (
            O => \N__54027\,
            I => \N__54024\
        );

    \I__12430\ : LocalMux
    port map (
            O => \N__54024\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1\
        );

    \I__12429\ : InMux
    port map (
            O => \N__54021\,
            I => \N__54018\
        );

    \I__12428\ : LocalMux
    port map (
            O => \N__54018\,
            I => \N__54015\
        );

    \I__12427\ : Span4Mux_v
    port map (
            O => \N__54015\,
            I => \N__54012\
        );

    \I__12426\ : Odrv4
    port map (
            O => \N__54012\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_0\
        );

    \I__12425\ : CascadeMux
    port map (
            O => \N__54009\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_cascade_\
        );

    \I__12424\ : InMux
    port map (
            O => \N__54006\,
            I => \N__53998\
        );

    \I__12423\ : InMux
    port map (
            O => \N__54005\,
            I => \N__53995\
        );

    \I__12422\ : InMux
    port map (
            O => \N__54004\,
            I => \N__53988\
        );

    \I__12421\ : InMux
    port map (
            O => \N__54003\,
            I => \N__53985\
        );

    \I__12420\ : InMux
    port map (
            O => \N__54002\,
            I => \N__53980\
        );

    \I__12419\ : InMux
    port map (
            O => \N__54001\,
            I => \N__53980\
        );

    \I__12418\ : LocalMux
    port map (
            O => \N__53998\,
            I => \N__53973\
        );

    \I__12417\ : LocalMux
    port map (
            O => \N__53995\,
            I => \N__53970\
        );

    \I__12416\ : CascadeMux
    port map (
            O => \N__53994\,
            I => \N__53963\
        );

    \I__12415\ : InMux
    port map (
            O => \N__53993\,
            I => \N__53956\
        );

    \I__12414\ : InMux
    port map (
            O => \N__53992\,
            I => \N__53953\
        );

    \I__12413\ : InMux
    port map (
            O => \N__53991\,
            I => \N__53950\
        );

    \I__12412\ : LocalMux
    port map (
            O => \N__53988\,
            I => \N__53945\
        );

    \I__12411\ : LocalMux
    port map (
            O => \N__53985\,
            I => \N__53942\
        );

    \I__12410\ : LocalMux
    port map (
            O => \N__53980\,
            I => \N__53939\
        );

    \I__12409\ : InMux
    port map (
            O => \N__53979\,
            I => \N__53934\
        );

    \I__12408\ : InMux
    port map (
            O => \N__53978\,
            I => \N__53934\
        );

    \I__12407\ : InMux
    port map (
            O => \N__53977\,
            I => \N__53931\
        );

    \I__12406\ : InMux
    port map (
            O => \N__53976\,
            I => \N__53928\
        );

    \I__12405\ : Span4Mux_v
    port map (
            O => \N__53973\,
            I => \N__53925\
        );

    \I__12404\ : Span4Mux_h
    port map (
            O => \N__53970\,
            I => \N__53922\
        );

    \I__12403\ : InMux
    port map (
            O => \N__53969\,
            I => \N__53919\
        );

    \I__12402\ : InMux
    port map (
            O => \N__53968\,
            I => \N__53914\
        );

    \I__12401\ : InMux
    port map (
            O => \N__53967\,
            I => \N__53914\
        );

    \I__12400\ : InMux
    port map (
            O => \N__53966\,
            I => \N__53911\
        );

    \I__12399\ : InMux
    port map (
            O => \N__53963\,
            I => \N__53908\
        );

    \I__12398\ : InMux
    port map (
            O => \N__53962\,
            I => \N__53905\
        );

    \I__12397\ : InMux
    port map (
            O => \N__53961\,
            I => \N__53902\
        );

    \I__12396\ : InMux
    port map (
            O => \N__53960\,
            I => \N__53899\
        );

    \I__12395\ : InMux
    port map (
            O => \N__53959\,
            I => \N__53896\
        );

    \I__12394\ : LocalMux
    port map (
            O => \N__53956\,
            I => \N__53893\
        );

    \I__12393\ : LocalMux
    port map (
            O => \N__53953\,
            I => \N__53888\
        );

    \I__12392\ : LocalMux
    port map (
            O => \N__53950\,
            I => \N__53888\
        );

    \I__12391\ : InMux
    port map (
            O => \N__53949\,
            I => \N__53885\
        );

    \I__12390\ : InMux
    port map (
            O => \N__53948\,
            I => \N__53882\
        );

    \I__12389\ : Span4Mux_v
    port map (
            O => \N__53945\,
            I => \N__53879\
        );

    \I__12388\ : Span4Mux_v
    port map (
            O => \N__53942\,
            I => \N__53874\
        );

    \I__12387\ : Span4Mux_v
    port map (
            O => \N__53939\,
            I => \N__53874\
        );

    \I__12386\ : LocalMux
    port map (
            O => \N__53934\,
            I => \N__53871\
        );

    \I__12385\ : LocalMux
    port map (
            O => \N__53931\,
            I => \N__53868\
        );

    \I__12384\ : LocalMux
    port map (
            O => \N__53928\,
            I => \N__53865\
        );

    \I__12383\ : Span4Mux_h
    port map (
            O => \N__53925\,
            I => \N__53858\
        );

    \I__12382\ : Span4Mux_v
    port map (
            O => \N__53922\,
            I => \N__53858\
        );

    \I__12381\ : LocalMux
    port map (
            O => \N__53919\,
            I => \N__53858\
        );

    \I__12380\ : LocalMux
    port map (
            O => \N__53914\,
            I => \N__53853\
        );

    \I__12379\ : LocalMux
    port map (
            O => \N__53911\,
            I => \N__53853\
        );

    \I__12378\ : LocalMux
    port map (
            O => \N__53908\,
            I => \N__53832\
        );

    \I__12377\ : LocalMux
    port map (
            O => \N__53905\,
            I => \N__53832\
        );

    \I__12376\ : LocalMux
    port map (
            O => \N__53902\,
            I => \N__53832\
        );

    \I__12375\ : LocalMux
    port map (
            O => \N__53899\,
            I => \N__53832\
        );

    \I__12374\ : LocalMux
    port map (
            O => \N__53896\,
            I => \N__53832\
        );

    \I__12373\ : Sp12to4
    port map (
            O => \N__53893\,
            I => \N__53832\
        );

    \I__12372\ : Span12Mux_v
    port map (
            O => \N__53888\,
            I => \N__53832\
        );

    \I__12371\ : LocalMux
    port map (
            O => \N__53885\,
            I => \N__53832\
        );

    \I__12370\ : LocalMux
    port map (
            O => \N__53882\,
            I => \N__53832\
        );

    \I__12369\ : Sp12to4
    port map (
            O => \N__53879\,
            I => \N__53832\
        );

    \I__12368\ : Span4Mux_h
    port map (
            O => \N__53874\,
            I => \N__53827\
        );

    \I__12367\ : Span4Mux_v
    port map (
            O => \N__53871\,
            I => \N__53827\
        );

    \I__12366\ : Span4Mux_h
    port map (
            O => \N__53868\,
            I => \N__53824\
        );

    \I__12365\ : Span4Mux_v
    port map (
            O => \N__53865\,
            I => \N__53819\
        );

    \I__12364\ : Span4Mux_h
    port map (
            O => \N__53858\,
            I => \N__53819\
        );

    \I__12363\ : Sp12to4
    port map (
            O => \N__53853\,
            I => \N__53816\
        );

    \I__12362\ : Span12Mux_h
    port map (
            O => \N__53832\,
            I => \N__53813\
        );

    \I__12361\ : Span4Mux_h
    port map (
            O => \N__53827\,
            I => \N__53810\
        );

    \I__12360\ : Span4Mux_v
    port map (
            O => \N__53824\,
            I => \N__53805\
        );

    \I__12359\ : Span4Mux_v
    port map (
            O => \N__53819\,
            I => \N__53805\
        );

    \I__12358\ : Span12Mux_v
    port map (
            O => \N__53816\,
            I => \N__53802\
        );

    \I__12357\ : Odrv12
    port map (
            O => \N__53813\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273\
        );

    \I__12356\ : Odrv4
    port map (
            O => \N__53810\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273\
        );

    \I__12355\ : Odrv4
    port map (
            O => \N__53805\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273\
        );

    \I__12354\ : Odrv12
    port map (
            O => \N__53802\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273\
        );

    \I__12353\ : CascadeMux
    port map (
            O => \N__53793\,
            I => \N__53789\
        );

    \I__12352\ : InMux
    port map (
            O => \N__53792\,
            I => \N__53785\
        );

    \I__12351\ : InMux
    port map (
            O => \N__53789\,
            I => \N__53782\
        );

    \I__12350\ : InMux
    port map (
            O => \N__53788\,
            I => \N__53779\
        );

    \I__12349\ : LocalMux
    port map (
            O => \N__53785\,
            I => \N__53776\
        );

    \I__12348\ : LocalMux
    port map (
            O => \N__53782\,
            I => \N__53773\
        );

    \I__12347\ : LocalMux
    port map (
            O => \N__53779\,
            I => \N__53770\
        );

    \I__12346\ : Span4Mux_v
    port map (
            O => \N__53776\,
            I => \N__53767\
        );

    \I__12345\ : Span4Mux_h
    port map (
            O => \N__53773\,
            I => \N__53764\
        );

    \I__12344\ : Span4Mux_v
    port map (
            O => \N__53770\,
            I => \N__53761\
        );

    \I__12343\ : Span4Mux_v
    port map (
            O => \N__53767\,
            I => \N__53756\
        );

    \I__12342\ : Span4Mux_h
    port map (
            O => \N__53764\,
            I => \N__53756\
        );

    \I__12341\ : Sp12to4
    port map (
            O => \N__53761\,
            I => \N__53753\
        );

    \I__12340\ : Span4Mux_v
    port map (
            O => \N__53756\,
            I => \N__53750\
        );

    \I__12339\ : Odrv12
    port map (
            O => \N__53753\,
            I => cemf_module_64ch_ctrl_inst1_data_config_2
        );

    \I__12338\ : Odrv4
    port map (
            O => \N__53750\,
            I => cemf_module_64ch_ctrl_inst1_data_config_2
        );

    \I__12337\ : CascadeMux
    port map (
            O => \N__53745\,
            I => \N__53742\
        );

    \I__12336\ : InMux
    port map (
            O => \N__53742\,
            I => \N__53739\
        );

    \I__12335\ : LocalMux
    port map (
            O => \N__53739\,
            I => \N__53736\
        );

    \I__12334\ : Span4Mux_h
    port map (
            O => \N__53736\,
            I => \N__53733\
        );

    \I__12333\ : Odrv4
    port map (
            O => \N__53733\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_2\
        );

    \I__12332\ : InMux
    port map (
            O => \N__53730\,
            I => \N__53727\
        );

    \I__12331\ : LocalMux
    port map (
            O => \N__53727\,
            I => \N__53724\
        );

    \I__12330\ : Odrv12
    port map (
            O => \N__53724\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_2\
        );

    \I__12329\ : InMux
    port map (
            O => \N__53721\,
            I => \N__53709\
        );

    \I__12328\ : InMux
    port map (
            O => \N__53720\,
            I => \N__53704\
        );

    \I__12327\ : InMux
    port map (
            O => \N__53719\,
            I => \N__53704\
        );

    \I__12326\ : InMux
    port map (
            O => \N__53718\,
            I => \N__53701\
        );

    \I__12325\ : InMux
    port map (
            O => \N__53717\,
            I => \N__53696\
        );

    \I__12324\ : InMux
    port map (
            O => \N__53716\,
            I => \N__53696\
        );

    \I__12323\ : InMux
    port map (
            O => \N__53715\,
            I => \N__53684\
        );

    \I__12322\ : InMux
    port map (
            O => \N__53714\,
            I => \N__53684\
        );

    \I__12321\ : InMux
    port map (
            O => \N__53713\,
            I => \N__53679\
        );

    \I__12320\ : InMux
    port map (
            O => \N__53712\,
            I => \N__53679\
        );

    \I__12319\ : LocalMux
    port map (
            O => \N__53709\,
            I => \N__53676\
        );

    \I__12318\ : LocalMux
    port map (
            O => \N__53704\,
            I => \N__53666\
        );

    \I__12317\ : LocalMux
    port map (
            O => \N__53701\,
            I => \N__53661\
        );

    \I__12316\ : LocalMux
    port map (
            O => \N__53696\,
            I => \N__53661\
        );

    \I__12315\ : InMux
    port map (
            O => \N__53695\,
            I => \N__53656\
        );

    \I__12314\ : InMux
    port map (
            O => \N__53694\,
            I => \N__53656\
        );

    \I__12313\ : InMux
    port map (
            O => \N__53693\,
            I => \N__53651\
        );

    \I__12312\ : InMux
    port map (
            O => \N__53692\,
            I => \N__53651\
        );

    \I__12311\ : InMux
    port map (
            O => \N__53691\,
            I => \N__53648\
        );

    \I__12310\ : InMux
    port map (
            O => \N__53690\,
            I => \N__53643\
        );

    \I__12309\ : InMux
    port map (
            O => \N__53689\,
            I => \N__53643\
        );

    \I__12308\ : LocalMux
    port map (
            O => \N__53684\,
            I => \N__53640\
        );

    \I__12307\ : LocalMux
    port map (
            O => \N__53679\,
            I => \N__53637\
        );

    \I__12306\ : Span4Mux_v
    port map (
            O => \N__53676\,
            I => \N__53634\
        );

    \I__12305\ : InMux
    port map (
            O => \N__53675\,
            I => \N__53629\
        );

    \I__12304\ : InMux
    port map (
            O => \N__53674\,
            I => \N__53629\
        );

    \I__12303\ : InMux
    port map (
            O => \N__53673\,
            I => \N__53626\
        );

    \I__12302\ : InMux
    port map (
            O => \N__53672\,
            I => \N__53623\
        );

    \I__12301\ : InMux
    port map (
            O => \N__53671\,
            I => \N__53620\
        );

    \I__12300\ : InMux
    port map (
            O => \N__53670\,
            I => \N__53615\
        );

    \I__12299\ : InMux
    port map (
            O => \N__53669\,
            I => \N__53615\
        );

    \I__12298\ : Span4Mux_h
    port map (
            O => \N__53666\,
            I => \N__53610\
        );

    \I__12297\ : Span4Mux_v
    port map (
            O => \N__53661\,
            I => \N__53610\
        );

    \I__12296\ : LocalMux
    port map (
            O => \N__53656\,
            I => \N__53607\
        );

    \I__12295\ : LocalMux
    port map (
            O => \N__53651\,
            I => \N__53596\
        );

    \I__12294\ : LocalMux
    port map (
            O => \N__53648\,
            I => \N__53596\
        );

    \I__12293\ : LocalMux
    port map (
            O => \N__53643\,
            I => \N__53596\
        );

    \I__12292\ : Span4Mux_v
    port map (
            O => \N__53640\,
            I => \N__53596\
        );

    \I__12291\ : Span4Mux_v
    port map (
            O => \N__53637\,
            I => \N__53596\
        );

    \I__12290\ : Span4Mux_h
    port map (
            O => \N__53634\,
            I => \N__53593\
        );

    \I__12289\ : LocalMux
    port map (
            O => \N__53629\,
            I => \N__53588\
        );

    \I__12288\ : LocalMux
    port map (
            O => \N__53626\,
            I => \N__53588\
        );

    \I__12287\ : LocalMux
    port map (
            O => \N__53623\,
            I => \N__53585\
        );

    \I__12286\ : LocalMux
    port map (
            O => \N__53620\,
            I => \N__53578\
        );

    \I__12285\ : LocalMux
    port map (
            O => \N__53615\,
            I => \N__53578\
        );

    \I__12284\ : Span4Mux_h
    port map (
            O => \N__53610\,
            I => \N__53578\
        );

    \I__12283\ : Span4Mux_v
    port map (
            O => \N__53607\,
            I => \N__53573\
        );

    \I__12282\ : Span4Mux_h
    port map (
            O => \N__53596\,
            I => \N__53573\
        );

    \I__12281\ : Span4Mux_v
    port map (
            O => \N__53593\,
            I => \N__53568\
        );

    \I__12280\ : Span4Mux_v
    port map (
            O => \N__53588\,
            I => \N__53568\
        );

    \I__12279\ : Sp12to4
    port map (
            O => \N__53585\,
            I => \N__53565\
        );

    \I__12278\ : Span4Mux_h
    port map (
            O => \N__53578\,
            I => \N__53562\
        );

    \I__12277\ : Span4Mux_v
    port map (
            O => \N__53573\,
            I => \N__53559\
        );

    \I__12276\ : Span4Mux_h
    port map (
            O => \N__53568\,
            I => \N__53556\
        );

    \I__12275\ : Odrv12
    port map (
            O => \N__53565\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i\
        );

    \I__12274\ : Odrv4
    port map (
            O => \N__53562\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i\
        );

    \I__12273\ : Odrv4
    port map (
            O => \N__53559\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i\
        );

    \I__12272\ : Odrv4
    port map (
            O => \N__53556\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i\
        );

    \I__12271\ : CascadeMux
    port map (
            O => \N__53547\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGHZ0Z5_cascade_\
        );

    \I__12270\ : InMux
    port map (
            O => \N__53544\,
            I => \N__53541\
        );

    \I__12269\ : LocalMux
    port map (
            O => \N__53541\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17\
        );

    \I__12268\ : CascadeMux
    port map (
            O => \N__53538\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17_cascade_\
        );

    \I__12267\ : InMux
    port map (
            O => \N__53535\,
            I => \N__53532\
        );

    \I__12266\ : LocalMux
    port map (
            O => \N__53532\,
            I => \N__53529\
        );

    \I__12265\ : Odrv12
    port map (
            O => \N__53529\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_17\
        );

    \I__12264\ : InMux
    port map (
            O => \N__53526\,
            I => \N__53521\
        );

    \I__12263\ : CascadeMux
    port map (
            O => \N__53525\,
            I => \N__53518\
        );

    \I__12262\ : InMux
    port map (
            O => \N__53524\,
            I => \N__53515\
        );

    \I__12261\ : LocalMux
    port map (
            O => \N__53521\,
            I => \N__53512\
        );

    \I__12260\ : InMux
    port map (
            O => \N__53518\,
            I => \N__53509\
        );

    \I__12259\ : LocalMux
    port map (
            O => \N__53515\,
            I => \N__53504\
        );

    \I__12258\ : Span4Mux_h
    port map (
            O => \N__53512\,
            I => \N__53504\
        );

    \I__12257\ : LocalMux
    port map (
            O => \N__53509\,
            I => \N__53501\
        );

    \I__12256\ : Odrv4
    port map (
            O => \N__53504\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_16
        );

    \I__12255\ : Odrv4
    port map (
            O => \N__53501\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_16
        );

    \I__12254\ : CascadeMux
    port map (
            O => \N__53496\,
            I => \N__53493\
        );

    \I__12253\ : InMux
    port map (
            O => \N__53493\,
            I => \N__53490\
        );

    \I__12252\ : LocalMux
    port map (
            O => \N__53490\,
            I => \N__53487\
        );

    \I__12251\ : Span4Mux_h
    port map (
            O => \N__53487\,
            I => \N__53484\
        );

    \I__12250\ : Odrv4
    port map (
            O => \N__53484\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_16\
        );

    \I__12249\ : InMux
    port map (
            O => \N__53481\,
            I => \N__53478\
        );

    \I__12248\ : LocalMux
    port map (
            O => \N__53478\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_16\
        );

    \I__12247\ : CascadeMux
    port map (
            O => \N__53475\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGHZ0Z5_cascade_\
        );

    \I__12246\ : InMux
    port map (
            O => \N__53472\,
            I => \N__53469\
        );

    \I__12245\ : LocalMux
    port map (
            O => \N__53469\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16\
        );

    \I__12244\ : InMux
    port map (
            O => \N__53466\,
            I => \N__53463\
        );

    \I__12243\ : LocalMux
    port map (
            O => \N__53463\,
            I => \N__53460\
        );

    \I__12242\ : Odrv12
    port map (
            O => \N__53460\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_15\
        );

    \I__12241\ : CascadeMux
    port map (
            O => \N__53457\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16_cascade_\
        );

    \I__12240\ : InMux
    port map (
            O => \N__53454\,
            I => \N__53451\
        );

    \I__12239\ : LocalMux
    port map (
            O => \N__53451\,
            I => \N__53448\
        );

    \I__12238\ : Odrv4
    port map (
            O => \N__53448\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_16\
        );

    \I__12237\ : InMux
    port map (
            O => \N__53445\,
            I => \N__53442\
        );

    \I__12236\ : LocalMux
    port map (
            O => \N__53442\,
            I => \N__53439\
        );

    \I__12235\ : Span12Mux_v
    port map (
            O => \N__53439\,
            I => \N__53436\
        );

    \I__12234\ : Span12Mux_h
    port map (
            O => \N__53436\,
            I => \N__53433\
        );

    \I__12233\ : Odrv12
    port map (
            O => \N__53433\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_31\
        );

    \I__12232\ : CascadeMux
    port map (
            O => \N__53430\,
            I => \N__53427\
        );

    \I__12231\ : InMux
    port map (
            O => \N__53427\,
            I => \N__53424\
        );

    \I__12230\ : LocalMux
    port map (
            O => \N__53424\,
            I => \N__53421\
        );

    \I__12229\ : Span4Mux_h
    port map (
            O => \N__53421\,
            I => \N__53416\
        );

    \I__12228\ : InMux
    port map (
            O => \N__53420\,
            I => \N__53413\
        );

    \I__12227\ : InMux
    port map (
            O => \N__53419\,
            I => \N__53410\
        );

    \I__12226\ : Span4Mux_h
    port map (
            O => \N__53416\,
            I => \N__53407\
        );

    \I__12225\ : LocalMux
    port map (
            O => \N__53413\,
            I => \N__53404\
        );

    \I__12224\ : LocalMux
    port map (
            O => \N__53410\,
            I => \N__53401\
        );

    \I__12223\ : Span4Mux_h
    port map (
            O => \N__53407\,
            I => \N__53398\
        );

    \I__12222\ : Span4Mux_v
    port map (
            O => \N__53404\,
            I => \N__53393\
        );

    \I__12221\ : Span4Mux_h
    port map (
            O => \N__53401\,
            I => \N__53393\
        );

    \I__12220\ : Span4Mux_h
    port map (
            O => \N__53398\,
            I => \N__53390\
        );

    \I__12219\ : Span4Mux_h
    port map (
            O => \N__53393\,
            I => \N__53387\
        );

    \I__12218\ : Odrv4
    port map (
            O => \N__53390\,
            I => cemf_module_64ch_ctrl_inst1_data_config_14
        );

    \I__12217\ : Odrv4
    port map (
            O => \N__53387\,
            I => cemf_module_64ch_ctrl_inst1_data_config_14
        );

    \I__12216\ : CascadeMux
    port map (
            O => \N__53382\,
            I => \N__53379\
        );

    \I__12215\ : InMux
    port map (
            O => \N__53379\,
            I => \N__53376\
        );

    \I__12214\ : LocalMux
    port map (
            O => \N__53376\,
            I => \N__53372\
        );

    \I__12213\ : InMux
    port map (
            O => \N__53375\,
            I => \N__53368\
        );

    \I__12212\ : Span4Mux_v
    port map (
            O => \N__53372\,
            I => \N__53365\
        );

    \I__12211\ : InMux
    port map (
            O => \N__53371\,
            I => \N__53362\
        );

    \I__12210\ : LocalMux
    port map (
            O => \N__53368\,
            I => \N__53359\
        );

    \I__12209\ : Span4Mux_h
    port map (
            O => \N__53365\,
            I => \N__53356\
        );

    \I__12208\ : LocalMux
    port map (
            O => \N__53362\,
            I => \N__53351\
        );

    \I__12207\ : Span4Mux_h
    port map (
            O => \N__53359\,
            I => \N__53351\
        );

    \I__12206\ : Span4Mux_h
    port map (
            O => \N__53356\,
            I => \N__53348\
        );

    \I__12205\ : Span4Mux_h
    port map (
            O => \N__53351\,
            I => \N__53345\
        );

    \I__12204\ : Odrv4
    port map (
            O => \N__53348\,
            I => cemf_module_64ch_ctrl_inst1_data_config_15
        );

    \I__12203\ : Odrv4
    port map (
            O => \N__53345\,
            I => cemf_module_64ch_ctrl_inst1_data_config_15
        );

    \I__12202\ : InMux
    port map (
            O => \N__53340\,
            I => \N__53337\
        );

    \I__12201\ : LocalMux
    port map (
            O => \N__53337\,
            I => \N__53334\
        );

    \I__12200\ : Odrv4
    port map (
            O => \N__53334\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_25\
        );

    \I__12199\ : InMux
    port map (
            O => \N__53331\,
            I => \N__53325\
        );

    \I__12198\ : CascadeMux
    port map (
            O => \N__53330\,
            I => \N__53320\
        );

    \I__12197\ : CascadeMux
    port map (
            O => \N__53329\,
            I => \N__53311\
        );

    \I__12196\ : CascadeMux
    port map (
            O => \N__53328\,
            I => \N__53307\
        );

    \I__12195\ : LocalMux
    port map (
            O => \N__53325\,
            I => \N__53303\
        );

    \I__12194\ : CascadeMux
    port map (
            O => \N__53324\,
            I => \N__53300\
        );

    \I__12193\ : CascadeMux
    port map (
            O => \N__53323\,
            I => \N__53297\
        );

    \I__12192\ : InMux
    port map (
            O => \N__53320\,
            I => \N__53293\
        );

    \I__12191\ : CascadeMux
    port map (
            O => \N__53319\,
            I => \N__53290\
        );

    \I__12190\ : CascadeMux
    port map (
            O => \N__53318\,
            I => \N__53287\
        );

    \I__12189\ : CascadeMux
    port map (
            O => \N__53317\,
            I => \N__53283\
        );

    \I__12188\ : CascadeMux
    port map (
            O => \N__53316\,
            I => \N__53278\
        );

    \I__12187\ : CascadeMux
    port map (
            O => \N__53315\,
            I => \N__53275\
        );

    \I__12186\ : InMux
    port map (
            O => \N__53314\,
            I => \N__53272\
        );

    \I__12185\ : InMux
    port map (
            O => \N__53311\,
            I => \N__53267\
        );

    \I__12184\ : CascadeMux
    port map (
            O => \N__53310\,
            I => \N__53263\
        );

    \I__12183\ : InMux
    port map (
            O => \N__53307\,
            I => \N__53259\
        );

    \I__12182\ : CascadeMux
    port map (
            O => \N__53306\,
            I => \N__53253\
        );

    \I__12181\ : Span4Mux_v
    port map (
            O => \N__53303\,
            I => \N__53250\
        );

    \I__12180\ : InMux
    port map (
            O => \N__53300\,
            I => \N__53247\
        );

    \I__12179\ : InMux
    port map (
            O => \N__53297\,
            I => \N__53244\
        );

    \I__12178\ : InMux
    port map (
            O => \N__53296\,
            I => \N__53241\
        );

    \I__12177\ : LocalMux
    port map (
            O => \N__53293\,
            I => \N__53238\
        );

    \I__12176\ : InMux
    port map (
            O => \N__53290\,
            I => \N__53235\
        );

    \I__12175\ : InMux
    port map (
            O => \N__53287\,
            I => \N__53232\
        );

    \I__12174\ : InMux
    port map (
            O => \N__53286\,
            I => \N__53229\
        );

    \I__12173\ : InMux
    port map (
            O => \N__53283\,
            I => \N__53226\
        );

    \I__12172\ : InMux
    port map (
            O => \N__53282\,
            I => \N__53223\
        );

    \I__12171\ : InMux
    port map (
            O => \N__53281\,
            I => \N__53220\
        );

    \I__12170\ : InMux
    port map (
            O => \N__53278\,
            I => \N__53217\
        );

    \I__12169\ : InMux
    port map (
            O => \N__53275\,
            I => \N__53214\
        );

    \I__12168\ : LocalMux
    port map (
            O => \N__53272\,
            I => \N__53211\
        );

    \I__12167\ : InMux
    port map (
            O => \N__53271\,
            I => \N__53208\
        );

    \I__12166\ : InMux
    port map (
            O => \N__53270\,
            I => \N__53205\
        );

    \I__12165\ : LocalMux
    port map (
            O => \N__53267\,
            I => \N__53202\
        );

    \I__12164\ : InMux
    port map (
            O => \N__53266\,
            I => \N__53199\
        );

    \I__12163\ : InMux
    port map (
            O => \N__53263\,
            I => \N__53196\
        );

    \I__12162\ : CascadeMux
    port map (
            O => \N__53262\,
            I => \N__53191\
        );

    \I__12161\ : LocalMux
    port map (
            O => \N__53259\,
            I => \N__53188\
        );

    \I__12160\ : InMux
    port map (
            O => \N__53258\,
            I => \N__53185\
        );

    \I__12159\ : InMux
    port map (
            O => \N__53257\,
            I => \N__53182\
        );

    \I__12158\ : CascadeMux
    port map (
            O => \N__53256\,
            I => \N__53176\
        );

    \I__12157\ : InMux
    port map (
            O => \N__53253\,
            I => \N__53172\
        );

    \I__12156\ : Span4Mux_h
    port map (
            O => \N__53250\,
            I => \N__53167\
        );

    \I__12155\ : LocalMux
    port map (
            O => \N__53247\,
            I => \N__53167\
        );

    \I__12154\ : LocalMux
    port map (
            O => \N__53244\,
            I => \N__53162\
        );

    \I__12153\ : LocalMux
    port map (
            O => \N__53241\,
            I => \N__53162\
        );

    \I__12152\ : Span4Mux_v
    port map (
            O => \N__53238\,
            I => \N__53157\
        );

    \I__12151\ : LocalMux
    port map (
            O => \N__53235\,
            I => \N__53157\
        );

    \I__12150\ : LocalMux
    port map (
            O => \N__53232\,
            I => \N__53154\
        );

    \I__12149\ : LocalMux
    port map (
            O => \N__53229\,
            I => \N__53147\
        );

    \I__12148\ : LocalMux
    port map (
            O => \N__53226\,
            I => \N__53147\
        );

    \I__12147\ : LocalMux
    port map (
            O => \N__53223\,
            I => \N__53147\
        );

    \I__12146\ : LocalMux
    port map (
            O => \N__53220\,
            I => \N__53142\
        );

    \I__12145\ : LocalMux
    port map (
            O => \N__53217\,
            I => \N__53142\
        );

    \I__12144\ : LocalMux
    port map (
            O => \N__53214\,
            I => \N__53137\
        );

    \I__12143\ : Span4Mux_h
    port map (
            O => \N__53211\,
            I => \N__53137\
        );

    \I__12142\ : LocalMux
    port map (
            O => \N__53208\,
            I => \N__53130\
        );

    \I__12141\ : LocalMux
    port map (
            O => \N__53205\,
            I => \N__53130\
        );

    \I__12140\ : Span4Mux_h
    port map (
            O => \N__53202\,
            I => \N__53130\
        );

    \I__12139\ : LocalMux
    port map (
            O => \N__53199\,
            I => \N__53127\
        );

    \I__12138\ : LocalMux
    port map (
            O => \N__53196\,
            I => \N__53124\
        );

    \I__12137\ : InMux
    port map (
            O => \N__53195\,
            I => \N__53119\
        );

    \I__12136\ : InMux
    port map (
            O => \N__53194\,
            I => \N__53119\
        );

    \I__12135\ : InMux
    port map (
            O => \N__53191\,
            I => \N__53116\
        );

    \I__12134\ : Span4Mux_h
    port map (
            O => \N__53188\,
            I => \N__53111\
        );

    \I__12133\ : LocalMux
    port map (
            O => \N__53185\,
            I => \N__53111\
        );

    \I__12132\ : LocalMux
    port map (
            O => \N__53182\,
            I => \N__53108\
        );

    \I__12131\ : InMux
    port map (
            O => \N__53181\,
            I => \N__53097\
        );

    \I__12130\ : InMux
    port map (
            O => \N__53180\,
            I => \N__53097\
        );

    \I__12129\ : InMux
    port map (
            O => \N__53179\,
            I => \N__53097\
        );

    \I__12128\ : InMux
    port map (
            O => \N__53176\,
            I => \N__53097\
        );

    \I__12127\ : InMux
    port map (
            O => \N__53175\,
            I => \N__53097\
        );

    \I__12126\ : LocalMux
    port map (
            O => \N__53172\,
            I => \N__53090\
        );

    \I__12125\ : Span4Mux_h
    port map (
            O => \N__53167\,
            I => \N__53090\
        );

    \I__12124\ : Span4Mux_h
    port map (
            O => \N__53162\,
            I => \N__53090\
        );

    \I__12123\ : Span4Mux_v
    port map (
            O => \N__53157\,
            I => \N__53087\
        );

    \I__12122\ : Span4Mux_v
    port map (
            O => \N__53154\,
            I => \N__53082\
        );

    \I__12121\ : Span4Mux_h
    port map (
            O => \N__53147\,
            I => \N__53082\
        );

    \I__12120\ : Span4Mux_v
    port map (
            O => \N__53142\,
            I => \N__53075\
        );

    \I__12119\ : Span4Mux_h
    port map (
            O => \N__53137\,
            I => \N__53075\
        );

    \I__12118\ : Span4Mux_v
    port map (
            O => \N__53130\,
            I => \N__53075\
        );

    \I__12117\ : Span4Mux_h
    port map (
            O => \N__53127\,
            I => \N__53068\
        );

    \I__12116\ : Span4Mux_v
    port map (
            O => \N__53124\,
            I => \N__53068\
        );

    \I__12115\ : LocalMux
    port map (
            O => \N__53119\,
            I => \N__53068\
        );

    \I__12114\ : LocalMux
    port map (
            O => \N__53116\,
            I => \N__53059\
        );

    \I__12113\ : Span4Mux_v
    port map (
            O => \N__53111\,
            I => \N__53059\
        );

    \I__12112\ : Span4Mux_h
    port map (
            O => \N__53108\,
            I => \N__53059\
        );

    \I__12111\ : LocalMux
    port map (
            O => \N__53097\,
            I => \N__53059\
        );

    \I__12110\ : Span4Mux_v
    port map (
            O => \N__53090\,
            I => \N__53056\
        );

    \I__12109\ : Sp12to4
    port map (
            O => \N__53087\,
            I => \N__53053\
        );

    \I__12108\ : Span4Mux_v
    port map (
            O => \N__53082\,
            I => \N__53048\
        );

    \I__12107\ : Span4Mux_h
    port map (
            O => \N__53075\,
            I => \N__53048\
        );

    \I__12106\ : Span4Mux_h
    port map (
            O => \N__53068\,
            I => \N__53043\
        );

    \I__12105\ : Span4Mux_h
    port map (
            O => \N__53059\,
            I => \N__53043\
        );

    \I__12104\ : Odrv4
    port map (
            O => \N__53056\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0\
        );

    \I__12103\ : Odrv12
    port map (
            O => \N__53053\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0\
        );

    \I__12102\ : Odrv4
    port map (
            O => \N__53048\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0\
        );

    \I__12101\ : Odrv4
    port map (
            O => \N__53043\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0\
        );

    \I__12100\ : CascadeMux
    port map (
            O => \N__53034\,
            I => \N__53031\
        );

    \I__12099\ : InMux
    port map (
            O => \N__53031\,
            I => \N__53028\
        );

    \I__12098\ : LocalMux
    port map (
            O => \N__53028\,
            I => \N__53025\
        );

    \I__12097\ : Span4Mux_v
    port map (
            O => \N__53025\,
            I => \N__53022\
        );

    \I__12096\ : Sp12to4
    port map (
            O => \N__53022\,
            I => \N__53019\
        );

    \I__12095\ : Odrv12
    port map (
            O => \N__53019\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_25\
        );

    \I__12094\ : InMux
    port map (
            O => \N__53016\,
            I => \N__53005\
        );

    \I__12093\ : InMux
    port map (
            O => \N__53015\,
            I => \N__53001\
        );

    \I__12092\ : InMux
    port map (
            O => \N__53014\,
            I => \N__52995\
        );

    \I__12091\ : CascadeMux
    port map (
            O => \N__53013\,
            I => \N__52991\
        );

    \I__12090\ : InMux
    port map (
            O => \N__53012\,
            I => \N__52984\
        );

    \I__12089\ : InMux
    port map (
            O => \N__53011\,
            I => \N__52979\
        );

    \I__12088\ : InMux
    port map (
            O => \N__53010\,
            I => \N__52976\
        );

    \I__12087\ : InMux
    port map (
            O => \N__53009\,
            I => \N__52973\
        );

    \I__12086\ : InMux
    port map (
            O => \N__53008\,
            I => \N__52970\
        );

    \I__12085\ : LocalMux
    port map (
            O => \N__53005\,
            I => \N__52967\
        );

    \I__12084\ : InMux
    port map (
            O => \N__53004\,
            I => \N__52964\
        );

    \I__12083\ : LocalMux
    port map (
            O => \N__53001\,
            I => \N__52961\
        );

    \I__12082\ : InMux
    port map (
            O => \N__53000\,
            I => \N__52958\
        );

    \I__12081\ : InMux
    port map (
            O => \N__52999\,
            I => \N__52955\
        );

    \I__12080\ : InMux
    port map (
            O => \N__52998\,
            I => \N__52952\
        );

    \I__12079\ : LocalMux
    port map (
            O => \N__52995\,
            I => \N__52949\
        );

    \I__12078\ : InMux
    port map (
            O => \N__52994\,
            I => \N__52946\
        );

    \I__12077\ : InMux
    port map (
            O => \N__52991\,
            I => \N__52943\
        );

    \I__12076\ : InMux
    port map (
            O => \N__52990\,
            I => \N__52940\
        );

    \I__12075\ : InMux
    port map (
            O => \N__52989\,
            I => \N__52937\
        );

    \I__12074\ : InMux
    port map (
            O => \N__52988\,
            I => \N__52934\
        );

    \I__12073\ : InMux
    port map (
            O => \N__52987\,
            I => \N__52931\
        );

    \I__12072\ : LocalMux
    port map (
            O => \N__52984\,
            I => \N__52928\
        );

    \I__12071\ : InMux
    port map (
            O => \N__52983\,
            I => \N__52919\
        );

    \I__12070\ : InMux
    port map (
            O => \N__52982\,
            I => \N__52916\
        );

    \I__12069\ : LocalMux
    port map (
            O => \N__52979\,
            I => \N__52911\
        );

    \I__12068\ : LocalMux
    port map (
            O => \N__52976\,
            I => \N__52911\
        );

    \I__12067\ : LocalMux
    port map (
            O => \N__52973\,
            I => \N__52908\
        );

    \I__12066\ : LocalMux
    port map (
            O => \N__52970\,
            I => \N__52905\
        );

    \I__12065\ : Span4Mux_h
    port map (
            O => \N__52967\,
            I => \N__52894\
        );

    \I__12064\ : LocalMux
    port map (
            O => \N__52964\,
            I => \N__52894\
        );

    \I__12063\ : Span4Mux_v
    port map (
            O => \N__52961\,
            I => \N__52894\
        );

    \I__12062\ : LocalMux
    port map (
            O => \N__52958\,
            I => \N__52885\
        );

    \I__12061\ : LocalMux
    port map (
            O => \N__52955\,
            I => \N__52885\
        );

    \I__12060\ : LocalMux
    port map (
            O => \N__52952\,
            I => \N__52885\
        );

    \I__12059\ : Span4Mux_v
    port map (
            O => \N__52949\,
            I => \N__52885\
        );

    \I__12058\ : LocalMux
    port map (
            O => \N__52946\,
            I => \N__52882\
        );

    \I__12057\ : LocalMux
    port map (
            O => \N__52943\,
            I => \N__52877\
        );

    \I__12056\ : LocalMux
    port map (
            O => \N__52940\,
            I => \N__52877\
        );

    \I__12055\ : LocalMux
    port map (
            O => \N__52937\,
            I => \N__52872\
        );

    \I__12054\ : LocalMux
    port map (
            O => \N__52934\,
            I => \N__52872\
        );

    \I__12053\ : LocalMux
    port map (
            O => \N__52931\,
            I => \N__52867\
        );

    \I__12052\ : Span4Mux_v
    port map (
            O => \N__52928\,
            I => \N__52867\
        );

    \I__12051\ : InMux
    port map (
            O => \N__52927\,
            I => \N__52854\
        );

    \I__12050\ : InMux
    port map (
            O => \N__52926\,
            I => \N__52854\
        );

    \I__12049\ : InMux
    port map (
            O => \N__52925\,
            I => \N__52854\
        );

    \I__12048\ : InMux
    port map (
            O => \N__52924\,
            I => \N__52854\
        );

    \I__12047\ : InMux
    port map (
            O => \N__52923\,
            I => \N__52854\
        );

    \I__12046\ : InMux
    port map (
            O => \N__52922\,
            I => \N__52854\
        );

    \I__12045\ : LocalMux
    port map (
            O => \N__52919\,
            I => \N__52847\
        );

    \I__12044\ : LocalMux
    port map (
            O => \N__52916\,
            I => \N__52847\
        );

    \I__12043\ : Span4Mux_h
    port map (
            O => \N__52911\,
            I => \N__52847\
        );

    \I__12042\ : Span4Mux_h
    port map (
            O => \N__52908\,
            I => \N__52842\
        );

    \I__12041\ : Span4Mux_v
    port map (
            O => \N__52905\,
            I => \N__52842\
        );

    \I__12040\ : InMux
    port map (
            O => \N__52904\,
            I => \N__52833\
        );

    \I__12039\ : InMux
    port map (
            O => \N__52903\,
            I => \N__52833\
        );

    \I__12038\ : InMux
    port map (
            O => \N__52902\,
            I => \N__52833\
        );

    \I__12037\ : InMux
    port map (
            O => \N__52901\,
            I => \N__52833\
        );

    \I__12036\ : Span4Mux_h
    port map (
            O => \N__52894\,
            I => \N__52830\
        );

    \I__12035\ : Span4Mux_h
    port map (
            O => \N__52885\,
            I => \N__52827\
        );

    \I__12034\ : Span4Mux_v
    port map (
            O => \N__52882\,
            I => \N__52816\
        );

    \I__12033\ : Span4Mux_v
    port map (
            O => \N__52877\,
            I => \N__52816\
        );

    \I__12032\ : Span4Mux_v
    port map (
            O => \N__52872\,
            I => \N__52816\
        );

    \I__12031\ : Span4Mux_h
    port map (
            O => \N__52867\,
            I => \N__52816\
        );

    \I__12030\ : LocalMux
    port map (
            O => \N__52854\,
            I => \N__52816\
        );

    \I__12029\ : Odrv4
    port map (
            O => \N__52847\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\
        );

    \I__12028\ : Odrv4
    port map (
            O => \N__52842\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\
        );

    \I__12027\ : LocalMux
    port map (
            O => \N__52833\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\
        );

    \I__12026\ : Odrv4
    port map (
            O => \N__52830\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\
        );

    \I__12025\ : Odrv4
    port map (
            O => \N__52827\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\
        );

    \I__12024\ : Odrv4
    port map (
            O => \N__52816\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\
        );

    \I__12023\ : InMux
    port map (
            O => \N__52803\,
            I => \N__52800\
        );

    \I__12022\ : LocalMux
    port map (
            O => \N__52800\,
            I => \N__52797\
        );

    \I__12021\ : Span4Mux_v
    port map (
            O => \N__52797\,
            I => \N__52794\
        );

    \I__12020\ : Span4Mux_h
    port map (
            O => \N__52794\,
            I => \N__52791\
        );

    \I__12019\ : Span4Mux_v
    port map (
            O => \N__52791\,
            I => \N__52788\
        );

    \I__12018\ : Sp12to4
    port map (
            O => \N__52788\,
            I => \N__52785\
        );

    \I__12017\ : Odrv12
    port map (
            O => \N__52785\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_25
        );

    \I__12016\ : InMux
    port map (
            O => \N__52782\,
            I => \N__52776\
        );

    \I__12015\ : InMux
    port map (
            O => \N__52781\,
            I => \N__52773\
        );

    \I__12014\ : InMux
    port map (
            O => \N__52780\,
            I => \N__52765\
        );

    \I__12013\ : InMux
    port map (
            O => \N__52779\,
            I => \N__52762\
        );

    \I__12012\ : LocalMux
    port map (
            O => \N__52776\,
            I => \N__52757\
        );

    \I__12011\ : LocalMux
    port map (
            O => \N__52773\,
            I => \N__52752\
        );

    \I__12010\ : InMux
    port map (
            O => \N__52772\,
            I => \N__52749\
        );

    \I__12009\ : InMux
    port map (
            O => \N__52771\,
            I => \N__52746\
        );

    \I__12008\ : InMux
    port map (
            O => \N__52770\,
            I => \N__52733\
        );

    \I__12007\ : InMux
    port map (
            O => \N__52769\,
            I => \N__52730\
        );

    \I__12006\ : InMux
    port map (
            O => \N__52768\,
            I => \N__52727\
        );

    \I__12005\ : LocalMux
    port map (
            O => \N__52765\,
            I => \N__52722\
        );

    \I__12004\ : LocalMux
    port map (
            O => \N__52762\,
            I => \N__52722\
        );

    \I__12003\ : InMux
    port map (
            O => \N__52761\,
            I => \N__52719\
        );

    \I__12002\ : InMux
    port map (
            O => \N__52760\,
            I => \N__52716\
        );

    \I__12001\ : Span4Mux_v
    port map (
            O => \N__52757\,
            I => \N__52713\
        );

    \I__12000\ : InMux
    port map (
            O => \N__52756\,
            I => \N__52710\
        );

    \I__11999\ : InMux
    port map (
            O => \N__52755\,
            I => \N__52707\
        );

    \I__11998\ : Span4Mux_h
    port map (
            O => \N__52752\,
            I => \N__52702\
        );

    \I__11997\ : LocalMux
    port map (
            O => \N__52749\,
            I => \N__52702\
        );

    \I__11996\ : LocalMux
    port map (
            O => \N__52746\,
            I => \N__52697\
        );

    \I__11995\ : InMux
    port map (
            O => \N__52745\,
            I => \N__52694\
        );

    \I__11994\ : InMux
    port map (
            O => \N__52744\,
            I => \N__52691\
        );

    \I__11993\ : InMux
    port map (
            O => \N__52743\,
            I => \N__52688\
        );

    \I__11992\ : InMux
    port map (
            O => \N__52742\,
            I => \N__52685\
        );

    \I__11991\ : InMux
    port map (
            O => \N__52741\,
            I => \N__52682\
        );

    \I__11990\ : InMux
    port map (
            O => \N__52740\,
            I => \N__52677\
        );

    \I__11989\ : InMux
    port map (
            O => \N__52739\,
            I => \N__52677\
        );

    \I__11988\ : InMux
    port map (
            O => \N__52738\,
            I => \N__52669\
        );

    \I__11987\ : InMux
    port map (
            O => \N__52737\,
            I => \N__52666\
        );

    \I__11986\ : InMux
    port map (
            O => \N__52736\,
            I => \N__52663\
        );

    \I__11985\ : LocalMux
    port map (
            O => \N__52733\,
            I => \N__52660\
        );

    \I__11984\ : LocalMux
    port map (
            O => \N__52730\,
            I => \N__52657\
        );

    \I__11983\ : LocalMux
    port map (
            O => \N__52727\,
            I => \N__52648\
        );

    \I__11982\ : Span4Mux_v
    port map (
            O => \N__52722\,
            I => \N__52648\
        );

    \I__11981\ : LocalMux
    port map (
            O => \N__52719\,
            I => \N__52648\
        );

    \I__11980\ : LocalMux
    port map (
            O => \N__52716\,
            I => \N__52648\
        );

    \I__11979\ : Span4Mux_h
    port map (
            O => \N__52713\,
            I => \N__52643\
        );

    \I__11978\ : LocalMux
    port map (
            O => \N__52710\,
            I => \N__52643\
        );

    \I__11977\ : LocalMux
    port map (
            O => \N__52707\,
            I => \N__52640\
        );

    \I__11976\ : Span4Mux_h
    port map (
            O => \N__52702\,
            I => \N__52637\
        );

    \I__11975\ : InMux
    port map (
            O => \N__52701\,
            I => \N__52634\
        );

    \I__11974\ : InMux
    port map (
            O => \N__52700\,
            I => \N__52631\
        );

    \I__11973\ : Span4Mux_v
    port map (
            O => \N__52697\,
            I => \N__52626\
        );

    \I__11972\ : LocalMux
    port map (
            O => \N__52694\,
            I => \N__52626\
        );

    \I__11971\ : LocalMux
    port map (
            O => \N__52691\,
            I => \N__52621\
        );

    \I__11970\ : LocalMux
    port map (
            O => \N__52688\,
            I => \N__52621\
        );

    \I__11969\ : LocalMux
    port map (
            O => \N__52685\,
            I => \N__52614\
        );

    \I__11968\ : LocalMux
    port map (
            O => \N__52682\,
            I => \N__52614\
        );

    \I__11967\ : LocalMux
    port map (
            O => \N__52677\,
            I => \N__52614\
        );

    \I__11966\ : InMux
    port map (
            O => \N__52676\,
            I => \N__52611\
        );

    \I__11965\ : InMux
    port map (
            O => \N__52675\,
            I => \N__52608\
        );

    \I__11964\ : InMux
    port map (
            O => \N__52674\,
            I => \N__52605\
        );

    \I__11963\ : InMux
    port map (
            O => \N__52673\,
            I => \N__52602\
        );

    \I__11962\ : InMux
    port map (
            O => \N__52672\,
            I => \N__52599\
        );

    \I__11961\ : LocalMux
    port map (
            O => \N__52669\,
            I => \N__52592\
        );

    \I__11960\ : LocalMux
    port map (
            O => \N__52666\,
            I => \N__52592\
        );

    \I__11959\ : LocalMux
    port map (
            O => \N__52663\,
            I => \N__52592\
        );

    \I__11958\ : Span4Mux_h
    port map (
            O => \N__52660\,
            I => \N__52585\
        );

    \I__11957\ : Span4Mux_v
    port map (
            O => \N__52657\,
            I => \N__52585\
        );

    \I__11956\ : Span4Mux_h
    port map (
            O => \N__52648\,
            I => \N__52585\
        );

    \I__11955\ : Span4Mux_h
    port map (
            O => \N__52643\,
            I => \N__52578\
        );

    \I__11954\ : Span4Mux_h
    port map (
            O => \N__52640\,
            I => \N__52578\
        );

    \I__11953\ : Span4Mux_h
    port map (
            O => \N__52637\,
            I => \N__52578\
        );

    \I__11952\ : LocalMux
    port map (
            O => \N__52634\,
            I => \N__52567\
        );

    \I__11951\ : LocalMux
    port map (
            O => \N__52631\,
            I => \N__52567\
        );

    \I__11950\ : Span4Mux_h
    port map (
            O => \N__52626\,
            I => \N__52567\
        );

    \I__11949\ : Span4Mux_v
    port map (
            O => \N__52621\,
            I => \N__52567\
        );

    \I__11948\ : Span4Mux_v
    port map (
            O => \N__52614\,
            I => \N__52567\
        );

    \I__11947\ : LocalMux
    port map (
            O => \N__52611\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11946\ : LocalMux
    port map (
            O => \N__52608\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11945\ : LocalMux
    port map (
            O => \N__52605\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11944\ : LocalMux
    port map (
            O => \N__52602\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11943\ : LocalMux
    port map (
            O => \N__52599\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11942\ : Odrv12
    port map (
            O => \N__52592\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11941\ : Odrv4
    port map (
            O => \N__52585\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11940\ : Odrv4
    port map (
            O => \N__52578\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11939\ : Odrv4
    port map (
            O => \N__52567\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\
        );

    \I__11938\ : CascadeMux
    port map (
            O => \N__52548\,
            I => \N__52545\
        );

    \I__11937\ : InMux
    port map (
            O => \N__52545\,
            I => \N__52542\
        );

    \I__11936\ : LocalMux
    port map (
            O => \N__52542\,
            I => \N__52539\
        );

    \I__11935\ : Span4Mux_v
    port map (
            O => \N__52539\,
            I => \N__52536\
        );

    \I__11934\ : Span4Mux_h
    port map (
            O => \N__52536\,
            I => \N__52533\
        );

    \I__11933\ : Sp12to4
    port map (
            O => \N__52533\,
            I => \N__52530\
        );

    \I__11932\ : Odrv12
    port map (
            O => \N__52530\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_25
        );

    \I__11931\ : InMux
    port map (
            O => \N__52527\,
            I => \N__52517\
        );

    \I__11930\ : InMux
    port map (
            O => \N__52526\,
            I => \N__52514\
        );

    \I__11929\ : InMux
    port map (
            O => \N__52525\,
            I => \N__52509\
        );

    \I__11928\ : InMux
    port map (
            O => \N__52524\,
            I => \N__52506\
        );

    \I__11927\ : InMux
    port map (
            O => \N__52523\,
            I => \N__52503\
        );

    \I__11926\ : InMux
    port map (
            O => \N__52522\,
            I => \N__52500\
        );

    \I__11925\ : InMux
    port map (
            O => \N__52521\,
            I => \N__52497\
        );

    \I__11924\ : InMux
    port map (
            O => \N__52520\,
            I => \N__52489\
        );

    \I__11923\ : LocalMux
    port map (
            O => \N__52517\,
            I => \N__52481\
        );

    \I__11922\ : LocalMux
    port map (
            O => \N__52514\,
            I => \N__52478\
        );

    \I__11921\ : InMux
    port map (
            O => \N__52513\,
            I => \N__52475\
        );

    \I__11920\ : InMux
    port map (
            O => \N__52512\,
            I => \N__52472\
        );

    \I__11919\ : LocalMux
    port map (
            O => \N__52509\,
            I => \N__52468\
        );

    \I__11918\ : LocalMux
    port map (
            O => \N__52506\,
            I => \N__52463\
        );

    \I__11917\ : LocalMux
    port map (
            O => \N__52503\,
            I => \N__52463\
        );

    \I__11916\ : LocalMux
    port map (
            O => \N__52500\,
            I => \N__52458\
        );

    \I__11915\ : LocalMux
    port map (
            O => \N__52497\,
            I => \N__52458\
        );

    \I__11914\ : InMux
    port map (
            O => \N__52496\,
            I => \N__52455\
        );

    \I__11913\ : InMux
    port map (
            O => \N__52495\,
            I => \N__52450\
        );

    \I__11912\ : InMux
    port map (
            O => \N__52494\,
            I => \N__52450\
        );

    \I__11911\ : InMux
    port map (
            O => \N__52493\,
            I => \N__52447\
        );

    \I__11910\ : InMux
    port map (
            O => \N__52492\,
            I => \N__52442\
        );

    \I__11909\ : LocalMux
    port map (
            O => \N__52489\,
            I => \N__52434\
        );

    \I__11908\ : InMux
    port map (
            O => \N__52488\,
            I => \N__52431\
        );

    \I__11907\ : InMux
    port map (
            O => \N__52487\,
            I => \N__52428\
        );

    \I__11906\ : InMux
    port map (
            O => \N__52486\,
            I => \N__52425\
        );

    \I__11905\ : InMux
    port map (
            O => \N__52485\,
            I => \N__52422\
        );

    \I__11904\ : InMux
    port map (
            O => \N__52484\,
            I => \N__52419\
        );

    \I__11903\ : Span4Mux_h
    port map (
            O => \N__52481\,
            I => \N__52410\
        );

    \I__11902\ : Span4Mux_h
    port map (
            O => \N__52478\,
            I => \N__52410\
        );

    \I__11901\ : LocalMux
    port map (
            O => \N__52475\,
            I => \N__52410\
        );

    \I__11900\ : LocalMux
    port map (
            O => \N__52472\,
            I => \N__52410\
        );

    \I__11899\ : InMux
    port map (
            O => \N__52471\,
            I => \N__52407\
        );

    \I__11898\ : Span4Mux_v
    port map (
            O => \N__52468\,
            I => \N__52404\
        );

    \I__11897\ : Span4Mux_v
    port map (
            O => \N__52463\,
            I => \N__52399\
        );

    \I__11896\ : Span4Mux_h
    port map (
            O => \N__52458\,
            I => \N__52399\
        );

    \I__11895\ : LocalMux
    port map (
            O => \N__52455\,
            I => \N__52396\
        );

    \I__11894\ : LocalMux
    port map (
            O => \N__52450\,
            I => \N__52391\
        );

    \I__11893\ : LocalMux
    port map (
            O => \N__52447\,
            I => \N__52391\
        );

    \I__11892\ : InMux
    port map (
            O => \N__52446\,
            I => \N__52388\
        );

    \I__11891\ : InMux
    port map (
            O => \N__52445\,
            I => \N__52385\
        );

    \I__11890\ : LocalMux
    port map (
            O => \N__52442\,
            I => \N__52382\
        );

    \I__11889\ : InMux
    port map (
            O => \N__52441\,
            I => \N__52378\
        );

    \I__11888\ : InMux
    port map (
            O => \N__52440\,
            I => \N__52375\
        );

    \I__11887\ : InMux
    port map (
            O => \N__52439\,
            I => \N__52372\
        );

    \I__11886\ : InMux
    port map (
            O => \N__52438\,
            I => \N__52367\
        );

    \I__11885\ : InMux
    port map (
            O => \N__52437\,
            I => \N__52364\
        );

    \I__11884\ : Span4Mux_h
    port map (
            O => \N__52434\,
            I => \N__52357\
        );

    \I__11883\ : LocalMux
    port map (
            O => \N__52431\,
            I => \N__52357\
        );

    \I__11882\ : LocalMux
    port map (
            O => \N__52428\,
            I => \N__52357\
        );

    \I__11881\ : LocalMux
    port map (
            O => \N__52425\,
            I => \N__52354\
        );

    \I__11880\ : LocalMux
    port map (
            O => \N__52422\,
            I => \N__52349\
        );

    \I__11879\ : LocalMux
    port map (
            O => \N__52419\,
            I => \N__52349\
        );

    \I__11878\ : Span4Mux_h
    port map (
            O => \N__52410\,
            I => \N__52344\
        );

    \I__11877\ : LocalMux
    port map (
            O => \N__52407\,
            I => \N__52344\
        );

    \I__11876\ : Span4Mux_h
    port map (
            O => \N__52404\,
            I => \N__52333\
        );

    \I__11875\ : Span4Mux_h
    port map (
            O => \N__52399\,
            I => \N__52333\
        );

    \I__11874\ : Span4Mux_v
    port map (
            O => \N__52396\,
            I => \N__52333\
        );

    \I__11873\ : Span4Mux_v
    port map (
            O => \N__52391\,
            I => \N__52333\
        );

    \I__11872\ : LocalMux
    port map (
            O => \N__52388\,
            I => \N__52333\
        );

    \I__11871\ : LocalMux
    port map (
            O => \N__52385\,
            I => \N__52330\
        );

    \I__11870\ : Span4Mux_h
    port map (
            O => \N__52382\,
            I => \N__52327\
        );

    \I__11869\ : InMux
    port map (
            O => \N__52381\,
            I => \N__52324\
        );

    \I__11868\ : LocalMux
    port map (
            O => \N__52378\,
            I => \N__52319\
        );

    \I__11867\ : LocalMux
    port map (
            O => \N__52375\,
            I => \N__52319\
        );

    \I__11866\ : LocalMux
    port map (
            O => \N__52372\,
            I => \N__52316\
        );

    \I__11865\ : InMux
    port map (
            O => \N__52371\,
            I => \N__52311\
        );

    \I__11864\ : InMux
    port map (
            O => \N__52370\,
            I => \N__52311\
        );

    \I__11863\ : LocalMux
    port map (
            O => \N__52367\,
            I => \N__52308\
        );

    \I__11862\ : LocalMux
    port map (
            O => \N__52364\,
            I => \N__52303\
        );

    \I__11861\ : Span4Mux_v
    port map (
            O => \N__52357\,
            I => \N__52303\
        );

    \I__11860\ : Span4Mux_h
    port map (
            O => \N__52354\,
            I => \N__52298\
        );

    \I__11859\ : Span4Mux_h
    port map (
            O => \N__52349\,
            I => \N__52298\
        );

    \I__11858\ : Span4Mux_v
    port map (
            O => \N__52344\,
            I => \N__52293\
        );

    \I__11857\ : Span4Mux_h
    port map (
            O => \N__52333\,
            I => \N__52293\
        );

    \I__11856\ : Span4Mux_h
    port map (
            O => \N__52330\,
            I => \N__52284\
        );

    \I__11855\ : Span4Mux_h
    port map (
            O => \N__52327\,
            I => \N__52284\
        );

    \I__11854\ : LocalMux
    port map (
            O => \N__52324\,
            I => \N__52284\
        );

    \I__11853\ : Span4Mux_v
    port map (
            O => \N__52319\,
            I => \N__52284\
        );

    \I__11852\ : Span4Mux_v
    port map (
            O => \N__52316\,
            I => \N__52279\
        );

    \I__11851\ : LocalMux
    port map (
            O => \N__52311\,
            I => \N__52279\
        );

    \I__11850\ : Span12Mux_v
    port map (
            O => \N__52308\,
            I => \N__52276\
        );

    \I__11849\ : Span4Mux_h
    port map (
            O => \N__52303\,
            I => \N__52271\
        );

    \I__11848\ : Span4Mux_v
    port map (
            O => \N__52298\,
            I => \N__52271\
        );

    \I__11847\ : Span4Mux_v
    port map (
            O => \N__52293\,
            I => \N__52268\
        );

    \I__11846\ : Span4Mux_v
    port map (
            O => \N__52284\,
            I => \N__52263\
        );

    \I__11845\ : Span4Mux_h
    port map (
            O => \N__52279\,
            I => \N__52263\
        );

    \I__11844\ : Odrv12
    port map (
            O => \N__52276\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314\
        );

    \I__11843\ : Odrv4
    port map (
            O => \N__52271\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314\
        );

    \I__11842\ : Odrv4
    port map (
            O => \N__52268\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314\
        );

    \I__11841\ : Odrv4
    port map (
            O => \N__52263\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314\
        );

    \I__11840\ : InMux
    port map (
            O => \N__52254\,
            I => \N__52251\
        );

    \I__11839\ : LocalMux
    port map (
            O => \N__52251\,
            I => \N__52248\
        );

    \I__11838\ : Span4Mux_h
    port map (
            O => \N__52248\,
            I => \N__52245\
        );

    \I__11837\ : Span4Mux_v
    port map (
            O => \N__52245\,
            I => \N__52242\
        );

    \I__11836\ : Odrv4
    port map (
            O => \N__52242\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_25\
        );

    \I__11835\ : CascadeMux
    port map (
            O => \N__52239\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_25_cascade_\
        );

    \I__11834\ : InMux
    port map (
            O => \N__52236\,
            I => \N__52228\
        );

    \I__11833\ : InMux
    port map (
            O => \N__52235\,
            I => \N__52224\
        );

    \I__11832\ : InMux
    port map (
            O => \N__52234\,
            I => \N__52217\
        );

    \I__11831\ : InMux
    port map (
            O => \N__52233\,
            I => \N__52210\
        );

    \I__11830\ : InMux
    port map (
            O => \N__52232\,
            I => \N__52207\
        );

    \I__11829\ : InMux
    port map (
            O => \N__52231\,
            I => \N__52200\
        );

    \I__11828\ : LocalMux
    port map (
            O => \N__52228\,
            I => \N__52195\
        );

    \I__11827\ : InMux
    port map (
            O => \N__52227\,
            I => \N__52192\
        );

    \I__11826\ : LocalMux
    port map (
            O => \N__52224\,
            I => \N__52188\
        );

    \I__11825\ : InMux
    port map (
            O => \N__52223\,
            I => \N__52183\
        );

    \I__11824\ : InMux
    port map (
            O => \N__52222\,
            I => \N__52179\
        );

    \I__11823\ : InMux
    port map (
            O => \N__52221\,
            I => \N__52176\
        );

    \I__11822\ : InMux
    port map (
            O => \N__52220\,
            I => \N__52173\
        );

    \I__11821\ : LocalMux
    port map (
            O => \N__52217\,
            I => \N__52170\
        );

    \I__11820\ : InMux
    port map (
            O => \N__52216\,
            I => \N__52167\
        );

    \I__11819\ : InMux
    port map (
            O => \N__52215\,
            I => \N__52164\
        );

    \I__11818\ : InMux
    port map (
            O => \N__52214\,
            I => \N__52161\
        );

    \I__11817\ : InMux
    port map (
            O => \N__52213\,
            I => \N__52158\
        );

    \I__11816\ : LocalMux
    port map (
            O => \N__52210\,
            I => \N__52153\
        );

    \I__11815\ : LocalMux
    port map (
            O => \N__52207\,
            I => \N__52153\
        );

    \I__11814\ : InMux
    port map (
            O => \N__52206\,
            I => \N__52150\
        );

    \I__11813\ : InMux
    port map (
            O => \N__52205\,
            I => \N__52147\
        );

    \I__11812\ : InMux
    port map (
            O => \N__52204\,
            I => \N__52142\
        );

    \I__11811\ : InMux
    port map (
            O => \N__52203\,
            I => \N__52139\
        );

    \I__11810\ : LocalMux
    port map (
            O => \N__52200\,
            I => \N__52136\
        );

    \I__11809\ : InMux
    port map (
            O => \N__52199\,
            I => \N__52133\
        );

    \I__11808\ : InMux
    port map (
            O => \N__52198\,
            I => \N__52130\
        );

    \I__11807\ : Span4Mux_h
    port map (
            O => \N__52195\,
            I => \N__52125\
        );

    \I__11806\ : LocalMux
    port map (
            O => \N__52192\,
            I => \N__52125\
        );

    \I__11805\ : InMux
    port map (
            O => \N__52191\,
            I => \N__52119\
        );

    \I__11804\ : Span4Mux_v
    port map (
            O => \N__52188\,
            I => \N__52116\
        );

    \I__11803\ : InMux
    port map (
            O => \N__52187\,
            I => \N__52113\
        );

    \I__11802\ : InMux
    port map (
            O => \N__52186\,
            I => \N__52110\
        );

    \I__11801\ : LocalMux
    port map (
            O => \N__52183\,
            I => \N__52107\
        );

    \I__11800\ : InMux
    port map (
            O => \N__52182\,
            I => \N__52104\
        );

    \I__11799\ : LocalMux
    port map (
            O => \N__52179\,
            I => \N__52099\
        );

    \I__11798\ : LocalMux
    port map (
            O => \N__52176\,
            I => \N__52099\
        );

    \I__11797\ : LocalMux
    port map (
            O => \N__52173\,
            I => \N__52090\
        );

    \I__11796\ : Span4Mux_h
    port map (
            O => \N__52170\,
            I => \N__52090\
        );

    \I__11795\ : LocalMux
    port map (
            O => \N__52167\,
            I => \N__52090\
        );

    \I__11794\ : LocalMux
    port map (
            O => \N__52164\,
            I => \N__52090\
        );

    \I__11793\ : LocalMux
    port map (
            O => \N__52161\,
            I => \N__52087\
        );

    \I__11792\ : LocalMux
    port map (
            O => \N__52158\,
            I => \N__52080\
        );

    \I__11791\ : Span4Mux_v
    port map (
            O => \N__52153\,
            I => \N__52080\
        );

    \I__11790\ : LocalMux
    port map (
            O => \N__52150\,
            I => \N__52080\
        );

    \I__11789\ : LocalMux
    port map (
            O => \N__52147\,
            I => \N__52077\
        );

    \I__11788\ : InMux
    port map (
            O => \N__52146\,
            I => \N__52074\
        );

    \I__11787\ : InMux
    port map (
            O => \N__52145\,
            I => \N__52071\
        );

    \I__11786\ : LocalMux
    port map (
            O => \N__52142\,
            I => \N__52066\
        );

    \I__11785\ : LocalMux
    port map (
            O => \N__52139\,
            I => \N__52066\
        );

    \I__11784\ : Span4Mux_h
    port map (
            O => \N__52136\,
            I => \N__52061\
        );

    \I__11783\ : LocalMux
    port map (
            O => \N__52133\,
            I => \N__52061\
        );

    \I__11782\ : LocalMux
    port map (
            O => \N__52130\,
            I => \N__52058\
        );

    \I__11781\ : Span4Mux_h
    port map (
            O => \N__52125\,
            I => \N__52055\
        );

    \I__11780\ : InMux
    port map (
            O => \N__52124\,
            I => \N__52051\
        );

    \I__11779\ : InMux
    port map (
            O => \N__52123\,
            I => \N__52048\
        );

    \I__11778\ : InMux
    port map (
            O => \N__52122\,
            I => \N__52045\
        );

    \I__11777\ : LocalMux
    port map (
            O => \N__52119\,
            I => \N__52038\
        );

    \I__11776\ : Sp12to4
    port map (
            O => \N__52116\,
            I => \N__52038\
        );

    \I__11775\ : LocalMux
    port map (
            O => \N__52113\,
            I => \N__52038\
        );

    \I__11774\ : LocalMux
    port map (
            O => \N__52110\,
            I => \N__52027\
        );

    \I__11773\ : Span4Mux_v
    port map (
            O => \N__52107\,
            I => \N__52027\
        );

    \I__11772\ : LocalMux
    port map (
            O => \N__52104\,
            I => \N__52027\
        );

    \I__11771\ : Span4Mux_h
    port map (
            O => \N__52099\,
            I => \N__52027\
        );

    \I__11770\ : Span4Mux_v
    port map (
            O => \N__52090\,
            I => \N__52027\
        );

    \I__11769\ : Span4Mux_h
    port map (
            O => \N__52087\,
            I => \N__52020\
        );

    \I__11768\ : Span4Mux_h
    port map (
            O => \N__52080\,
            I => \N__52020\
        );

    \I__11767\ : Span4Mux_h
    port map (
            O => \N__52077\,
            I => \N__52020\
        );

    \I__11766\ : LocalMux
    port map (
            O => \N__52074\,
            I => \N__52017\
        );

    \I__11765\ : LocalMux
    port map (
            O => \N__52071\,
            I => \N__52006\
        );

    \I__11764\ : Span4Mux_h
    port map (
            O => \N__52066\,
            I => \N__52006\
        );

    \I__11763\ : Span4Mux_h
    port map (
            O => \N__52061\,
            I => \N__52006\
        );

    \I__11762\ : Span4Mux_h
    port map (
            O => \N__52058\,
            I => \N__52006\
        );

    \I__11761\ : Span4Mux_h
    port map (
            O => \N__52055\,
            I => \N__52006\
        );

    \I__11760\ : InMux
    port map (
            O => \N__52054\,
            I => \N__52003\
        );

    \I__11759\ : LocalMux
    port map (
            O => \N__52051\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11758\ : LocalMux
    port map (
            O => \N__52048\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11757\ : LocalMux
    port map (
            O => \N__52045\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11756\ : Odrv12
    port map (
            O => \N__52038\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11755\ : Odrv4
    port map (
            O => \N__52027\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11754\ : Odrv4
    port map (
            O => \N__52020\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11753\ : Odrv4
    port map (
            O => \N__52017\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11752\ : Odrv4
    port map (
            O => \N__52006\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11751\ : LocalMux
    port map (
            O => \N__52003\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\
        );

    \I__11750\ : InMux
    port map (
            O => \N__51984\,
            I => \N__51981\
        );

    \I__11749\ : LocalMux
    port map (
            O => \N__51981\,
            I => \N__51978\
        );

    \I__11748\ : Odrv12
    port map (
            O => \N__51978\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_25\
        );

    \I__11747\ : InMux
    port map (
            O => \N__51975\,
            I => \N__51972\
        );

    \I__11746\ : LocalMux
    port map (
            O => \N__51972\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_25\
        );

    \I__11745\ : CascadeMux
    port map (
            O => \N__51969\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_25_cascade_\
        );

    \I__11744\ : InMux
    port map (
            O => \N__51966\,
            I => \N__51963\
        );

    \I__11743\ : LocalMux
    port map (
            O => \N__51963\,
            I => \N__51960\
        );

    \I__11742\ : Span4Mux_h
    port map (
            O => \N__51960\,
            I => \N__51957\
        );

    \I__11741\ : Span4Mux_h
    port map (
            O => \N__51957\,
            I => \N__51954\
        );

    \I__11740\ : Odrv4
    port map (
            O => \N__51954\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_665\
        );

    \I__11739\ : CascadeMux
    port map (
            O => \N__51951\,
            I => \N__51947\
        );

    \I__11738\ : InMux
    port map (
            O => \N__51950\,
            I => \N__51943\
        );

    \I__11737\ : InMux
    port map (
            O => \N__51947\,
            I => \N__51940\
        );

    \I__11736\ : CascadeMux
    port map (
            O => \N__51946\,
            I => \N__51937\
        );

    \I__11735\ : LocalMux
    port map (
            O => \N__51943\,
            I => \N__51931\
        );

    \I__11734\ : LocalMux
    port map (
            O => \N__51940\,
            I => \N__51931\
        );

    \I__11733\ : InMux
    port map (
            O => \N__51937\,
            I => \N__51928\
        );

    \I__11732\ : InMux
    port map (
            O => \N__51936\,
            I => \N__51916\
        );

    \I__11731\ : Span4Mux_v
    port map (
            O => \N__51931\,
            I => \N__51910\
        );

    \I__11730\ : LocalMux
    port map (
            O => \N__51928\,
            I => \N__51910\
        );

    \I__11729\ : InMux
    port map (
            O => \N__51927\,
            I => \N__51907\
        );

    \I__11728\ : CascadeMux
    port map (
            O => \N__51926\,
            I => \N__51899\
        );

    \I__11727\ : InMux
    port map (
            O => \N__51925\,
            I => \N__51896\
        );

    \I__11726\ : InMux
    port map (
            O => \N__51924\,
            I => \N__51893\
        );

    \I__11725\ : InMux
    port map (
            O => \N__51923\,
            I => \N__51887\
        );

    \I__11724\ : InMux
    port map (
            O => \N__51922\,
            I => \N__51884\
        );

    \I__11723\ : InMux
    port map (
            O => \N__51921\,
            I => \N__51881\
        );

    \I__11722\ : InMux
    port map (
            O => \N__51920\,
            I => \N__51878\
        );

    \I__11721\ : InMux
    port map (
            O => \N__51919\,
            I => \N__51875\
        );

    \I__11720\ : LocalMux
    port map (
            O => \N__51916\,
            I => \N__51872\
        );

    \I__11719\ : CascadeMux
    port map (
            O => \N__51915\,
            I => \N__51868\
        );

    \I__11718\ : Span4Mux_h
    port map (
            O => \N__51910\,
            I => \N__51861\
        );

    \I__11717\ : LocalMux
    port map (
            O => \N__51907\,
            I => \N__51861\
        );

    \I__11716\ : InMux
    port map (
            O => \N__51906\,
            I => \N__51856\
        );

    \I__11715\ : CascadeMux
    port map (
            O => \N__51905\,
            I => \N__51853\
        );

    \I__11714\ : InMux
    port map (
            O => \N__51904\,
            I => \N__51850\
        );

    \I__11713\ : InMux
    port map (
            O => \N__51903\,
            I => \N__51847\
        );

    \I__11712\ : InMux
    port map (
            O => \N__51902\,
            I => \N__51843\
        );

    \I__11711\ : InMux
    port map (
            O => \N__51899\,
            I => \N__51840\
        );

    \I__11710\ : LocalMux
    port map (
            O => \N__51896\,
            I => \N__51837\
        );

    \I__11709\ : LocalMux
    port map (
            O => \N__51893\,
            I => \N__51834\
        );

    \I__11708\ : InMux
    port map (
            O => \N__51892\,
            I => \N__51831\
        );

    \I__11707\ : InMux
    port map (
            O => \N__51891\,
            I => \N__51828\
        );

    \I__11706\ : InMux
    port map (
            O => \N__51890\,
            I => \N__51825\
        );

    \I__11705\ : LocalMux
    port map (
            O => \N__51887\,
            I => \N__51821\
        );

    \I__11704\ : LocalMux
    port map (
            O => \N__51884\,
            I => \N__51814\
        );

    \I__11703\ : LocalMux
    port map (
            O => \N__51881\,
            I => \N__51814\
        );

    \I__11702\ : LocalMux
    port map (
            O => \N__51878\,
            I => \N__51814\
        );

    \I__11701\ : LocalMux
    port map (
            O => \N__51875\,
            I => \N__51809\
        );

    \I__11700\ : Span4Mux_h
    port map (
            O => \N__51872\,
            I => \N__51809\
        );

    \I__11699\ : InMux
    port map (
            O => \N__51871\,
            I => \N__51804\
        );

    \I__11698\ : InMux
    port map (
            O => \N__51868\,
            I => \N__51804\
        );

    \I__11697\ : CascadeMux
    port map (
            O => \N__51867\,
            I => \N__51801\
        );

    \I__11696\ : InMux
    port map (
            O => \N__51866\,
            I => \N__51798\
        );

    \I__11695\ : Span4Mux_v
    port map (
            O => \N__51861\,
            I => \N__51795\
        );

    \I__11694\ : InMux
    port map (
            O => \N__51860\,
            I => \N__51792\
        );

    \I__11693\ : InMux
    port map (
            O => \N__51859\,
            I => \N__51787\
        );

    \I__11692\ : LocalMux
    port map (
            O => \N__51856\,
            I => \N__51784\
        );

    \I__11691\ : InMux
    port map (
            O => \N__51853\,
            I => \N__51781\
        );

    \I__11690\ : LocalMux
    port map (
            O => \N__51850\,
            I => \N__51776\
        );

    \I__11689\ : LocalMux
    port map (
            O => \N__51847\,
            I => \N__51776\
        );

    \I__11688\ : InMux
    port map (
            O => \N__51846\,
            I => \N__51773\
        );

    \I__11687\ : LocalMux
    port map (
            O => \N__51843\,
            I => \N__51770\
        );

    \I__11686\ : LocalMux
    port map (
            O => \N__51840\,
            I => \N__51765\
        );

    \I__11685\ : Span4Mux_h
    port map (
            O => \N__51837\,
            I => \N__51765\
        );

    \I__11684\ : Span4Mux_v
    port map (
            O => \N__51834\,
            I => \N__51760\
        );

    \I__11683\ : LocalMux
    port map (
            O => \N__51831\,
            I => \N__51760\
        );

    \I__11682\ : LocalMux
    port map (
            O => \N__51828\,
            I => \N__51755\
        );

    \I__11681\ : LocalMux
    port map (
            O => \N__51825\,
            I => \N__51755\
        );

    \I__11680\ : InMux
    port map (
            O => \N__51824\,
            I => \N__51752\
        );

    \I__11679\ : Span4Mux_h
    port map (
            O => \N__51821\,
            I => \N__51743\
        );

    \I__11678\ : Span4Mux_v
    port map (
            O => \N__51814\,
            I => \N__51743\
        );

    \I__11677\ : Span4Mux_h
    port map (
            O => \N__51809\,
            I => \N__51743\
        );

    \I__11676\ : LocalMux
    port map (
            O => \N__51804\,
            I => \N__51743\
        );

    \I__11675\ : InMux
    port map (
            O => \N__51801\,
            I => \N__51740\
        );

    \I__11674\ : LocalMux
    port map (
            O => \N__51798\,
            I => \N__51733\
        );

    \I__11673\ : Sp12to4
    port map (
            O => \N__51795\,
            I => \N__51733\
        );

    \I__11672\ : LocalMux
    port map (
            O => \N__51792\,
            I => \N__51733\
        );

    \I__11671\ : InMux
    port map (
            O => \N__51791\,
            I => \N__51730\
        );

    \I__11670\ : InMux
    port map (
            O => \N__51790\,
            I => \N__51727\
        );

    \I__11669\ : LocalMux
    port map (
            O => \N__51787\,
            I => \N__51718\
        );

    \I__11668\ : Span4Mux_v
    port map (
            O => \N__51784\,
            I => \N__51718\
        );

    \I__11667\ : LocalMux
    port map (
            O => \N__51781\,
            I => \N__51718\
        );

    \I__11666\ : Span4Mux_v
    port map (
            O => \N__51776\,
            I => \N__51718\
        );

    \I__11665\ : LocalMux
    port map (
            O => \N__51773\,
            I => \N__51707\
        );

    \I__11664\ : Span4Mux_v
    port map (
            O => \N__51770\,
            I => \N__51707\
        );

    \I__11663\ : Span4Mux_v
    port map (
            O => \N__51765\,
            I => \N__51707\
        );

    \I__11662\ : Span4Mux_h
    port map (
            O => \N__51760\,
            I => \N__51707\
        );

    \I__11661\ : Span4Mux_v
    port map (
            O => \N__51755\,
            I => \N__51707\
        );

    \I__11660\ : LocalMux
    port map (
            O => \N__51752\,
            I => \N__51702\
        );

    \I__11659\ : Span4Mux_h
    port map (
            O => \N__51743\,
            I => \N__51702\
        );

    \I__11658\ : LocalMux
    port map (
            O => \N__51740\,
            I => \N__51697\
        );

    \I__11657\ : Span12Mux_h
    port map (
            O => \N__51733\,
            I => \N__51697\
        );

    \I__11656\ : LocalMux
    port map (
            O => \N__51730\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\
        );

    \I__11655\ : LocalMux
    port map (
            O => \N__51727\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\
        );

    \I__11654\ : Odrv4
    port map (
            O => \N__51718\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\
        );

    \I__11653\ : Odrv4
    port map (
            O => \N__51707\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\
        );

    \I__11652\ : Odrv4
    port map (
            O => \N__51702\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\
        );

    \I__11651\ : Odrv12
    port map (
            O => \N__51697\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\
        );

    \I__11650\ : CascadeMux
    port map (
            O => \N__51684\,
            I => \N__51681\
        );

    \I__11649\ : InMux
    port map (
            O => \N__51681\,
            I => \N__51678\
        );

    \I__11648\ : LocalMux
    port map (
            O => \N__51678\,
            I => \N__51675\
        );

    \I__11647\ : Odrv4
    port map (
            O => \N__51675\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_25\
        );

    \I__11646\ : InMux
    port map (
            O => \N__51672\,
            I => \N__51669\
        );

    \I__11645\ : LocalMux
    port map (
            O => \N__51669\,
            I => \N__51666\
        );

    \I__11644\ : Odrv12
    port map (
            O => \N__51666\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_25\
        );

    \I__11643\ : InMux
    port map (
            O => \N__51663\,
            I => \N__51660\
        );

    \I__11642\ : LocalMux
    port map (
            O => \N__51660\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_25\
        );

    \I__11641\ : InMux
    port map (
            O => \N__51657\,
            I => \N__51653\
        );

    \I__11640\ : CascadeMux
    port map (
            O => \N__51656\,
            I => \N__51649\
        );

    \I__11639\ : LocalMux
    port map (
            O => \N__51653\,
            I => \N__51646\
        );

    \I__11638\ : InMux
    port map (
            O => \N__51652\,
            I => \N__51643\
        );

    \I__11637\ : InMux
    port map (
            O => \N__51649\,
            I => \N__51640\
        );

    \I__11636\ : Span4Mux_h
    port map (
            O => \N__51646\,
            I => \N__51637\
        );

    \I__11635\ : LocalMux
    port map (
            O => \N__51643\,
            I => \N__51634\
        );

    \I__11634\ : LocalMux
    port map (
            O => \N__51640\,
            I => \N__51631\
        );

    \I__11633\ : Odrv4
    port map (
            O => \N__51637\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_16
        );

    \I__11632\ : Odrv4
    port map (
            O => \N__51634\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_16
        );

    \I__11631\ : Odrv4
    port map (
            O => \N__51631\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_16
        );

    \I__11630\ : InMux
    port map (
            O => \N__51624\,
            I => \N__51621\
        );

    \I__11629\ : LocalMux
    port map (
            O => \N__51621\,
            I => \N__51617\
        );

    \I__11628\ : CascadeMux
    port map (
            O => \N__51620\,
            I => \N__51614\
        );

    \I__11627\ : Span4Mux_v
    port map (
            O => \N__51617\,
            I => \N__51611\
        );

    \I__11626\ : InMux
    port map (
            O => \N__51614\,
            I => \N__51607\
        );

    \I__11625\ : Span4Mux_h
    port map (
            O => \N__51611\,
            I => \N__51604\
        );

    \I__11624\ : InMux
    port map (
            O => \N__51610\,
            I => \N__51601\
        );

    \I__11623\ : LocalMux
    port map (
            O => \N__51607\,
            I => \N__51598\
        );

    \I__11622\ : Span4Mux_h
    port map (
            O => \N__51604\,
            I => \N__51591\
        );

    \I__11621\ : LocalMux
    port map (
            O => \N__51601\,
            I => \N__51591\
        );

    \I__11620\ : Span4Mux_h
    port map (
            O => \N__51598\,
            I => \N__51591\
        );

    \I__11619\ : Odrv4
    port map (
            O => \N__51591\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_17
        );

    \I__11618\ : CascadeMux
    port map (
            O => \N__51588\,
            I => \N__51583\
        );

    \I__11617\ : InMux
    port map (
            O => \N__51587\,
            I => \N__51580\
        );

    \I__11616\ : InMux
    port map (
            O => \N__51586\,
            I => \N__51577\
        );

    \I__11615\ : InMux
    port map (
            O => \N__51583\,
            I => \N__51574\
        );

    \I__11614\ : LocalMux
    port map (
            O => \N__51580\,
            I => \N__51571\
        );

    \I__11613\ : LocalMux
    port map (
            O => \N__51577\,
            I => \N__51568\
        );

    \I__11612\ : LocalMux
    port map (
            O => \N__51574\,
            I => \N__51565\
        );

    \I__11611\ : Span4Mux_h
    port map (
            O => \N__51571\,
            I => \N__51562\
        );

    \I__11610\ : Odrv12
    port map (
            O => \N__51568\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_17
        );

    \I__11609\ : Odrv4
    port map (
            O => \N__51565\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_17
        );

    \I__11608\ : Odrv4
    port map (
            O => \N__51562\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_17
        );

    \I__11607\ : CascadeMux
    port map (
            O => \N__51555\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_17_cascade_\
        );

    \I__11606\ : InMux
    port map (
            O => \N__51552\,
            I => \N__51549\
        );

    \I__11605\ : LocalMux
    port map (
            O => \N__51549\,
            I => \N__51546\
        );

    \I__11604\ : Odrv4
    port map (
            O => \N__51546\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_17\
        );

    \I__11603\ : InMux
    port map (
            O => \N__51543\,
            I => \N__51540\
        );

    \I__11602\ : LocalMux
    port map (
            O => \N__51540\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_19\
        );

    \I__11601\ : CascadeMux
    port map (
            O => \N__51537\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HHZ0Z5_cascade_\
        );

    \I__11600\ : InMux
    port map (
            O => \N__51534\,
            I => \N__51531\
        );

    \I__11599\ : LocalMux
    port map (
            O => \N__51531\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19\
        );

    \I__11598\ : CascadeMux
    port map (
            O => \N__51528\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19_cascade_\
        );

    \I__11597\ : InMux
    port map (
            O => \N__51525\,
            I => \N__51522\
        );

    \I__11596\ : LocalMux
    port map (
            O => \N__51522\,
            I => \N__51519\
        );

    \I__11595\ : Span4Mux_h
    port map (
            O => \N__51519\,
            I => \N__51516\
        );

    \I__11594\ : Span4Mux_h
    port map (
            O => \N__51516\,
            I => \N__51513\
        );

    \I__11593\ : Odrv4
    port map (
            O => \N__51513\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_19\
        );

    \I__11592\ : InMux
    port map (
            O => \N__51510\,
            I => \N__51507\
        );

    \I__11591\ : LocalMux
    port map (
            O => \N__51507\,
            I => \N__51502\
        );

    \I__11590\ : CascadeMux
    port map (
            O => \N__51506\,
            I => \N__51499\
        );

    \I__11589\ : CascadeMux
    port map (
            O => \N__51505\,
            I => \N__51496\
        );

    \I__11588\ : Span4Mux_v
    port map (
            O => \N__51502\,
            I => \N__51493\
        );

    \I__11587\ : InMux
    port map (
            O => \N__51499\,
            I => \N__51490\
        );

    \I__11586\ : InMux
    port map (
            O => \N__51496\,
            I => \N__51487\
        );

    \I__11585\ : Span4Mux_h
    port map (
            O => \N__51493\,
            I => \N__51482\
        );

    \I__11584\ : LocalMux
    port map (
            O => \N__51490\,
            I => \N__51482\
        );

    \I__11583\ : LocalMux
    port map (
            O => \N__51487\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_19
        );

    \I__11582\ : Odrv4
    port map (
            O => \N__51482\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_19
        );

    \I__11581\ : InMux
    port map (
            O => \N__51477\,
            I => \N__51473\
        );

    \I__11580\ : InMux
    port map (
            O => \N__51476\,
            I => \N__51470\
        );

    \I__11579\ : LocalMux
    port map (
            O => \N__51473\,
            I => \N__51467\
        );

    \I__11578\ : LocalMux
    port map (
            O => \N__51470\,
            I => \N__51464\
        );

    \I__11577\ : Span4Mux_h
    port map (
            O => \N__51467\,
            I => \N__51460\
        );

    \I__11576\ : Span4Mux_h
    port map (
            O => \N__51464\,
            I => \N__51457\
        );

    \I__11575\ : InMux
    port map (
            O => \N__51463\,
            I => \N__51454\
        );

    \I__11574\ : Odrv4
    port map (
            O => \N__51460\,
            I => cemf_module_64ch_ctrl_inst1_data_config_19
        );

    \I__11573\ : Odrv4
    port map (
            O => \N__51457\,
            I => cemf_module_64ch_ctrl_inst1_data_config_19
        );

    \I__11572\ : LocalMux
    port map (
            O => \N__51454\,
            I => cemf_module_64ch_ctrl_inst1_data_config_19
        );

    \I__11571\ : CascadeMux
    port map (
            O => \N__51447\,
            I => \N__51444\
        );

    \I__11570\ : InMux
    port map (
            O => \N__51444\,
            I => \N__51441\
        );

    \I__11569\ : LocalMux
    port map (
            O => \N__51441\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_19\
        );

    \I__11568\ : InMux
    port map (
            O => \N__51438\,
            I => \N__51435\
        );

    \I__11567\ : LocalMux
    port map (
            O => \N__51435\,
            I => \N__51431\
        );

    \I__11566\ : CascadeMux
    port map (
            O => \N__51434\,
            I => \N__51427\
        );

    \I__11565\ : Span4Mux_h
    port map (
            O => \N__51431\,
            I => \N__51424\
        );

    \I__11564\ : CascadeMux
    port map (
            O => \N__51430\,
            I => \N__51421\
        );

    \I__11563\ : InMux
    port map (
            O => \N__51427\,
            I => \N__51418\
        );

    \I__11562\ : Span4Mux_h
    port map (
            O => \N__51424\,
            I => \N__51415\
        );

    \I__11561\ : InMux
    port map (
            O => \N__51421\,
            I => \N__51412\
        );

    \I__11560\ : LocalMux
    port map (
            O => \N__51418\,
            I => \N__51409\
        );

    \I__11559\ : Odrv4
    port map (
            O => \N__51415\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_18
        );

    \I__11558\ : LocalMux
    port map (
            O => \N__51412\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_18
        );

    \I__11557\ : Odrv4
    port map (
            O => \N__51409\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_18
        );

    \I__11556\ : InMux
    port map (
            O => \N__51402\,
            I => \N__51399\
        );

    \I__11555\ : LocalMux
    port map (
            O => \N__51399\,
            I => \N__51396\
        );

    \I__11554\ : Span4Mux_v
    port map (
            O => \N__51396\,
            I => \N__51392\
        );

    \I__11553\ : InMux
    port map (
            O => \N__51395\,
            I => \N__51389\
        );

    \I__11552\ : Span4Mux_h
    port map (
            O => \N__51392\,
            I => \N__51386\
        );

    \I__11551\ : LocalMux
    port map (
            O => \N__51389\,
            I => \N__51383\
        );

    \I__11550\ : Span4Mux_h
    port map (
            O => \N__51386\,
            I => \N__51377\
        );

    \I__11549\ : Span4Mux_v
    port map (
            O => \N__51383\,
            I => \N__51377\
        );

    \I__11548\ : InMux
    port map (
            O => \N__51382\,
            I => \N__51374\
        );

    \I__11547\ : Odrv4
    port map (
            O => \N__51377\,
            I => cemf_module_64ch_ctrl_inst1_data_config_18
        );

    \I__11546\ : LocalMux
    port map (
            O => \N__51374\,
            I => cemf_module_64ch_ctrl_inst1_data_config_18
        );

    \I__11545\ : InMux
    port map (
            O => \N__51369\,
            I => \N__51365\
        );

    \I__11544\ : InMux
    port map (
            O => \N__51368\,
            I => \N__51361\
        );

    \I__11543\ : LocalMux
    port map (
            O => \N__51365\,
            I => \N__51358\
        );

    \I__11542\ : InMux
    port map (
            O => \N__51364\,
            I => \N__51355\
        );

    \I__11541\ : LocalMux
    port map (
            O => \N__51361\,
            I => \N__51352\
        );

    \I__11540\ : Span4Mux_v
    port map (
            O => \N__51358\,
            I => \N__51347\
        );

    \I__11539\ : LocalMux
    port map (
            O => \N__51355\,
            I => \N__51347\
        );

    \I__11538\ : Odrv4
    port map (
            O => \N__51352\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_18
        );

    \I__11537\ : Odrv4
    port map (
            O => \N__51347\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_18
        );

    \I__11536\ : CascadeMux
    port map (
            O => \N__51342\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_18_cascade_\
        );

    \I__11535\ : InMux
    port map (
            O => \N__51339\,
            I => \N__51336\
        );

    \I__11534\ : LocalMux
    port map (
            O => \N__51336\,
            I => \N__51333\
        );

    \I__11533\ : Span4Mux_h
    port map (
            O => \N__51333\,
            I => \N__51330\
        );

    \I__11532\ : Odrv4
    port map (
            O => \N__51330\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_18\
        );

    \I__11531\ : CascadeMux
    port map (
            O => \N__51327\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGHZ0Z5_cascade_\
        );

    \I__11530\ : InMux
    port map (
            O => \N__51324\,
            I => \N__51321\
        );

    \I__11529\ : LocalMux
    port map (
            O => \N__51321\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18\
        );

    \I__11528\ : CascadeMux
    port map (
            O => \N__51318\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18_cascade_\
        );

    \I__11527\ : InMux
    port map (
            O => \N__51315\,
            I => \N__51312\
        );

    \I__11526\ : LocalMux
    port map (
            O => \N__51312\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_18\
        );

    \I__11525\ : InMux
    port map (
            O => \N__51309\,
            I => \N__51306\
        );

    \I__11524\ : LocalMux
    port map (
            O => \N__51306\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_1\
        );

    \I__11523\ : InMux
    port map (
            O => \N__51303\,
            I => \N__51300\
        );

    \I__11522\ : LocalMux
    port map (
            O => \N__51300\,
            I => \N__51296\
        );

    \I__11521\ : InMux
    port map (
            O => \N__51299\,
            I => \N__51293\
        );

    \I__11520\ : Span12Mux_v
    port map (
            O => \N__51296\,
            I => \N__51290\
        );

    \I__11519\ : LocalMux
    port map (
            O => \N__51293\,
            I => \I2C_top_level_inst1.s_r_w\
        );

    \I__11518\ : Odrv12
    port map (
            O => \N__51290\,
            I => \I2C_top_level_inst1.s_r_w\
        );

    \I__11517\ : InMux
    port map (
            O => \N__51285\,
            I => \N__51282\
        );

    \I__11516\ : LocalMux
    port map (
            O => \N__51282\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_0\
        );

    \I__11515\ : InMux
    port map (
            O => \N__51279\,
            I => \N__51276\
        );

    \I__11514\ : LocalMux
    port map (
            O => \N__51276\,
            I => \N__51273\
        );

    \I__11513\ : Span4Mux_v
    port map (
            O => \N__51273\,
            I => \N__51270\
        );

    \I__11512\ : Span4Mux_h
    port map (
            O => \N__51270\,
            I => \N__51267\
        );

    \I__11511\ : Odrv4
    port map (
            O => \N__51267\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_27\
        );

    \I__11510\ : InMux
    port map (
            O => \N__51264\,
            I => \N__51261\
        );

    \I__11509\ : LocalMux
    port map (
            O => \N__51261\,
            I => \N__51258\
        );

    \I__11508\ : Span4Mux_h
    port map (
            O => \N__51258\,
            I => \N__51255\
        );

    \I__11507\ : Odrv4
    port map (
            O => \N__51255\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_29\
        );

    \I__11506\ : InMux
    port map (
            O => \N__51252\,
            I => \N__51248\
        );

    \I__11505\ : InMux
    port map (
            O => \N__51251\,
            I => \N__51245\
        );

    \I__11504\ : LocalMux
    port map (
            O => \N__51248\,
            I => \N__51242\
        );

    \I__11503\ : LocalMux
    port map (
            O => \N__51245\,
            I => \N__51238\
        );

    \I__11502\ : Span4Mux_v
    port map (
            O => \N__51242\,
            I => \N__51235\
        );

    \I__11501\ : InMux
    port map (
            O => \N__51241\,
            I => \N__51232\
        );

    \I__11500\ : Span4Mux_v
    port map (
            O => \N__51238\,
            I => \N__51229\
        );

    \I__11499\ : Span4Mux_h
    port map (
            O => \N__51235\,
            I => \N__51224\
        );

    \I__11498\ : LocalMux
    port map (
            O => \N__51232\,
            I => \N__51224\
        );

    \I__11497\ : Span4Mux_h
    port map (
            O => \N__51229\,
            I => \N__51221\
        );

    \I__11496\ : Span4Mux_v
    port map (
            O => \N__51224\,
            I => \N__51218\
        );

    \I__11495\ : Odrv4
    port map (
            O => \N__51221\,
            I => cemf_module_64ch_ctrl_inst1_data_config_23
        );

    \I__11494\ : Odrv4
    port map (
            O => \N__51218\,
            I => cemf_module_64ch_ctrl_inst1_data_config_23
        );

    \I__11493\ : InMux
    port map (
            O => \N__51213\,
            I => \N__51210\
        );

    \I__11492\ : LocalMux
    port map (
            O => \N__51210\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_1\
        );

    \I__11491\ : IoInMux
    port map (
            O => \N__51207\,
            I => \N__51203\
        );

    \I__11490\ : InMux
    port map (
            O => \N__51206\,
            I => \N__51200\
        );

    \I__11489\ : LocalMux
    port map (
            O => \N__51203\,
            I => \N__51197\
        );

    \I__11488\ : LocalMux
    port map (
            O => \N__51200\,
            I => \N__51194\
        );

    \I__11487\ : IoSpan4Mux
    port map (
            O => \N__51197\,
            I => \N__51191\
        );

    \I__11486\ : Span4Mux_h
    port map (
            O => \N__51194\,
            I => \N__51187\
        );

    \I__11485\ : Span4Mux_s2_v
    port map (
            O => \N__51191\,
            I => \N__51183\
        );

    \I__11484\ : InMux
    port map (
            O => \N__51190\,
            I => \N__51180\
        );

    \I__11483\ : Span4Mux_v
    port map (
            O => \N__51187\,
            I => \N__51177\
        );

    \I__11482\ : InMux
    port map (
            O => \N__51186\,
            I => \N__51174\
        );

    \I__11481\ : Sp12to4
    port map (
            O => \N__51183\,
            I => \N__51171\
        );

    \I__11480\ : LocalMux
    port map (
            O => \N__51180\,
            I => \N__51168\
        );

    \I__11479\ : Span4Mux_h
    port map (
            O => \N__51177\,
            I => \N__51163\
        );

    \I__11478\ : LocalMux
    port map (
            O => \N__51174\,
            I => \N__51163\
        );

    \I__11477\ : Span12Mux_h
    port map (
            O => \N__51171\,
            I => \N__51160\
        );

    \I__11476\ : Span4Mux_v
    port map (
            O => \N__51168\,
            I => \N__51157\
        );

    \I__11475\ : Span4Mux_h
    port map (
            O => \N__51163\,
            I => \N__51154\
        );

    \I__11474\ : Span12Mux_v
    port map (
            O => \N__51160\,
            I => \N__51151\
        );

    \I__11473\ : Span4Mux_h
    port map (
            O => \N__51157\,
            I => \N__51148\
        );

    \I__11472\ : Span4Mux_v
    port map (
            O => \N__51154\,
            I => \N__51145\
        );

    \I__11471\ : Span12Mux_v
    port map (
            O => \N__51151\,
            I => \N__51142\
        );

    \I__11470\ : Sp12to4
    port map (
            O => \N__51148\,
            I => \N__51139\
        );

    \I__11469\ : IoSpan4Mux
    port map (
            O => \N__51145\,
            I => \N__51136\
        );

    \I__11468\ : Odrv12
    port map (
            O => \N__51142\,
            I => scl_c
        );

    \I__11467\ : Odrv12
    port map (
            O => \N__51139\,
            I => scl_c
        );

    \I__11466\ : Odrv4
    port map (
            O => \N__51136\,
            I => scl_c
        );

    \I__11465\ : InMux
    port map (
            O => \N__51129\,
            I => \N__51126\
        );

    \I__11464\ : LocalMux
    port map (
            O => \N__51126\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_0\
        );

    \I__11463\ : InMux
    port map (
            O => \N__51123\,
            I => \N__51113\
        );

    \I__11462\ : InMux
    port map (
            O => \N__51122\,
            I => \N__51113\
        );

    \I__11461\ : InMux
    port map (
            O => \N__51121\,
            I => \N__51104\
        );

    \I__11460\ : InMux
    port map (
            O => \N__51120\,
            I => \N__51104\
        );

    \I__11459\ : InMux
    port map (
            O => \N__51119\,
            I => \N__51104\
        );

    \I__11458\ : InMux
    port map (
            O => \N__51118\,
            I => \N__51104\
        );

    \I__11457\ : LocalMux
    port map (
            O => \N__51113\,
            I => \N__51101\
        );

    \I__11456\ : LocalMux
    port map (
            O => \N__51104\,
            I => \N__51098\
        );

    \I__11455\ : Span4Mux_v
    port map (
            O => \N__51101\,
            I => \N__51095\
        );

    \I__11454\ : Span4Mux_v
    port map (
            O => \N__51098\,
            I => \N__51092\
        );

    \I__11453\ : Span4Mux_h
    port map (
            O => \N__51095\,
            I => \N__51089\
        );

    \I__11452\ : Span4Mux_h
    port map (
            O => \N__51092\,
            I => \N__51086\
        );

    \I__11451\ : Odrv4
    port map (
            O => \N__51089\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0\
        );

    \I__11450\ : Odrv4
    port map (
            O => \N__51086\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0\
        );

    \I__11449\ : InMux
    port map (
            O => \N__51081\,
            I => \N__51070\
        );

    \I__11448\ : InMux
    port map (
            O => \N__51080\,
            I => \N__51070\
        );

    \I__11447\ : InMux
    port map (
            O => \N__51079\,
            I => \N__51059\
        );

    \I__11446\ : InMux
    port map (
            O => \N__51078\,
            I => \N__51059\
        );

    \I__11445\ : InMux
    port map (
            O => \N__51077\,
            I => \N__51059\
        );

    \I__11444\ : InMux
    port map (
            O => \N__51076\,
            I => \N__51059\
        );

    \I__11443\ : InMux
    port map (
            O => \N__51075\,
            I => \N__51059\
        );

    \I__11442\ : LocalMux
    port map (
            O => \N__51070\,
            I => \I2C_top_level_inst1.s_command_1\
        );

    \I__11441\ : LocalMux
    port map (
            O => \N__51059\,
            I => \I2C_top_level_inst1.s_command_1\
        );

    \I__11440\ : CascadeMux
    port map (
            O => \N__51054\,
            I => \N__51049\
        );

    \I__11439\ : CascadeMux
    port map (
            O => \N__51053\,
            I => \N__51045\
        );

    \I__11438\ : InMux
    port map (
            O => \N__51052\,
            I => \N__51037\
        );

    \I__11437\ : InMux
    port map (
            O => \N__51049\,
            I => \N__51037\
        );

    \I__11436\ : InMux
    port map (
            O => \N__51048\,
            I => \N__51037\
        );

    \I__11435\ : InMux
    port map (
            O => \N__51045\,
            I => \N__51032\
        );

    \I__11434\ : InMux
    port map (
            O => \N__51044\,
            I => \N__51032\
        );

    \I__11433\ : LocalMux
    port map (
            O => \N__51037\,
            I => \N__51029\
        );

    \I__11432\ : LocalMux
    port map (
            O => \N__51032\,
            I => \I2C_top_level_inst1.s_command_2\
        );

    \I__11431\ : Odrv4
    port map (
            O => \N__51029\,
            I => \I2C_top_level_inst1.s_command_2\
        );

    \I__11430\ : CascadeMux
    port map (
            O => \N__51024\,
            I => \N__51019\
        );

    \I__11429\ : CascadeMux
    port map (
            O => \N__51023\,
            I => \N__51016\
        );

    \I__11428\ : InMux
    port map (
            O => \N__51022\,
            I => \N__51008\
        );

    \I__11427\ : InMux
    port map (
            O => \N__51019\,
            I => \N__51008\
        );

    \I__11426\ : InMux
    port map (
            O => \N__51016\,
            I => \N__50999\
        );

    \I__11425\ : InMux
    port map (
            O => \N__51015\,
            I => \N__50999\
        );

    \I__11424\ : InMux
    port map (
            O => \N__51014\,
            I => \N__50999\
        );

    \I__11423\ : InMux
    port map (
            O => \N__51013\,
            I => \N__50999\
        );

    \I__11422\ : LocalMux
    port map (
            O => \N__51008\,
            I => \I2C_top_level_inst1.s_command_3\
        );

    \I__11421\ : LocalMux
    port map (
            O => \N__50999\,
            I => \I2C_top_level_inst1.s_command_3\
        );

    \I__11420\ : InMux
    port map (
            O => \N__50994\,
            I => \N__50990\
        );

    \I__11419\ : InMux
    port map (
            O => \N__50993\,
            I => \N__50987\
        );

    \I__11418\ : LocalMux
    port map (
            O => \N__50990\,
            I => \N__50984\
        );

    \I__11417\ : LocalMux
    port map (
            O => \N__50987\,
            I => \N__50980\
        );

    \I__11416\ : Span4Mux_h
    port map (
            O => \N__50984\,
            I => \N__50976\
        );

    \I__11415\ : InMux
    port map (
            O => \N__50983\,
            I => \N__50973\
        );

    \I__11414\ : Span4Mux_h
    port map (
            O => \N__50980\,
            I => \N__50970\
        );

    \I__11413\ : InMux
    port map (
            O => \N__50979\,
            I => \N__50967\
        );

    \I__11412\ : Span4Mux_v
    port map (
            O => \N__50976\,
            I => \N__50960\
        );

    \I__11411\ : LocalMux
    port map (
            O => \N__50973\,
            I => \N__50960\
        );

    \I__11410\ : Span4Mux_v
    port map (
            O => \N__50970\,
            I => \N__50960\
        );

    \I__11409\ : LocalMux
    port map (
            O => \N__50967\,
            I => \I2C_top_level_inst1.s_load_wdata\
        );

    \I__11408\ : Odrv4
    port map (
            O => \N__50960\,
            I => \I2C_top_level_inst1.s_load_wdata\
        );

    \I__11407\ : InMux
    port map (
            O => \N__50955\,
            I => \N__50952\
        );

    \I__11406\ : LocalMux
    port map (
            O => \N__50952\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_0\
        );

    \I__11405\ : InMux
    port map (
            O => \N__50949\,
            I => \N__50946\
        );

    \I__11404\ : LocalMux
    port map (
            O => \N__50946\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_1\
        );

    \I__11403\ : InMux
    port map (
            O => \N__50943\,
            I => \N__50940\
        );

    \I__11402\ : LocalMux
    port map (
            O => \N__50940\,
            I => \N__50937\
        );

    \I__11401\ : Span4Mux_v
    port map (
            O => \N__50937\,
            I => \N__50934\
        );

    \I__11400\ : Span4Mux_v
    port map (
            O => \N__50934\,
            I => \N__50927\
        );

    \I__11399\ : InMux
    port map (
            O => \N__50933\,
            I => \N__50924\
        );

    \I__11398\ : InMux
    port map (
            O => \N__50932\,
            I => \N__50914\
        );

    \I__11397\ : InMux
    port map (
            O => \N__50931\,
            I => \N__50914\
        );

    \I__11396\ : InMux
    port map (
            O => \N__50930\,
            I => \N__50914\
        );

    \I__11395\ : Span4Mux_h
    port map (
            O => \N__50927\,
            I => \N__50909\
        );

    \I__11394\ : LocalMux
    port map (
            O => \N__50924\,
            I => \N__50909\
        );

    \I__11393\ : InMux
    port map (
            O => \N__50923\,
            I => \N__50902\
        );

    \I__11392\ : InMux
    port map (
            O => \N__50922\,
            I => \N__50902\
        );

    \I__11391\ : InMux
    port map (
            O => \N__50921\,
            I => \N__50902\
        );

    \I__11390\ : LocalMux
    port map (
            O => \N__50914\,
            I => \N__50899\
        );

    \I__11389\ : Span4Mux_h
    port map (
            O => \N__50909\,
            I => \N__50896\
        );

    \I__11388\ : LocalMux
    port map (
            O => \N__50902\,
            I => \N__50893\
        );

    \I__11387\ : Odrv4
    port map (
            O => \N__50899\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2\
        );

    \I__11386\ : Odrv4
    port map (
            O => \N__50896\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2\
        );

    \I__11385\ : Odrv4
    port map (
            O => \N__50893\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2\
        );

    \I__11384\ : InMux
    port map (
            O => \N__50886\,
            I => \N__50878\
        );

    \I__11383\ : CascadeMux
    port map (
            O => \N__50885\,
            I => \N__50875\
        );

    \I__11382\ : InMux
    port map (
            O => \N__50884\,
            I => \N__50866\
        );

    \I__11381\ : InMux
    port map (
            O => \N__50883\,
            I => \N__50866\
        );

    \I__11380\ : InMux
    port map (
            O => \N__50882\,
            I => \N__50861\
        );

    \I__11379\ : InMux
    port map (
            O => \N__50881\,
            I => \N__50858\
        );

    \I__11378\ : LocalMux
    port map (
            O => \N__50878\,
            I => \N__50855\
        );

    \I__11377\ : InMux
    port map (
            O => \N__50875\,
            I => \N__50844\
        );

    \I__11376\ : InMux
    port map (
            O => \N__50874\,
            I => \N__50844\
        );

    \I__11375\ : InMux
    port map (
            O => \N__50873\,
            I => \N__50844\
        );

    \I__11374\ : InMux
    port map (
            O => \N__50872\,
            I => \N__50844\
        );

    \I__11373\ : InMux
    port map (
            O => \N__50871\,
            I => \N__50844\
        );

    \I__11372\ : LocalMux
    port map (
            O => \N__50866\,
            I => \N__50841\
        );

    \I__11371\ : InMux
    port map (
            O => \N__50865\,
            I => \N__50836\
        );

    \I__11370\ : InMux
    port map (
            O => \N__50864\,
            I => \N__50836\
        );

    \I__11369\ : LocalMux
    port map (
            O => \N__50861\,
            I => \N__50833\
        );

    \I__11368\ : LocalMux
    port map (
            O => \N__50858\,
            I => \N__50830\
        );

    \I__11367\ : Span4Mux_h
    port map (
            O => \N__50855\,
            I => \N__50821\
        );

    \I__11366\ : LocalMux
    port map (
            O => \N__50844\,
            I => \N__50821\
        );

    \I__11365\ : Span4Mux_v
    port map (
            O => \N__50841\,
            I => \N__50821\
        );

    \I__11364\ : LocalMux
    port map (
            O => \N__50836\,
            I => \N__50821\
        );

    \I__11363\ : Span4Mux_v
    port map (
            O => \N__50833\,
            I => \N__50817\
        );

    \I__11362\ : Span4Mux_h
    port map (
            O => \N__50830\,
            I => \N__50814\
        );

    \I__11361\ : Span4Mux_h
    port map (
            O => \N__50821\,
            I => \N__50811\
        );

    \I__11360\ : InMux
    port map (
            O => \N__50820\,
            I => \N__50808\
        );

    \I__11359\ : Sp12to4
    port map (
            O => \N__50817\,
            I => \N__50805\
        );

    \I__11358\ : Span4Mux_v
    port map (
            O => \N__50814\,
            I => \N__50802\
        );

    \I__11357\ : Span4Mux_v
    port map (
            O => \N__50811\,
            I => \N__50797\
        );

    \I__11356\ : LocalMux
    port map (
            O => \N__50808\,
            I => \N__50797\
        );

    \I__11355\ : Odrv12
    port map (
            O => \N__50805\,
            I => \I2C_top_level_inst1.s_start\
        );

    \I__11354\ : Odrv4
    port map (
            O => \N__50802\,
            I => \I2C_top_level_inst1.s_start\
        );

    \I__11353\ : Odrv4
    port map (
            O => \N__50797\,
            I => \I2C_top_level_inst1.s_start\
        );

    \I__11352\ : InMux
    port map (
            O => \N__50790\,
            I => \N__50787\
        );

    \I__11351\ : LocalMux
    port map (
            O => \N__50787\,
            I => \N__50784\
        );

    \I__11350\ : Span4Mux_h
    port map (
            O => \N__50784\,
            I => \N__50781\
        );

    \I__11349\ : Span4Mux_h
    port map (
            O => \N__50781\,
            I => \N__50778\
        );

    \I__11348\ : Odrv4
    port map (
            O => \N__50778\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_0\
        );

    \I__11347\ : CascadeMux
    port map (
            O => \N__50775\,
            I => \N__50772\
        );

    \I__11346\ : InMux
    port map (
            O => \N__50772\,
            I => \N__50769\
        );

    \I__11345\ : LocalMux
    port map (
            O => \N__50769\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_86_0\
        );

    \I__11344\ : InMux
    port map (
            O => \N__50766\,
            I => \N__50763\
        );

    \I__11343\ : LocalMux
    port map (
            O => \N__50763\,
            I => \N__50760\
        );

    \I__11342\ : Odrv4
    port map (
            O => \N__50760\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_95_0\
        );

    \I__11341\ : InMux
    port map (
            O => \N__50757\,
            I => \N__50754\
        );

    \I__11340\ : LocalMux
    port map (
            O => \N__50754\,
            I => \N__50751\
        );

    \I__11339\ : Span4Mux_h
    port map (
            O => \N__50751\,
            I => \N__50748\
        );

    \I__11338\ : Span4Mux_h
    port map (
            O => \N__50748\,
            I => \N__50743\
        );

    \I__11337\ : InMux
    port map (
            O => \N__50747\,
            I => \N__50738\
        );

    \I__11336\ : InMux
    port map (
            O => \N__50746\,
            I => \N__50738\
        );

    \I__11335\ : Span4Mux_h
    port map (
            O => \N__50743\,
            I => \N__50735\
        );

    \I__11334\ : LocalMux
    port map (
            O => \N__50738\,
            I => \N__50732\
        );

    \I__11333\ : Odrv4
    port map (
            O => \N__50735\,
            I => \I2C_top_level_inst1.s_stop\
        );

    \I__11332\ : Odrv4
    port map (
            O => \N__50732\,
            I => \I2C_top_level_inst1.s_stop\
        );

    \I__11331\ : InMux
    port map (
            O => \N__50727\,
            I => \N__50724\
        );

    \I__11330\ : LocalMux
    port map (
            O => \N__50724\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_0\
        );

    \I__11329\ : InMux
    port map (
            O => \N__50721\,
            I => \N__50718\
        );

    \I__11328\ : LocalMux
    port map (
            O => \N__50718\,
            I => \N__50711\
        );

    \I__11327\ : InMux
    port map (
            O => \N__50717\,
            I => \N__50706\
        );

    \I__11326\ : InMux
    port map (
            O => \N__50716\,
            I => \N__50706\
        );

    \I__11325\ : InMux
    port map (
            O => \N__50715\,
            I => \N__50701\
        );

    \I__11324\ : InMux
    port map (
            O => \N__50714\,
            I => \N__50701\
        );

    \I__11323\ : Span4Mux_v
    port map (
            O => \N__50711\,
            I => \N__50698\
        );

    \I__11322\ : LocalMux
    port map (
            O => \N__50706\,
            I => \N__50693\
        );

    \I__11321\ : LocalMux
    port map (
            O => \N__50701\,
            I => \N__50693\
        );

    \I__11320\ : Span4Mux_h
    port map (
            O => \N__50698\,
            I => \N__50690\
        );

    \I__11319\ : Span12Mux_v
    port map (
            O => \N__50693\,
            I => \N__50687\
        );

    \I__11318\ : Odrv4
    port map (
            O => \N__50690\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2\
        );

    \I__11317\ : Odrv12
    port map (
            O => \N__50687\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2\
        );

    \I__11316\ : InMux
    port map (
            O => \N__50682\,
            I => \N__50678\
        );

    \I__11315\ : InMux
    port map (
            O => \N__50681\,
            I => \N__50675\
        );

    \I__11314\ : LocalMux
    port map (
            O => \N__50678\,
            I => \N__50670\
        );

    \I__11313\ : LocalMux
    port map (
            O => \N__50675\,
            I => \N__50670\
        );

    \I__11312\ : Odrv4
    port map (
            O => \N__50670\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_844_2\
        );

    \I__11311\ : InMux
    port map (
            O => \N__50667\,
            I => \N__50663\
        );

    \I__11310\ : InMux
    port map (
            O => \N__50666\,
            I => \N__50660\
        );

    \I__11309\ : LocalMux
    port map (
            O => \N__50663\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2\
        );

    \I__11308\ : LocalMux
    port map (
            O => \N__50660\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2\
        );

    \I__11307\ : InMux
    port map (
            O => \N__50655\,
            I => \N__50652\
        );

    \I__11306\ : LocalMux
    port map (
            O => \N__50652\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_1\
        );

    \I__11305\ : InMux
    port map (
            O => \N__50649\,
            I => \N__50646\
        );

    \I__11304\ : LocalMux
    port map (
            O => \N__50646\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_1\
        );

    \I__11303\ : InMux
    port map (
            O => \N__50643\,
            I => \N__50637\
        );

    \I__11302\ : InMux
    port map (
            O => \N__50642\,
            I => \N__50637\
        );

    \I__11301\ : LocalMux
    port map (
            O => \N__50637\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1754_1\
        );

    \I__11300\ : CascadeMux
    port map (
            O => \N__50634\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0_cascade_\
        );

    \I__11299\ : InMux
    port map (
            O => \N__50631\,
            I => \N__50628\
        );

    \I__11298\ : LocalMux
    port map (
            O => \N__50628\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_25\
        );

    \I__11297\ : CascadeMux
    port map (
            O => \N__50625\,
            I => \N__50622\
        );

    \I__11296\ : InMux
    port map (
            O => \N__50622\,
            I => \N__50618\
        );

    \I__11295\ : InMux
    port map (
            O => \N__50621\,
            I => \N__50615\
        );

    \I__11294\ : LocalMux
    port map (
            O => \N__50618\,
            I => \N__50612\
        );

    \I__11293\ : LocalMux
    port map (
            O => \N__50615\,
            I => \N__50608\
        );

    \I__11292\ : Span4Mux_h
    port map (
            O => \N__50612\,
            I => \N__50605\
        );

    \I__11291\ : InMux
    port map (
            O => \N__50611\,
            I => \N__50602\
        );

    \I__11290\ : Span4Mux_v
    port map (
            O => \N__50608\,
            I => \N__50597\
        );

    \I__11289\ : Span4Mux_h
    port map (
            O => \N__50605\,
            I => \N__50597\
        );

    \I__11288\ : LocalMux
    port map (
            O => \N__50602\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2\
        );

    \I__11287\ : Odrv4
    port map (
            O => \N__50597\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2\
        );

    \I__11286\ : InMux
    port map (
            O => \N__50592\,
            I => \N__50589\
        );

    \I__11285\ : LocalMux
    port map (
            O => \N__50589\,
            I => \N__50586\
        );

    \I__11284\ : Span4Mux_h
    port map (
            O => \N__50586\,
            I => \N__50582\
        );

    \I__11283\ : InMux
    port map (
            O => \N__50585\,
            I => \N__50578\
        );

    \I__11282\ : Span4Mux_v
    port map (
            O => \N__50582\,
            I => \N__50575\
        );

    \I__11281\ : InMux
    port map (
            O => \N__50581\,
            I => \N__50572\
        );

    \I__11280\ : LocalMux
    port map (
            O => \N__50578\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i\
        );

    \I__11279\ : Odrv4
    port map (
            O => \N__50575\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i\
        );

    \I__11278\ : LocalMux
    port map (
            O => \N__50572\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i\
        );

    \I__11277\ : CascadeMux
    port map (
            O => \N__50565\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_24_cascade_\
        );

    \I__11276\ : CascadeMux
    port map (
            O => \N__50562\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_11_cascade_\
        );

    \I__11275\ : InMux
    port map (
            O => \N__50559\,
            I => \N__50555\
        );

    \I__11274\ : InMux
    port map (
            O => \N__50558\,
            I => \N__50552\
        );

    \I__11273\ : LocalMux
    port map (
            O => \N__50555\,
            I => \N__50546\
        );

    \I__11272\ : LocalMux
    port map (
            O => \N__50552\,
            I => \N__50546\
        );

    \I__11271\ : InMux
    port map (
            O => \N__50551\,
            I => \N__50540\
        );

    \I__11270\ : Span4Mux_v
    port map (
            O => \N__50546\,
            I => \N__50533\
        );

    \I__11269\ : InMux
    port map (
            O => \N__50545\,
            I => \N__50530\
        );

    \I__11268\ : InMux
    port map (
            O => \N__50544\,
            I => \N__50525\
        );

    \I__11267\ : InMux
    port map (
            O => \N__50543\,
            I => \N__50525\
        );

    \I__11266\ : LocalMux
    port map (
            O => \N__50540\,
            I => \N__50522\
        );

    \I__11265\ : InMux
    port map (
            O => \N__50539\,
            I => \N__50517\
        );

    \I__11264\ : InMux
    port map (
            O => \N__50538\,
            I => \N__50517\
        );

    \I__11263\ : InMux
    port map (
            O => \N__50537\,
            I => \N__50512\
        );

    \I__11262\ : InMux
    port map (
            O => \N__50536\,
            I => \N__50512\
        );

    \I__11261\ : Span4Mux_h
    port map (
            O => \N__50533\,
            I => \N__50509\
        );

    \I__11260\ : LocalMux
    port map (
            O => \N__50530\,
            I => \N__50506\
        );

    \I__11259\ : LocalMux
    port map (
            O => \N__50525\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\
        );

    \I__11258\ : Odrv4
    port map (
            O => \N__50522\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\
        );

    \I__11257\ : LocalMux
    port map (
            O => \N__50517\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\
        );

    \I__11256\ : LocalMux
    port map (
            O => \N__50512\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\
        );

    \I__11255\ : Odrv4
    port map (
            O => \N__50509\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\
        );

    \I__11254\ : Odrv12
    port map (
            O => \N__50506\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\
        );

    \I__11253\ : CascadeMux
    port map (
            O => \N__50493\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_11_cascade_\
        );

    \I__11252\ : CascadeMux
    port map (
            O => \N__50490\,
            I => \N__50487\
        );

    \I__11251\ : InMux
    port map (
            O => \N__50487\,
            I => \N__50484\
        );

    \I__11250\ : LocalMux
    port map (
            O => \N__50484\,
            I => \N__50481\
        );

    \I__11249\ : Span4Mux_v
    port map (
            O => \N__50481\,
            I => \N__50478\
        );

    \I__11248\ : Span4Mux_h
    port map (
            O => \N__50478\,
            I => \N__50475\
        );

    \I__11247\ : Span4Mux_h
    port map (
            O => \N__50475\,
            I => \N__50472\
        );

    \I__11246\ : Odrv4
    port map (
            O => \N__50472\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_2_11\
        );

    \I__11245\ : CascadeMux
    port map (
            O => \N__50469\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_1_2_0_cascade_\
        );

    \I__11244\ : CascadeMux
    port map (
            O => \N__50466\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i_cascade_\
        );

    \I__11243\ : CascadeMux
    port map (
            O => \N__50463\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_372_cascade_\
        );

    \I__11242\ : InMux
    port map (
            O => \N__50460\,
            I => \N__50457\
        );

    \I__11241\ : LocalMux
    port map (
            O => \N__50457\,
            I => \N__50453\
        );

    \I__11240\ : InMux
    port map (
            O => \N__50456\,
            I => \N__50450\
        );

    \I__11239\ : Span4Mux_h
    port map (
            O => \N__50453\,
            I => \N__50446\
        );

    \I__11238\ : LocalMux
    port map (
            O => \N__50450\,
            I => \N__50443\
        );

    \I__11237\ : InMux
    port map (
            O => \N__50449\,
            I => \N__50440\
        );

    \I__11236\ : Span4Mux_h
    port map (
            O => \N__50446\,
            I => \N__50437\
        );

    \I__11235\ : Span12Mux_h
    port map (
            O => \N__50443\,
            I => \N__50434\
        );

    \I__11234\ : LocalMux
    port map (
            O => \N__50440\,
            I => \N_409\
        );

    \I__11233\ : Odrv4
    port map (
            O => \N__50437\,
            I => \N_409\
        );

    \I__11232\ : Odrv12
    port map (
            O => \N__50434\,
            I => \N_409\
        );

    \I__11231\ : InMux
    port map (
            O => \N__50427\,
            I => \N__50424\
        );

    \I__11230\ : LocalMux
    port map (
            O => \N__50424\,
            I => \N__50421\
        );

    \I__11229\ : Odrv4
    port map (
            O => \N__50421\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_a3_1_0_14\
        );

    \I__11228\ : CascadeMux
    port map (
            O => \N__50418\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_412_0_cascade_\
        );

    \I__11227\ : InMux
    port map (
            O => \N__50415\,
            I => \N__50412\
        );

    \I__11226\ : LocalMux
    port map (
            O => \N__50412\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_1_14\
        );

    \I__11225\ : CascadeMux
    port map (
            O => \N__50409\,
            I => \N__50398\
        );

    \I__11224\ : InMux
    port map (
            O => \N__50408\,
            I => \N__50381\
        );

    \I__11223\ : InMux
    port map (
            O => \N__50407\,
            I => \N__50381\
        );

    \I__11222\ : InMux
    port map (
            O => \N__50406\,
            I => \N__50368\
        );

    \I__11221\ : InMux
    port map (
            O => \N__50405\,
            I => \N__50368\
        );

    \I__11220\ : InMux
    port map (
            O => \N__50404\,
            I => \N__50368\
        );

    \I__11219\ : InMux
    port map (
            O => \N__50403\,
            I => \N__50368\
        );

    \I__11218\ : InMux
    port map (
            O => \N__50402\,
            I => \N__50368\
        );

    \I__11217\ : InMux
    port map (
            O => \N__50401\,
            I => \N__50359\
        );

    \I__11216\ : InMux
    port map (
            O => \N__50398\,
            I => \N__50359\
        );

    \I__11215\ : InMux
    port map (
            O => \N__50397\,
            I => \N__50359\
        );

    \I__11214\ : InMux
    port map (
            O => \N__50396\,
            I => \N__50359\
        );

    \I__11213\ : CascadeMux
    port map (
            O => \N__50395\,
            I => \N__50356\
        );

    \I__11212\ : InMux
    port map (
            O => \N__50394\,
            I => \N__50334\
        );

    \I__11211\ : InMux
    port map (
            O => \N__50393\,
            I => \N__50334\
        );

    \I__11210\ : InMux
    port map (
            O => \N__50392\,
            I => \N__50334\
        );

    \I__11209\ : InMux
    port map (
            O => \N__50391\,
            I => \N__50334\
        );

    \I__11208\ : InMux
    port map (
            O => \N__50390\,
            I => \N__50334\
        );

    \I__11207\ : InMux
    port map (
            O => \N__50389\,
            I => \N__50334\
        );

    \I__11206\ : InMux
    port map (
            O => \N__50388\,
            I => \N__50329\
        );

    \I__11205\ : InMux
    port map (
            O => \N__50387\,
            I => \N__50329\
        );

    \I__11204\ : CascadeMux
    port map (
            O => \N__50386\,
            I => \N__50326\
        );

    \I__11203\ : LocalMux
    port map (
            O => \N__50381\,
            I => \N__50323\
        );

    \I__11202\ : InMux
    port map (
            O => \N__50380\,
            I => \N__50318\
        );

    \I__11201\ : InMux
    port map (
            O => \N__50379\,
            I => \N__50318\
        );

    \I__11200\ : LocalMux
    port map (
            O => \N__50368\,
            I => \N__50313\
        );

    \I__11199\ : LocalMux
    port map (
            O => \N__50359\,
            I => \N__50313\
        );

    \I__11198\ : InMux
    port map (
            O => \N__50356\,
            I => \N__50308\
        );

    \I__11197\ : InMux
    port map (
            O => \N__50355\,
            I => \N__50308\
        );

    \I__11196\ : InMux
    port map (
            O => \N__50354\,
            I => \N__50301\
        );

    \I__11195\ : InMux
    port map (
            O => \N__50353\,
            I => \N__50301\
        );

    \I__11194\ : InMux
    port map (
            O => \N__50352\,
            I => \N__50301\
        );

    \I__11193\ : InMux
    port map (
            O => \N__50351\,
            I => \N__50290\
        );

    \I__11192\ : InMux
    port map (
            O => \N__50350\,
            I => \N__50290\
        );

    \I__11191\ : InMux
    port map (
            O => \N__50349\,
            I => \N__50290\
        );

    \I__11190\ : InMux
    port map (
            O => \N__50348\,
            I => \N__50290\
        );

    \I__11189\ : InMux
    port map (
            O => \N__50347\,
            I => \N__50290\
        );

    \I__11188\ : LocalMux
    port map (
            O => \N__50334\,
            I => \N__50285\
        );

    \I__11187\ : LocalMux
    port map (
            O => \N__50329\,
            I => \N__50285\
        );

    \I__11186\ : InMux
    port map (
            O => \N__50326\,
            I => \N__50282\
        );

    \I__11185\ : Span4Mux_v
    port map (
            O => \N__50323\,
            I => \N__50277\
        );

    \I__11184\ : LocalMux
    port map (
            O => \N__50318\,
            I => \N__50277\
        );

    \I__11183\ : Span4Mux_h
    port map (
            O => \N__50313\,
            I => \N__50274\
        );

    \I__11182\ : LocalMux
    port map (
            O => \N__50308\,
            I => \N__50265\
        );

    \I__11181\ : LocalMux
    port map (
            O => \N__50301\,
            I => \N__50265\
        );

    \I__11180\ : LocalMux
    port map (
            O => \N__50290\,
            I => \N__50265\
        );

    \I__11179\ : Span4Mux_v
    port map (
            O => \N__50285\,
            I => \N__50265\
        );

    \I__11178\ : LocalMux
    port map (
            O => \N__50282\,
            I => \N__50262\
        );

    \I__11177\ : Span4Mux_h
    port map (
            O => \N__50277\,
            I => \N__50257\
        );

    \I__11176\ : Span4Mux_v
    port map (
            O => \N__50274\,
            I => \N__50257\
        );

    \I__11175\ : Span4Mux_h
    port map (
            O => \N__50265\,
            I => \N__50254\
        );

    \I__11174\ : Span4Mux_h
    port map (
            O => \N__50262\,
            I => \N__50251\
        );

    \I__11173\ : Span4Mux_v
    port map (
            O => \N__50257\,
            I => \N__50248\
        );

    \I__11172\ : Span4Mux_v
    port map (
            O => \N__50254\,
            I => \N__50245\
        );

    \I__11171\ : Span4Mux_h
    port map (
            O => \N__50251\,
            I => \N__50239\
        );

    \I__11170\ : Span4Mux_h
    port map (
            O => \N__50248\,
            I => \N__50239\
        );

    \I__11169\ : Span4Mux_h
    port map (
            O => \N__50245\,
            I => \N__50236\
        );

    \I__11168\ : InMux
    port map (
            O => \N__50244\,
            I => \N__50233\
        );

    \I__11167\ : Odrv4
    port map (
            O => \N__50239\,
            I => \N_410\
        );

    \I__11166\ : Odrv4
    port map (
            O => \N__50236\,
            I => \N_410\
        );

    \I__11165\ : LocalMux
    port map (
            O => \N__50233\,
            I => \N_410\
        );

    \I__11164\ : InMux
    port map (
            O => \N__50226\,
            I => \N__50223\
        );

    \I__11163\ : LocalMux
    port map (
            O => \N__50223\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_1_0_14\
        );

    \I__11162\ : CascadeMux
    port map (
            O => \N__50220\,
            I => \N__50215\
        );

    \I__11161\ : InMux
    port map (
            O => \N__50219\,
            I => \N__50208\
        );

    \I__11160\ : InMux
    port map (
            O => \N__50218\,
            I => \N__50208\
        );

    \I__11159\ : InMux
    port map (
            O => \N__50215\,
            I => \N__50208\
        );

    \I__11158\ : LocalMux
    port map (
            O => \N__50208\,
            I => \N__50205\
        );

    \I__11157\ : Span4Mux_v
    port map (
            O => \N__50205\,
            I => \N__50202\
        );

    \I__11156\ : Span4Mux_h
    port map (
            O => \N__50202\,
            I => \N__50199\
        );

    \I__11155\ : Odrv4
    port map (
            O => \N__50199\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_322\
        );

    \I__11154\ : CascadeMux
    port map (
            O => \N__50196\,
            I => \N__50193\
        );

    \I__11153\ : InMux
    port map (
            O => \N__50193\,
            I => \N__50188\
        );

    \I__11152\ : InMux
    port map (
            O => \N__50192\,
            I => \N__50185\
        );

    \I__11151\ : InMux
    port map (
            O => \N__50191\,
            I => \N__50182\
        );

    \I__11150\ : LocalMux
    port map (
            O => \N__50188\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0\
        );

    \I__11149\ : LocalMux
    port map (
            O => \N__50185\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0\
        );

    \I__11148\ : LocalMux
    port map (
            O => \N__50182\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0\
        );

    \I__11147\ : InMux
    port map (
            O => \N__50175\,
            I => \N__50172\
        );

    \I__11146\ : LocalMux
    port map (
            O => \N__50172\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0\
        );

    \I__11145\ : CascadeMux
    port map (
            O => \N__50169\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0_cascade_\
        );

    \I__11144\ : InMux
    port map (
            O => \N__50166\,
            I => \N__50163\
        );

    \I__11143\ : LocalMux
    port map (
            O => \N__50163\,
            I => \N__50160\
        );

    \I__11142\ : Span4Mux_v
    port map (
            O => \N__50160\,
            I => \N__50157\
        );

    \I__11141\ : Odrv4
    port map (
            O => \N__50157\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_267\
        );

    \I__11140\ : InMux
    port map (
            O => \N__50154\,
            I => \N__50151\
        );

    \I__11139\ : LocalMux
    port map (
            O => \N__50151\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_394\
        );

    \I__11138\ : CascadeMux
    port map (
            O => \N__50148\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_267_cascade_\
        );

    \I__11137\ : InMux
    port map (
            O => \N__50145\,
            I => \N__50142\
        );

    \I__11136\ : LocalMux
    port map (
            O => \N__50142\,
            I => \N__50134\
        );

    \I__11135\ : InMux
    port map (
            O => \N__50141\,
            I => \N__50131\
        );

    \I__11134\ : InMux
    port map (
            O => \N__50140\,
            I => \N__50126\
        );

    \I__11133\ : InMux
    port map (
            O => \N__50139\,
            I => \N__50126\
        );

    \I__11132\ : InMux
    port map (
            O => \N__50138\,
            I => \N__50121\
        );

    \I__11131\ : InMux
    port map (
            O => \N__50137\,
            I => \N__50121\
        );

    \I__11130\ : Span4Mux_h
    port map (
            O => \N__50134\,
            I => \N__50114\
        );

    \I__11129\ : LocalMux
    port map (
            O => \N__50131\,
            I => \N__50114\
        );

    \I__11128\ : LocalMux
    port map (
            O => \N__50126\,
            I => \N__50114\
        );

    \I__11127\ : LocalMux
    port map (
            O => \N__50121\,
            I => \N__50109\
        );

    \I__11126\ : Span4Mux_v
    port map (
            O => \N__50114\,
            I => \N__50106\
        );

    \I__11125\ : InMux
    port map (
            O => \N__50113\,
            I => \N__50103\
        );

    \I__11124\ : InMux
    port map (
            O => \N__50112\,
            I => \N__50100\
        );

    \I__11123\ : Odrv4
    port map (
            O => \N__50109\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0\
        );

    \I__11122\ : Odrv4
    port map (
            O => \N__50106\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0\
        );

    \I__11121\ : LocalMux
    port map (
            O => \N__50103\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0\
        );

    \I__11120\ : LocalMux
    port map (
            O => \N__50100\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0\
        );

    \I__11119\ : CEMux
    port map (
            O => \N__50091\,
            I => \N__50088\
        );

    \I__11118\ : LocalMux
    port map (
            O => \N__50088\,
            I => \N__50084\
        );

    \I__11117\ : CEMux
    port map (
            O => \N__50087\,
            I => \N__50081\
        );

    \I__11116\ : Span4Mux_h
    port map (
            O => \N__50084\,
            I => \N__50077\
        );

    \I__11115\ : LocalMux
    port map (
            O => \N__50081\,
            I => \N__50073\
        );

    \I__11114\ : CEMux
    port map (
            O => \N__50080\,
            I => \N__50070\
        );

    \I__11113\ : Span4Mux_v
    port map (
            O => \N__50077\,
            I => \N__50067\
        );

    \I__11112\ : CEMux
    port map (
            O => \N__50076\,
            I => \N__50064\
        );

    \I__11111\ : Span4Mux_h
    port map (
            O => \N__50073\,
            I => \N__50061\
        );

    \I__11110\ : LocalMux
    port map (
            O => \N__50070\,
            I => \N__50058\
        );

    \I__11109\ : Span4Mux_v
    port map (
            O => \N__50067\,
            I => \N__50053\
        );

    \I__11108\ : LocalMux
    port map (
            O => \N__50064\,
            I => \N__50053\
        );

    \I__11107\ : Span4Mux_h
    port map (
            O => \N__50061\,
            I => \N__50046\
        );

    \I__11106\ : Span4Mux_h
    port map (
            O => \N__50058\,
            I => \N__50043\
        );

    \I__11105\ : Span4Mux_h
    port map (
            O => \N__50053\,
            I => \N__50040\
        );

    \I__11104\ : CEMux
    port map (
            O => \N__50052\,
            I => \N__50037\
        );

    \I__11103\ : InMux
    port map (
            O => \N__50051\,
            I => \N__50030\
        );

    \I__11102\ : InMux
    port map (
            O => \N__50050\,
            I => \N__50030\
        );

    \I__11101\ : InMux
    port map (
            O => \N__50049\,
            I => \N__50030\
        );

    \I__11100\ : Odrv4
    port map (
            O => \N__50046\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\
        );

    \I__11099\ : Odrv4
    port map (
            O => \N__50043\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\
        );

    \I__11098\ : Odrv4
    port map (
            O => \N__50040\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\
        );

    \I__11097\ : LocalMux
    port map (
            O => \N__50037\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\
        );

    \I__11096\ : LocalMux
    port map (
            O => \N__50030\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\
        );

    \I__11095\ : CascadeMux
    port map (
            O => \N__50019\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_1_1_i_m2_1_9_cascade_\
        );

    \I__11094\ : InMux
    port map (
            O => \N__50016\,
            I => \N__50012\
        );

    \I__11093\ : InMux
    port map (
            O => \N__50015\,
            I => \N__50009\
        );

    \I__11092\ : LocalMux
    port map (
            O => \N__50012\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_101\
        );

    \I__11091\ : LocalMux
    port map (
            O => \N__50009\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_101\
        );

    \I__11090\ : InMux
    port map (
            O => \N__50004\,
            I => \N__50001\
        );

    \I__11089\ : LocalMux
    port map (
            O => \N__50001\,
            I => \N__49998\
        );

    \I__11088\ : Span4Mux_v
    port map (
            O => \N__49998\,
            I => \N__49994\
        );

    \I__11087\ : InMux
    port map (
            O => \N__49997\,
            I => \N__49991\
        );

    \I__11086\ : Odrv4
    port map (
            O => \N__49994\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0\
        );

    \I__11085\ : LocalMux
    port map (
            O => \N__49991\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0\
        );

    \I__11084\ : CascadeMux
    port map (
            O => \N__49986\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3_cascade_\
        );

    \I__11083\ : InMux
    port map (
            O => \N__49983\,
            I => \N__49980\
        );

    \I__11082\ : LocalMux
    port map (
            O => \N__49980\,
            I => \N__49977\
        );

    \I__11081\ : Span4Mux_v
    port map (
            O => \N__49977\,
            I => \N__49974\
        );

    \I__11080\ : Span4Mux_h
    port map (
            O => \N__49974\,
            I => \N__49971\
        );

    \I__11079\ : Span4Mux_h
    port map (
            O => \N__49971\,
            I => \N__49968\
        );

    \I__11078\ : Odrv4
    port map (
            O => \N__49968\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_3\
        );

    \I__11077\ : InMux
    port map (
            O => \N__49965\,
            I => \N__49962\
        );

    \I__11076\ : LocalMux
    port map (
            O => \N__49962\,
            I => \N__49958\
        );

    \I__11075\ : InMux
    port map (
            O => \N__49961\,
            I => \N__49955\
        );

    \I__11074\ : Span4Mux_h
    port map (
            O => \N__49958\,
            I => \N__49952\
        );

    \I__11073\ : LocalMux
    port map (
            O => \N__49955\,
            I => \N__49949\
        );

    \I__11072\ : Span4Mux_v
    port map (
            O => \N__49952\,
            I => \N__49943\
        );

    \I__11071\ : Span4Mux_h
    port map (
            O => \N__49949\,
            I => \N__49943\
        );

    \I__11070\ : InMux
    port map (
            O => \N__49948\,
            I => \N__49940\
        );

    \I__11069\ : Odrv4
    port map (
            O => \N__49943\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_2
        );

    \I__11068\ : LocalMux
    port map (
            O => \N__49940\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_2
        );

    \I__11067\ : CascadeMux
    port map (
            O => \N__49935\,
            I => \N__49932\
        );

    \I__11066\ : InMux
    port map (
            O => \N__49932\,
            I => \N__49929\
        );

    \I__11065\ : LocalMux
    port map (
            O => \N__49929\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_2\
        );

    \I__11064\ : InMux
    port map (
            O => \N__49926\,
            I => \N__49923\
        );

    \I__11063\ : LocalMux
    port map (
            O => \N__49923\,
            I => \N__49920\
        );

    \I__11062\ : Odrv4
    port map (
            O => \N__49920\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_2\
        );

    \I__11061\ : CascadeMux
    port map (
            O => \N__49917\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2QZ0Z5_cascade_\
        );

    \I__11060\ : InMux
    port map (
            O => \N__49914\,
            I => \N__49911\
        );

    \I__11059\ : LocalMux
    port map (
            O => \N__49911\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2\
        );

    \I__11058\ : CascadeMux
    port map (
            O => \N__49908\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2_cascade_\
        );

    \I__11057\ : InMux
    port map (
            O => \N__49905\,
            I => \N__49902\
        );

    \I__11056\ : LocalMux
    port map (
            O => \N__49902\,
            I => \N__49899\
        );

    \I__11055\ : Sp12to4
    port map (
            O => \N__49899\,
            I => \N__49896\
        );

    \I__11054\ : Odrv12
    port map (
            O => \N__49896\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_2\
        );

    \I__11053\ : CascadeMux
    port map (
            O => \N__49893\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_6_0_0_cascade_\
        );

    \I__11052\ : InMux
    port map (
            O => \N__49890\,
            I => \N__49887\
        );

    \I__11051\ : LocalMux
    port map (
            O => \N__49887\,
            I => \N__49884\
        );

    \I__11050\ : Span12Mux_v
    port map (
            O => \N__49884\,
            I => \N__49881\
        );

    \I__11049\ : Odrv12
    port map (
            O => \N__49881\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_607\
        );

    \I__11048\ : CascadeMux
    port map (
            O => \N__49878\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_15_cascade_\
        );

    \I__11047\ : InMux
    port map (
            O => \N__49875\,
            I => \N__49872\
        );

    \I__11046\ : LocalMux
    port map (
            O => \N__49872\,
            I => \N__49869\
        );

    \I__11045\ : Span4Mux_h
    port map (
            O => \N__49869\,
            I => \N__49866\
        );

    \I__11044\ : Span4Mux_h
    port map (
            O => \N__49866\,
            I => \N__49863\
        );

    \I__11043\ : Odrv4
    port map (
            O => \N__49863\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_1_15\
        );

    \I__11042\ : CascadeMux
    port map (
            O => \N__49860\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10_cascade_\
        );

    \I__11041\ : InMux
    port map (
            O => \N__49857\,
            I => \N__49854\
        );

    \I__11040\ : LocalMux
    port map (
            O => \N__49854\,
            I => \N__49851\
        );

    \I__11039\ : Span4Mux_v
    port map (
            O => \N__49851\,
            I => \N__49848\
        );

    \I__11038\ : Span4Mux_h
    port map (
            O => \N__49848\,
            I => \N__49845\
        );

    \I__11037\ : Odrv4
    port map (
            O => \N__49845\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_10\
        );

    \I__11036\ : InMux
    port map (
            O => \N__49842\,
            I => \N__49839\
        );

    \I__11035\ : LocalMux
    port map (
            O => \N__49839\,
            I => \N__49836\
        );

    \I__11034\ : Span4Mux_h
    port map (
            O => \N__49836\,
            I => \N__49833\
        );

    \I__11033\ : Span4Mux_v
    port map (
            O => \N__49833\,
            I => \N__49829\
        );

    \I__11032\ : InMux
    port map (
            O => \N__49832\,
            I => \N__49826\
        );

    \I__11031\ : Sp12to4
    port map (
            O => \N__49829\,
            I => \N__49823\
        );

    \I__11030\ : LocalMux
    port map (
            O => \N__49826\,
            I => \N__49820\
        );

    \I__11029\ : Span12Mux_h
    port map (
            O => \N__49823\,
            I => \N__49816\
        );

    \I__11028\ : Span4Mux_v
    port map (
            O => \N__49820\,
            I => \N__49813\
        );

    \I__11027\ : InMux
    port map (
            O => \N__49819\,
            I => \N__49810\
        );

    \I__11026\ : Odrv12
    port map (
            O => \N__49816\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_9
        );

    \I__11025\ : Odrv4
    port map (
            O => \N__49813\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_9
        );

    \I__11024\ : LocalMux
    port map (
            O => \N__49810\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_9
        );

    \I__11023\ : CascadeMux
    port map (
            O => \N__49803\,
            I => \N__49800\
        );

    \I__11022\ : InMux
    port map (
            O => \N__49800\,
            I => \N__49797\
        );

    \I__11021\ : LocalMux
    port map (
            O => \N__49797\,
            I => \N__49794\
        );

    \I__11020\ : Odrv4
    port map (
            O => \N__49794\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_9\
        );

    \I__11019\ : InMux
    port map (
            O => \N__49791\,
            I => \N__49788\
        );

    \I__11018\ : LocalMux
    port map (
            O => \N__49788\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_9\
        );

    \I__11017\ : CascadeMux
    port map (
            O => \N__49785\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044QZ0Z5_cascade_\
        );

    \I__11016\ : InMux
    port map (
            O => \N__49782\,
            I => \N__49779\
        );

    \I__11015\ : LocalMux
    port map (
            O => \N__49779\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9\
        );

    \I__11014\ : InMux
    port map (
            O => \N__49776\,
            I => \N__49773\
        );

    \I__11013\ : LocalMux
    port map (
            O => \N__49773\,
            I => \N__49770\
        );

    \I__11012\ : Span4Mux_v
    port map (
            O => \N__49770\,
            I => \N__49767\
        );

    \I__11011\ : Span4Mux_v
    port map (
            O => \N__49767\,
            I => \N__49764\
        );

    \I__11010\ : Odrv4
    port map (
            O => \N__49764\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_8\
        );

    \I__11009\ : CascadeMux
    port map (
            O => \N__49761\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9_cascade_\
        );

    \I__11008\ : InMux
    port map (
            O => \N__49758\,
            I => \N__49755\
        );

    \I__11007\ : LocalMux
    port map (
            O => \N__49755\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_9\
        );

    \I__11006\ : InMux
    port map (
            O => \N__49752\,
            I => \N__49748\
        );

    \I__11005\ : InMux
    port map (
            O => \N__49751\,
            I => \N__49744\
        );

    \I__11004\ : LocalMux
    port map (
            O => \N__49748\,
            I => \N__49741\
        );

    \I__11003\ : CascadeMux
    port map (
            O => \N__49747\,
            I => \N__49738\
        );

    \I__11002\ : LocalMux
    port map (
            O => \N__49744\,
            I => \N__49735\
        );

    \I__11001\ : Span12Mux_v
    port map (
            O => \N__49741\,
            I => \N__49732\
        );

    \I__11000\ : InMux
    port map (
            O => \N__49738\,
            I => \N__49729\
        );

    \I__10999\ : Span4Mux_v
    port map (
            O => \N__49735\,
            I => \N__49726\
        );

    \I__10998\ : Odrv12
    port map (
            O => \N__49732\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_2
        );

    \I__10997\ : LocalMux
    port map (
            O => \N__49729\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_2
        );

    \I__10996\ : Odrv4
    port map (
            O => \N__49726\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_2
        );

    \I__10995\ : InMux
    port map (
            O => \N__49719\,
            I => \N__49715\
        );

    \I__10994\ : CascadeMux
    port map (
            O => \N__49718\,
            I => \N__49712\
        );

    \I__10993\ : LocalMux
    port map (
            O => \N__49715\,
            I => \N__49709\
        );

    \I__10992\ : InMux
    port map (
            O => \N__49712\,
            I => \N__49706\
        );

    \I__10991\ : Span4Mux_v
    port map (
            O => \N__49709\,
            I => \N__49703\
        );

    \I__10990\ : LocalMux
    port map (
            O => \N__49706\,
            I => \N__49700\
        );

    \I__10989\ : Sp12to4
    port map (
            O => \N__49703\,
            I => \N__49697\
        );

    \I__10988\ : Span4Mux_h
    port map (
            O => \N__49700\,
            I => \N__49694\
        );

    \I__10987\ : Span12Mux_h
    port map (
            O => \N__49697\,
            I => \N__49690\
        );

    \I__10986\ : Span4Mux_v
    port map (
            O => \N__49694\,
            I => \N__49687\
        );

    \I__10985\ : InMux
    port map (
            O => \N__49693\,
            I => \N__49684\
        );

    \I__10984\ : Odrv12
    port map (
            O => \N__49690\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_3
        );

    \I__10983\ : Odrv4
    port map (
            O => \N__49687\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_3
        );

    \I__10982\ : LocalMux
    port map (
            O => \N__49684\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_3
        );

    \I__10981\ : InMux
    port map (
            O => \N__49677\,
            I => \N__49673\
        );

    \I__10980\ : InMux
    port map (
            O => \N__49676\,
            I => \N__49670\
        );

    \I__10979\ : LocalMux
    port map (
            O => \N__49673\,
            I => \N__49666\
        );

    \I__10978\ : LocalMux
    port map (
            O => \N__49670\,
            I => \N__49663\
        );

    \I__10977\ : InMux
    port map (
            O => \N__49669\,
            I => \N__49660\
        );

    \I__10976\ : Span4Mux_v
    port map (
            O => \N__49666\,
            I => \N__49657\
        );

    \I__10975\ : Span4Mux_v
    port map (
            O => \N__49663\,
            I => \N__49654\
        );

    \I__10974\ : LocalMux
    port map (
            O => \N__49660\,
            I => \N__49651\
        );

    \I__10973\ : Span4Mux_h
    port map (
            O => \N__49657\,
            I => \N__49648\
        );

    \I__10972\ : Odrv4
    port map (
            O => \N__49654\,
            I => cemf_module_64ch_ctrl_inst1_data_config_3
        );

    \I__10971\ : Odrv4
    port map (
            O => \N__49651\,
            I => cemf_module_64ch_ctrl_inst1_data_config_3
        );

    \I__10970\ : Odrv4
    port map (
            O => \N__49648\,
            I => cemf_module_64ch_ctrl_inst1_data_config_3
        );

    \I__10969\ : InMux
    port map (
            O => \N__49641\,
            I => \N__49638\
        );

    \I__10968\ : LocalMux
    port map (
            O => \N__49638\,
            I => \N__49633\
        );

    \I__10967\ : InMux
    port map (
            O => \N__49637\,
            I => \N__49630\
        );

    \I__10966\ : CascadeMux
    port map (
            O => \N__49636\,
            I => \N__49627\
        );

    \I__10965\ : Span4Mux_v
    port map (
            O => \N__49633\,
            I => \N__49624\
        );

    \I__10964\ : LocalMux
    port map (
            O => \N__49630\,
            I => \N__49621\
        );

    \I__10963\ : InMux
    port map (
            O => \N__49627\,
            I => \N__49618\
        );

    \I__10962\ : Span4Mux_h
    port map (
            O => \N__49624\,
            I => \N__49615\
        );

    \I__10961\ : Span4Mux_v
    port map (
            O => \N__49621\,
            I => \N__49612\
        );

    \I__10960\ : LocalMux
    port map (
            O => \N__49618\,
            I => \N__49609\
        );

    \I__10959\ : Span4Mux_h
    port map (
            O => \N__49615\,
            I => \N__49602\
        );

    \I__10958\ : Span4Mux_v
    port map (
            O => \N__49612\,
            I => \N__49602\
        );

    \I__10957\ : Span4Mux_v
    port map (
            O => \N__49609\,
            I => \N__49602\
        );

    \I__10956\ : Odrv4
    port map (
            O => \N__49602\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_3
        );

    \I__10955\ : CascadeMux
    port map (
            O => \N__49599\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_3_cascade_\
        );

    \I__10954\ : InMux
    port map (
            O => \N__49596\,
            I => \N__49593\
        );

    \I__10953\ : LocalMux
    port map (
            O => \N__49593\,
            I => \N__49590\
        );

    \I__10952\ : Span4Mux_h
    port map (
            O => \N__49590\,
            I => \N__49587\
        );

    \I__10951\ : Span4Mux_h
    port map (
            O => \N__49587\,
            I => \N__49584\
        );

    \I__10950\ : Odrv4
    port map (
            O => \N__49584\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_3\
        );

    \I__10949\ : CascadeMux
    port map (
            O => \N__49581\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253QZ0Z5_cascade_\
        );

    \I__10948\ : InMux
    port map (
            O => \N__49578\,
            I => \N__49575\
        );

    \I__10947\ : LocalMux
    port map (
            O => \N__49575\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3\
        );

    \I__10946\ : CascadeMux
    port map (
            O => \N__49572\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLHZ0Z5_cascade_\
        );

    \I__10945\ : InMux
    port map (
            O => \N__49569\,
            I => \N__49566\
        );

    \I__10944\ : LocalMux
    port map (
            O => \N__49566\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23\
        );

    \I__10943\ : CascadeMux
    port map (
            O => \N__49563\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23_cascade_\
        );

    \I__10942\ : InMux
    port map (
            O => \N__49560\,
            I => \N__49557\
        );

    \I__10941\ : LocalMux
    port map (
            O => \N__49557\,
            I => \N__49554\
        );

    \I__10940\ : Span4Mux_v
    port map (
            O => \N__49554\,
            I => \N__49551\
        );

    \I__10939\ : Span4Mux_v
    port map (
            O => \N__49551\,
            I => \N__49548\
        );

    \I__10938\ : Sp12to4
    port map (
            O => \N__49548\,
            I => \N__49545\
        );

    \I__10937\ : Span12Mux_h
    port map (
            O => \N__49545\,
            I => \N__49542\
        );

    \I__10936\ : Odrv12
    port map (
            O => \N__49542\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.dout_conf\
        );

    \I__10935\ : CascadeMux
    port map (
            O => \N__49539\,
            I => \N__49536\
        );

    \I__10934\ : InMux
    port map (
            O => \N__49536\,
            I => \N__49533\
        );

    \I__10933\ : LocalMux
    port map (
            O => \N__49533\,
            I => \N__49530\
        );

    \I__10932\ : Odrv12
    port map (
            O => \N__49530\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALHZ0Z5\
        );

    \I__10931\ : InMux
    port map (
            O => \N__49527\,
            I => \N__49524\
        );

    \I__10930\ : LocalMux
    port map (
            O => \N__49524\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22\
        );

    \I__10929\ : InMux
    port map (
            O => \N__49521\,
            I => \N__49518\
        );

    \I__10928\ : LocalMux
    port map (
            O => \N__49518\,
            I => \N__49515\
        );

    \I__10927\ : Span4Mux_v
    port map (
            O => \N__49515\,
            I => \N__49512\
        );

    \I__10926\ : Sp12to4
    port map (
            O => \N__49512\,
            I => \N__49509\
        );

    \I__10925\ : Odrv12
    port map (
            O => \N__49509\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_21\
        );

    \I__10924\ : CascadeMux
    port map (
            O => \N__49506\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22_cascade_\
        );

    \I__10923\ : InMux
    port map (
            O => \N__49503\,
            I => \N__49500\
        );

    \I__10922\ : LocalMux
    port map (
            O => \N__49500\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_22\
        );

    \I__10921\ : InMux
    port map (
            O => \N__49497\,
            I => \N__49494\
        );

    \I__10920\ : LocalMux
    port map (
            O => \N__49494\,
            I => \N__49490\
        );

    \I__10919\ : CascadeMux
    port map (
            O => \N__49493\,
            I => \N__49487\
        );

    \I__10918\ : Span4Mux_h
    port map (
            O => \N__49490\,
            I => \N__49484\
        );

    \I__10917\ : InMux
    port map (
            O => \N__49487\,
            I => \N__49481\
        );

    \I__10916\ : Span4Mux_v
    port map (
            O => \N__49484\,
            I => \N__49477\
        );

    \I__10915\ : LocalMux
    port map (
            O => \N__49481\,
            I => \N__49474\
        );

    \I__10914\ : InMux
    port map (
            O => \N__49480\,
            I => \N__49471\
        );

    \I__10913\ : Odrv4
    port map (
            O => \N__49477\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_23
        );

    \I__10912\ : Odrv12
    port map (
            O => \N__49474\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_23
        );

    \I__10911\ : LocalMux
    port map (
            O => \N__49471\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_23
        );

    \I__10910\ : InMux
    port map (
            O => \N__49464\,
            I => \N__49461\
        );

    \I__10909\ : LocalMux
    port map (
            O => \N__49461\,
            I => \N__49458\
        );

    \I__10908\ : Span4Mux_h
    port map (
            O => \N__49458\,
            I => \N__49455\
        );

    \I__10907\ : Span4Mux_v
    port map (
            O => \N__49455\,
            I => \N__49450\
        );

    \I__10906\ : InMux
    port map (
            O => \N__49454\,
            I => \N__49447\
        );

    \I__10905\ : InMux
    port map (
            O => \N__49453\,
            I => \N__49444\
        );

    \I__10904\ : Odrv4
    port map (
            O => \N__49450\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_23
        );

    \I__10903\ : LocalMux
    port map (
            O => \N__49447\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_23
        );

    \I__10902\ : LocalMux
    port map (
            O => \N__49444\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_23
        );

    \I__10901\ : InMux
    port map (
            O => \N__49437\,
            I => \N__49434\
        );

    \I__10900\ : LocalMux
    port map (
            O => \N__49434\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_23\
        );

    \I__10899\ : CascadeMux
    port map (
            O => \N__49431\,
            I => \N__49428\
        );

    \I__10898\ : InMux
    port map (
            O => \N__49428\,
            I => \N__49424\
        );

    \I__10897\ : InMux
    port map (
            O => \N__49427\,
            I => \N__49420\
        );

    \I__10896\ : LocalMux
    port map (
            O => \N__49424\,
            I => \N__49417\
        );

    \I__10895\ : InMux
    port map (
            O => \N__49423\,
            I => \N__49414\
        );

    \I__10894\ : LocalMux
    port map (
            O => \N__49420\,
            I => \N__49411\
        );

    \I__10893\ : Span4Mux_h
    port map (
            O => \N__49417\,
            I => \N__49408\
        );

    \I__10892\ : LocalMux
    port map (
            O => \N__49414\,
            I => \N__49405\
        );

    \I__10891\ : Span4Mux_v
    port map (
            O => \N__49411\,
            I => \N__49402\
        );

    \I__10890\ : Span4Mux_v
    port map (
            O => \N__49408\,
            I => \N__49399\
        );

    \I__10889\ : Span4Mux_v
    port map (
            O => \N__49405\,
            I => \N__49394\
        );

    \I__10888\ : Span4Mux_h
    port map (
            O => \N__49402\,
            I => \N__49394\
        );

    \I__10887\ : Span4Mux_h
    port map (
            O => \N__49399\,
            I => \N__49391\
        );

    \I__10886\ : Odrv4
    port map (
            O => \N__49394\,
            I => cemf_module_64ch_ctrl_inst1_data_config_9
        );

    \I__10885\ : Odrv4
    port map (
            O => \N__49391\,
            I => cemf_module_64ch_ctrl_inst1_data_config_9
        );

    \I__10884\ : InMux
    port map (
            O => \N__49386\,
            I => \N__49383\
        );

    \I__10883\ : LocalMux
    port map (
            O => \N__49383\,
            I => \N__49379\
        );

    \I__10882\ : CascadeMux
    port map (
            O => \N__49382\,
            I => \N__49375\
        );

    \I__10881\ : Span4Mux_v
    port map (
            O => \N__49379\,
            I => \N__49372\
        );

    \I__10880\ : InMux
    port map (
            O => \N__49378\,
            I => \N__49369\
        );

    \I__10879\ : InMux
    port map (
            O => \N__49375\,
            I => \N__49366\
        );

    \I__10878\ : Span4Mux_h
    port map (
            O => \N__49372\,
            I => \N__49363\
        );

    \I__10877\ : LocalMux
    port map (
            O => \N__49369\,
            I => \N__49360\
        );

    \I__10876\ : LocalMux
    port map (
            O => \N__49366\,
            I => \N__49357\
        );

    \I__10875\ : Span4Mux_v
    port map (
            O => \N__49363\,
            I => \N__49354\
        );

    \I__10874\ : Span4Mux_h
    port map (
            O => \N__49360\,
            I => \N__49349\
        );

    \I__10873\ : Span4Mux_h
    port map (
            O => \N__49357\,
            I => \N__49349\
        );

    \I__10872\ : Odrv4
    port map (
            O => \N__49354\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_9
        );

    \I__10871\ : Odrv4
    port map (
            O => \N__49349\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_9
        );

    \I__10870\ : CascadeMux
    port map (
            O => \N__49344\,
            I => \N__49341\
        );

    \I__10869\ : InMux
    port map (
            O => \N__49341\,
            I => \N__49336\
        );

    \I__10868\ : InMux
    port map (
            O => \N__49340\,
            I => \N__49333\
        );

    \I__10867\ : CascadeMux
    port map (
            O => \N__49339\,
            I => \N__49330\
        );

    \I__10866\ : LocalMux
    port map (
            O => \N__49336\,
            I => \N__49327\
        );

    \I__10865\ : LocalMux
    port map (
            O => \N__49333\,
            I => \N__49324\
        );

    \I__10864\ : InMux
    port map (
            O => \N__49330\,
            I => \N__49321\
        );

    \I__10863\ : Span4Mux_h
    port map (
            O => \N__49327\,
            I => \N__49318\
        );

    \I__10862\ : Span12Mux_v
    port map (
            O => \N__49324\,
            I => \N__49313\
        );

    \I__10861\ : LocalMux
    port map (
            O => \N__49321\,
            I => \N__49313\
        );

    \I__10860\ : Odrv4
    port map (
            O => \N__49318\,
            I => cemf_module_64ch_ctrl_inst1_data_config_10
        );

    \I__10859\ : Odrv12
    port map (
            O => \N__49313\,
            I => cemf_module_64ch_ctrl_inst1_data_config_10
        );

    \I__10858\ : InMux
    port map (
            O => \N__49308\,
            I => \N__49304\
        );

    \I__10857\ : InMux
    port map (
            O => \N__49307\,
            I => \N__49301\
        );

    \I__10856\ : LocalMux
    port map (
            O => \N__49304\,
            I => \N__49298\
        );

    \I__10855\ : LocalMux
    port map (
            O => \N__49301\,
            I => \N__49295\
        );

    \I__10854\ : Span4Mux_v
    port map (
            O => \N__49298\,
            I => \N__49292\
        );

    \I__10853\ : Span4Mux_h
    port map (
            O => \N__49295\,
            I => \N__49289\
        );

    \I__10852\ : Span4Mux_h
    port map (
            O => \N__49292\,
            I => \N__49286\
        );

    \I__10851\ : Span4Mux_h
    port map (
            O => \N__49289\,
            I => \N__49282\
        );

    \I__10850\ : Sp12to4
    port map (
            O => \N__49286\,
            I => \N__49279\
        );

    \I__10849\ : InMux
    port map (
            O => \N__49285\,
            I => \N__49276\
        );

    \I__10848\ : Odrv4
    port map (
            O => \N__49282\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_10
        );

    \I__10847\ : Odrv12
    port map (
            O => \N__49279\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_10
        );

    \I__10846\ : LocalMux
    port map (
            O => \N__49276\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_10
        );

    \I__10845\ : InMux
    port map (
            O => \N__49269\,
            I => \N__49265\
        );

    \I__10844\ : InMux
    port map (
            O => \N__49268\,
            I => \N__49262\
        );

    \I__10843\ : LocalMux
    port map (
            O => \N__49265\,
            I => \N__49259\
        );

    \I__10842\ : LocalMux
    port map (
            O => \N__49262\,
            I => \N__49256\
        );

    \I__10841\ : Span4Mux_v
    port map (
            O => \N__49259\,
            I => \N__49252\
        );

    \I__10840\ : Span4Mux_v
    port map (
            O => \N__49256\,
            I => \N__49249\
        );

    \I__10839\ : CascadeMux
    port map (
            O => \N__49255\,
            I => \N__49246\
        );

    \I__10838\ : Span4Mux_h
    port map (
            O => \N__49252\,
            I => \N__49241\
        );

    \I__10837\ : Span4Mux_h
    port map (
            O => \N__49249\,
            I => \N__49241\
        );

    \I__10836\ : InMux
    port map (
            O => \N__49246\,
            I => \N__49238\
        );

    \I__10835\ : Odrv4
    port map (
            O => \N__49241\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_10
        );

    \I__10834\ : LocalMux
    port map (
            O => \N__49238\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_10
        );

    \I__10833\ : CascadeMux
    port map (
            O => \N__49233\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_10_cascade_\
        );

    \I__10832\ : InMux
    port map (
            O => \N__49230\,
            I => \N__49227\
        );

    \I__10831\ : LocalMux
    port map (
            O => \N__49227\,
            I => \N__49224\
        );

    \I__10830\ : Span4Mux_v
    port map (
            O => \N__49224\,
            I => \N__49221\
        );

    \I__10829\ : Odrv4
    port map (
            O => \N__49221\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_10\
        );

    \I__10828\ : CascadeMux
    port map (
            O => \N__49218\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFHZ0Z5_cascade_\
        );

    \I__10827\ : InMux
    port map (
            O => \N__49215\,
            I => \N__49212\
        );

    \I__10826\ : LocalMux
    port map (
            O => \N__49212\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10\
        );

    \I__10825\ : CascadeMux
    port map (
            O => \N__49209\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9DZ0Z7_cascade_\
        );

    \I__10824\ : InMux
    port map (
            O => \N__49206\,
            I => \N__49203\
        );

    \I__10823\ : LocalMux
    port map (
            O => \N__49203\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19\
        );

    \I__10822\ : CascadeMux
    port map (
            O => \N__49200\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19_cascade_\
        );

    \I__10821\ : InMux
    port map (
            O => \N__49197\,
            I => \N__49194\
        );

    \I__10820\ : LocalMux
    port map (
            O => \N__49194\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_18\
        );

    \I__10819\ : InMux
    port map (
            O => \N__49191\,
            I => \N__49188\
        );

    \I__10818\ : LocalMux
    port map (
            O => \N__49188\,
            I => \N__49185\
        );

    \I__10817\ : Span4Mux_h
    port map (
            O => \N__49185\,
            I => \N__49182\
        );

    \I__10816\ : Span4Mux_h
    port map (
            O => \N__49182\,
            I => \N__49179\
        );

    \I__10815\ : Span4Mux_v
    port map (
            O => \N__49179\,
            I => \N__49176\
        );

    \I__10814\ : Odrv4
    port map (
            O => \N__49176\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_19\
        );

    \I__10813\ : InMux
    port map (
            O => \N__49173\,
            I => \N__49170\
        );

    \I__10812\ : LocalMux
    port map (
            O => \N__49170\,
            I => \N__49167\
        );

    \I__10811\ : Span4Mux_h
    port map (
            O => \N__49167\,
            I => \N__49164\
        );

    \I__10810\ : Span4Mux_h
    port map (
            O => \N__49164\,
            I => \N__49160\
        );

    \I__10809\ : CascadeMux
    port map (
            O => \N__49163\,
            I => \N__49157\
        );

    \I__10808\ : Span4Mux_h
    port map (
            O => \N__49160\,
            I => \N__49153\
        );

    \I__10807\ : InMux
    port map (
            O => \N__49157\,
            I => \N__49148\
        );

    \I__10806\ : InMux
    port map (
            O => \N__49156\,
            I => \N__49148\
        );

    \I__10805\ : Odrv4
    port map (
            O => \N__49153\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_18
        );

    \I__10804\ : LocalMux
    port map (
            O => \N__49148\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_18
        );

    \I__10803\ : InMux
    port map (
            O => \N__49143\,
            I => \N__49140\
        );

    \I__10802\ : LocalMux
    port map (
            O => \N__49140\,
            I => \N__49137\
        );

    \I__10801\ : Span4Mux_v
    port map (
            O => \N__49137\,
            I => \N__49134\
        );

    \I__10800\ : Span4Mux_v
    port map (
            O => \N__49134\,
            I => \N__49131\
        );

    \I__10799\ : Odrv4
    port map (
            O => \N__49131\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_27\
        );

    \I__10798\ : InMux
    port map (
            O => \N__49128\,
            I => \N__49125\
        );

    \I__10797\ : LocalMux
    port map (
            O => \N__49125\,
            I => \N__49122\
        );

    \I__10796\ : Span4Mux_h
    port map (
            O => \N__49122\,
            I => \N__49119\
        );

    \I__10795\ : Span4Mux_h
    port map (
            O => \N__49119\,
            I => \N__49116\
        );

    \I__10794\ : Span4Mux_h
    port map (
            O => \N__49116\,
            I => \N__49113\
        );

    \I__10793\ : Odrv4
    port map (
            O => \N__49113\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_28\
        );

    \I__10792\ : InMux
    port map (
            O => \N__49110\,
            I => \N__49107\
        );

    \I__10791\ : LocalMux
    port map (
            O => \N__49107\,
            I => \N__49104\
        );

    \I__10790\ : Span4Mux_h
    port map (
            O => \N__49104\,
            I => \N__49101\
        );

    \I__10789\ : Span4Mux_v
    port map (
            O => \N__49101\,
            I => \N__49098\
        );

    \I__10788\ : Odrv4
    port map (
            O => \N__49098\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_29\
        );

    \I__10787\ : CEMux
    port map (
            O => \N__49095\,
            I => \N__49090\
        );

    \I__10786\ : CEMux
    port map (
            O => \N__49094\,
            I => \N__49087\
        );

    \I__10785\ : CEMux
    port map (
            O => \N__49093\,
            I => \N__49084\
        );

    \I__10784\ : LocalMux
    port map (
            O => \N__49090\,
            I => \N__49080\
        );

    \I__10783\ : LocalMux
    port map (
            O => \N__49087\,
            I => \N__49075\
        );

    \I__10782\ : LocalMux
    port map (
            O => \N__49084\,
            I => \N__49075\
        );

    \I__10781\ : CEMux
    port map (
            O => \N__49083\,
            I => \N__49072\
        );

    \I__10780\ : Span4Mux_v
    port map (
            O => \N__49080\,
            I => \N__49064\
        );

    \I__10779\ : Span4Mux_v
    port map (
            O => \N__49075\,
            I => \N__49064\
        );

    \I__10778\ : LocalMux
    port map (
            O => \N__49072\,
            I => \N__49064\
        );

    \I__10777\ : CEMux
    port map (
            O => \N__49071\,
            I => \N__49060\
        );

    \I__10776\ : Span4Mux_h
    port map (
            O => \N__49064\,
            I => \N__49056\
        );

    \I__10775\ : CEMux
    port map (
            O => \N__49063\,
            I => \N__49053\
        );

    \I__10774\ : LocalMux
    port map (
            O => \N__49060\,
            I => \N__49050\
        );

    \I__10773\ : CEMux
    port map (
            O => \N__49059\,
            I => \N__49047\
        );

    \I__10772\ : Span4Mux_v
    port map (
            O => \N__49056\,
            I => \N__49044\
        );

    \I__10771\ : LocalMux
    port map (
            O => \N__49053\,
            I => \N__49041\
        );

    \I__10770\ : Span4Mux_v
    port map (
            O => \N__49050\,
            I => \N__49038\
        );

    \I__10769\ : LocalMux
    port map (
            O => \N__49047\,
            I => \N__49035\
        );

    \I__10768\ : Span4Mux_h
    port map (
            O => \N__49044\,
            I => \N__49028\
        );

    \I__10767\ : Span4Mux_h
    port map (
            O => \N__49041\,
            I => \N__49028\
        );

    \I__10766\ : Span4Mux_h
    port map (
            O => \N__49038\,
            I => \N__49023\
        );

    \I__10765\ : Span4Mux_h
    port map (
            O => \N__49035\,
            I => \N__49023\
        );

    \I__10764\ : CEMux
    port map (
            O => \N__49034\,
            I => \N__49020\
        );

    \I__10763\ : CEMux
    port map (
            O => \N__49033\,
            I => \N__49017\
        );

    \I__10762\ : Odrv4
    port map (
            O => \N__49028\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0\
        );

    \I__10761\ : Odrv4
    port map (
            O => \N__49023\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0\
        );

    \I__10760\ : LocalMux
    port map (
            O => \N__49020\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0\
        );

    \I__10759\ : LocalMux
    port map (
            O => \N__49017\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0\
        );

    \I__10758\ : CascadeMux
    port map (
            O => \N__49008\,
            I => \N__49005\
        );

    \I__10757\ : InMux
    port map (
            O => \N__49005\,
            I => \N__49000\
        );

    \I__10756\ : InMux
    port map (
            O => \N__49004\,
            I => \N__48997\
        );

    \I__10755\ : InMux
    port map (
            O => \N__49003\,
            I => \N__48994\
        );

    \I__10754\ : LocalMux
    port map (
            O => \N__49000\,
            I => \N__48991\
        );

    \I__10753\ : LocalMux
    port map (
            O => \N__48997\,
            I => \N__48988\
        );

    \I__10752\ : LocalMux
    port map (
            O => \N__48994\,
            I => \N__48985\
        );

    \I__10751\ : Span4Mux_h
    port map (
            O => \N__48991\,
            I => \N__48982\
        );

    \I__10750\ : Odrv12
    port map (
            O => \N__48988\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_23
        );

    \I__10749\ : Odrv4
    port map (
            O => \N__48985\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_23
        );

    \I__10748\ : Odrv4
    port map (
            O => \N__48982\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_23
        );

    \I__10747\ : InMux
    port map (
            O => \N__48975\,
            I => \N__48971\
        );

    \I__10746\ : InMux
    port map (
            O => \N__48974\,
            I => \N__48968\
        );

    \I__10745\ : LocalMux
    port map (
            O => \N__48971\,
            I => \N__48965\
        );

    \I__10744\ : LocalMux
    port map (
            O => \N__48968\,
            I => \N__48961\
        );

    \I__10743\ : Span4Mux_h
    port map (
            O => \N__48965\,
            I => \N__48958\
        );

    \I__10742\ : InMux
    port map (
            O => \N__48964\,
            I => \N__48955\
        );

    \I__10741\ : Span4Mux_h
    port map (
            O => \N__48961\,
            I => \N__48950\
        );

    \I__10740\ : Span4Mux_h
    port map (
            O => \N__48958\,
            I => \N__48950\
        );

    \I__10739\ : LocalMux
    port map (
            O => \N__48955\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_23
        );

    \I__10738\ : Odrv4
    port map (
            O => \N__48950\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_23
        );

    \I__10737\ : CascadeMux
    port map (
            O => \N__48945\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_23_cascade_\
        );

    \I__10736\ : InMux
    port map (
            O => \N__48942\,
            I => \N__48939\
        );

    \I__10735\ : LocalMux
    port map (
            O => \N__48939\,
            I => \N__48936\
        );

    \I__10734\ : Span4Mux_h
    port map (
            O => \N__48936\,
            I => \N__48931\
        );

    \I__10733\ : InMux
    port map (
            O => \N__48935\,
            I => \N__48926\
        );

    \I__10732\ : InMux
    port map (
            O => \N__48934\,
            I => \N__48926\
        );

    \I__10731\ : Odrv4
    port map (
            O => \N__48931\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_0
        );

    \I__10730\ : LocalMux
    port map (
            O => \N__48926\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_0
        );

    \I__10729\ : InMux
    port map (
            O => \N__48921\,
            I => \N__48918\
        );

    \I__10728\ : LocalMux
    port map (
            O => \N__48918\,
            I => \N__48915\
        );

    \I__10727\ : Span4Mux_h
    port map (
            O => \N__48915\,
            I => \N__48911\
        );

    \I__10726\ : CascadeMux
    port map (
            O => \N__48914\,
            I => \N__48907\
        );

    \I__10725\ : Span4Mux_h
    port map (
            O => \N__48911\,
            I => \N__48904\
        );

    \I__10724\ : InMux
    port map (
            O => \N__48910\,
            I => \N__48901\
        );

    \I__10723\ : InMux
    port map (
            O => \N__48907\,
            I => \N__48898\
        );

    \I__10722\ : Odrv4
    port map (
            O => \N__48904\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_0
        );

    \I__10721\ : LocalMux
    port map (
            O => \N__48901\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_0
        );

    \I__10720\ : LocalMux
    port map (
            O => \N__48898\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_0
        );

    \I__10719\ : InMux
    port map (
            O => \N__48891\,
            I => \N__48888\
        );

    \I__10718\ : LocalMux
    port map (
            O => \N__48888\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_0\
        );

    \I__10717\ : CascadeMux
    port map (
            O => \N__48885\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_0_cascade_\
        );

    \I__10716\ : CascadeMux
    port map (
            O => \N__48882\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQLZ0Z7_cascade_\
        );

    \I__10715\ : InMux
    port map (
            O => \N__48879\,
            I => \N__48875\
        );

    \I__10714\ : InMux
    port map (
            O => \N__48878\,
            I => \N__48872\
        );

    \I__10713\ : LocalMux
    port map (
            O => \N__48875\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0\
        );

    \I__10712\ : LocalMux
    port map (
            O => \N__48872\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0\
        );

    \I__10711\ : CascadeMux
    port map (
            O => \N__48867\,
            I => \N__48863\
        );

    \I__10710\ : InMux
    port map (
            O => \N__48866\,
            I => \N__48859\
        );

    \I__10709\ : InMux
    port map (
            O => \N__48863\,
            I => \N__48856\
        );

    \I__10708\ : InMux
    port map (
            O => \N__48862\,
            I => \N__48853\
        );

    \I__10707\ : LocalMux
    port map (
            O => \N__48859\,
            I => \N__48848\
        );

    \I__10706\ : LocalMux
    port map (
            O => \N__48856\,
            I => \N__48848\
        );

    \I__10705\ : LocalMux
    port map (
            O => \N__48853\,
            I => \N__48845\
        );

    \I__10704\ : Span4Mux_v
    port map (
            O => \N__48848\,
            I => \N__48842\
        );

    \I__10703\ : Odrv12
    port map (
            O => \N__48845\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_18
        );

    \I__10702\ : Odrv4
    port map (
            O => \N__48842\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_18
        );

    \I__10701\ : CascadeMux
    port map (
            O => \N__48837\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_18_cascade_\
        );

    \I__10700\ : InMux
    port map (
            O => \N__48834\,
            I => \N__48831\
        );

    \I__10699\ : LocalMux
    port map (
            O => \N__48831\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_18\
        );

    \I__10698\ : CascadeMux
    port map (
            O => \N__48828\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579DZ0Z7_cascade_\
        );

    \I__10697\ : InMux
    port map (
            O => \N__48825\,
            I => \N__48822\
        );

    \I__10696\ : LocalMux
    port map (
            O => \N__48822\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18\
        );

    \I__10695\ : InMux
    port map (
            O => \N__48819\,
            I => \N__48816\
        );

    \I__10694\ : LocalMux
    port map (
            O => \N__48816\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_17\
        );

    \I__10693\ : CascadeMux
    port map (
            O => \N__48813\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18_cascade_\
        );

    \I__10692\ : CascadeMux
    port map (
            O => \N__48810\,
            I => \N__48807\
        );

    \I__10691\ : InMux
    port map (
            O => \N__48807\,
            I => \N__48804\
        );

    \I__10690\ : LocalMux
    port map (
            O => \N__48804\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_19\
        );

    \I__10689\ : InMux
    port map (
            O => \N__48801\,
            I => \N__48798\
        );

    \I__10688\ : LocalMux
    port map (
            O => \N__48798\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_19\
        );

    \I__10687\ : CascadeMux
    port map (
            O => \N__48795\,
            I => \N__48792\
        );

    \I__10686\ : InMux
    port map (
            O => \N__48792\,
            I => \N__48789\
        );

    \I__10685\ : LocalMux
    port map (
            O => \N__48789\,
            I => \N__48786\
        );

    \I__10684\ : Span4Mux_v
    port map (
            O => \N__48786\,
            I => \N__48783\
        );

    \I__10683\ : Span4Mux_h
    port map (
            O => \N__48783\,
            I => \N__48780\
        );

    \I__10682\ : Span4Mux_h
    port map (
            O => \N__48780\,
            I => \N__48777\
        );

    \I__10681\ : Odrv4
    port map (
            O => \N__48777\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_28\
        );

    \I__10680\ : CascadeMux
    port map (
            O => \N__48774\,
            I => \N__48771\
        );

    \I__10679\ : InMux
    port map (
            O => \N__48771\,
            I => \N__48768\
        );

    \I__10678\ : LocalMux
    port map (
            O => \N__48768\,
            I => \N__48765\
        );

    \I__10677\ : Span4Mux_h
    port map (
            O => \N__48765\,
            I => \N__48762\
        );

    \I__10676\ : Odrv4
    port map (
            O => \N__48762\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_29\
        );

    \I__10675\ : InMux
    port map (
            O => \N__48759\,
            I => \N__48756\
        );

    \I__10674\ : LocalMux
    port map (
            O => \N__48756\,
            I => \N__48753\
        );

    \I__10673\ : Span4Mux_v
    port map (
            O => \N__48753\,
            I => \N__48750\
        );

    \I__10672\ : Sp12to4
    port map (
            O => \N__48750\,
            I => \N__48746\
        );

    \I__10671\ : InMux
    port map (
            O => \N__48749\,
            I => \N__48742\
        );

    \I__10670\ : Span12Mux_h
    port map (
            O => \N__48746\,
            I => \N__48739\
        );

    \I__10669\ : InMux
    port map (
            O => \N__48745\,
            I => \N__48736\
        );

    \I__10668\ : LocalMux
    port map (
            O => \N__48742\,
            I => \N__48733\
        );

    \I__10667\ : Odrv12
    port map (
            O => \N__48739\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_7
        );

    \I__10666\ : LocalMux
    port map (
            O => \N__48736\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_7
        );

    \I__10665\ : Odrv4
    port map (
            O => \N__48733\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_7
        );

    \I__10664\ : CEMux
    port map (
            O => \N__48726\,
            I => \N__48711\
        );

    \I__10663\ : CEMux
    port map (
            O => \N__48725\,
            I => \N__48711\
        );

    \I__10662\ : CEMux
    port map (
            O => \N__48724\,
            I => \N__48711\
        );

    \I__10661\ : CEMux
    port map (
            O => \N__48723\,
            I => \N__48711\
        );

    \I__10660\ : CEMux
    port map (
            O => \N__48722\,
            I => \N__48711\
        );

    \I__10659\ : GlobalMux
    port map (
            O => \N__48711\,
            I => \N__48708\
        );

    \I__10658\ : gio2CtrlBuf
    port map (
            O => \N__48708\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g\
        );

    \I__10657\ : InMux
    port map (
            O => \N__48705\,
            I => \N__48702\
        );

    \I__10656\ : LocalMux
    port map (
            O => \N__48702\,
            I => \N__48698\
        );

    \I__10655\ : CascadeMux
    port map (
            O => \N__48701\,
            I => \N__48695\
        );

    \I__10654\ : Span4Mux_v
    port map (
            O => \N__48698\,
            I => \N__48691\
        );

    \I__10653\ : InMux
    port map (
            O => \N__48695\,
            I => \N__48686\
        );

    \I__10652\ : InMux
    port map (
            O => \N__48694\,
            I => \N__48686\
        );

    \I__10651\ : Odrv4
    port map (
            O => \N__48691\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_19
        );

    \I__10650\ : LocalMux
    port map (
            O => \N__48686\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_19
        );

    \I__10649\ : InMux
    port map (
            O => \N__48681\,
            I => \N__48678\
        );

    \I__10648\ : LocalMux
    port map (
            O => \N__48678\,
            I => \N__48674\
        );

    \I__10647\ : CascadeMux
    port map (
            O => \N__48677\,
            I => \N__48671\
        );

    \I__10646\ : Span12Mux_s10_v
    port map (
            O => \N__48674\,
            I => \N__48667\
        );

    \I__10645\ : InMux
    port map (
            O => \N__48671\,
            I => \N__48664\
        );

    \I__10644\ : InMux
    port map (
            O => \N__48670\,
            I => \N__48661\
        );

    \I__10643\ : Odrv12
    port map (
            O => \N__48667\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_19
        );

    \I__10642\ : LocalMux
    port map (
            O => \N__48664\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_19
        );

    \I__10641\ : LocalMux
    port map (
            O => \N__48661\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_19
        );

    \I__10640\ : InMux
    port map (
            O => \N__48654\,
            I => \N__48642\
        );

    \I__10639\ : InMux
    port map (
            O => \N__48653\,
            I => \N__48642\
        );

    \I__10638\ : InMux
    port map (
            O => \N__48652\,
            I => \N__48642\
        );

    \I__10637\ : InMux
    port map (
            O => \N__48651\,
            I => \N__48642\
        );

    \I__10636\ : LocalMux
    port map (
            O => \N__48642\,
            I => \N__48635\
        );

    \I__10635\ : InMux
    port map (
            O => \N__48641\,
            I => \N__48626\
        );

    \I__10634\ : InMux
    port map (
            O => \N__48640\,
            I => \N__48626\
        );

    \I__10633\ : InMux
    port map (
            O => \N__48639\,
            I => \N__48626\
        );

    \I__10632\ : InMux
    port map (
            O => \N__48638\,
            I => \N__48626\
        );

    \I__10631\ : Odrv4
    port map (
            O => \N__48635\,
            I => \serializer_mod_inst.next_state32_i\
        );

    \I__10630\ : LocalMux
    port map (
            O => \N__48626\,
            I => \serializer_mod_inst.next_state32_i\
        );

    \I__10629\ : InMux
    port map (
            O => \N__48621\,
            I => \serializer_mod_inst.counter_sr_cry_6\
        );

    \I__10628\ : InMux
    port map (
            O => \N__48618\,
            I => \N__48613\
        );

    \I__10627\ : InMux
    port map (
            O => \N__48617\,
            I => \N__48610\
        );

    \I__10626\ : InMux
    port map (
            O => \N__48616\,
            I => \N__48607\
        );

    \I__10625\ : LocalMux
    port map (
            O => \N__48613\,
            I => \serializer_mod_inst.counter_srZ0Z_7\
        );

    \I__10624\ : LocalMux
    port map (
            O => \N__48610\,
            I => \serializer_mod_inst.counter_srZ0Z_7\
        );

    \I__10623\ : LocalMux
    port map (
            O => \N__48607\,
            I => \serializer_mod_inst.counter_srZ0Z_7\
        );

    \I__10622\ : CEMux
    port map (
            O => \N__48600\,
            I => \N__48597\
        );

    \I__10621\ : LocalMux
    port map (
            O => \N__48597\,
            I => \N__48594\
        );

    \I__10620\ : Span4Mux_v
    port map (
            O => \N__48594\,
            I => \N__48591\
        );

    \I__10619\ : Span4Mux_h
    port map (
            O => \N__48591\,
            I => \N__48588\
        );

    \I__10618\ : Odrv4
    port map (
            O => \N__48588\,
            I => \serializer_mod_inst.counter_sre_0_i\
        );

    \I__10617\ : CascadeMux
    port map (
            O => \N__48585\,
            I => \N__48582\
        );

    \I__10616\ : InMux
    port map (
            O => \N__48582\,
            I => \N__48578\
        );

    \I__10615\ : InMux
    port map (
            O => \N__48581\,
            I => \N__48575\
        );

    \I__10614\ : LocalMux
    port map (
            O => \N__48578\,
            I => \N__48572\
        );

    \I__10613\ : LocalMux
    port map (
            O => \N__48575\,
            I => \N__48569\
        );

    \I__10612\ : Span4Mux_v
    port map (
            O => \N__48572\,
            I => \N__48566\
        );

    \I__10611\ : Span4Mux_v
    port map (
            O => \N__48569\,
            I => \N__48562\
        );

    \I__10610\ : Span4Mux_v
    port map (
            O => \N__48566\,
            I => \N__48559\
        );

    \I__10609\ : CascadeMux
    port map (
            O => \N__48565\,
            I => \N__48556\
        );

    \I__10608\ : Span4Mux_h
    port map (
            O => \N__48562\,
            I => \N__48551\
        );

    \I__10607\ : Span4Mux_h
    port map (
            O => \N__48559\,
            I => \N__48551\
        );

    \I__10606\ : InMux
    port map (
            O => \N__48556\,
            I => \N__48548\
        );

    \I__10605\ : Span4Mux_h
    port map (
            O => \N__48551\,
            I => \N__48545\
        );

    \I__10604\ : LocalMux
    port map (
            O => \N__48548\,
            I => \N__48542\
        );

    \I__10603\ : Odrv4
    port map (
            O => \N__48545\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_15
        );

    \I__10602\ : Odrv4
    port map (
            O => \N__48542\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_15
        );

    \I__10601\ : CascadeMux
    port map (
            O => \N__48537\,
            I => \N__48534\
        );

    \I__10600\ : InMux
    port map (
            O => \N__48534\,
            I => \N__48531\
        );

    \I__10599\ : LocalMux
    port map (
            O => \N__48531\,
            I => \N__48528\
        );

    \I__10598\ : Span4Mux_v
    port map (
            O => \N__48528\,
            I => \N__48525\
        );

    \I__10597\ : Span4Mux_h
    port map (
            O => \N__48525\,
            I => \N__48522\
        );

    \I__10596\ : Odrv4
    port map (
            O => \N__48522\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_24\
        );

    \I__10595\ : InMux
    port map (
            O => \N__48519\,
            I => \N__48516\
        );

    \I__10594\ : LocalMux
    port map (
            O => \N__48516\,
            I => \N__48513\
        );

    \I__10593\ : Span4Mux_v
    port map (
            O => \N__48513\,
            I => \N__48510\
        );

    \I__10592\ : Span4Mux_h
    port map (
            O => \N__48510\,
            I => \N__48507\
        );

    \I__10591\ : Odrv4
    port map (
            O => \N__48507\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_2Z0Z_26\
        );

    \I__10590\ : CascadeMux
    port map (
            O => \N__48504\,
            I => \N__48501\
        );

    \I__10589\ : InMux
    port map (
            O => \N__48501\,
            I => \N__48498\
        );

    \I__10588\ : LocalMux
    port map (
            O => \N__48498\,
            I => \N__48495\
        );

    \I__10587\ : Span4Mux_h
    port map (
            O => \N__48495\,
            I => \N__48492\
        );

    \I__10586\ : Odrv4
    port map (
            O => \N__48492\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_27\
        );

    \I__10585\ : InMux
    port map (
            O => \N__48489\,
            I => \N__48486\
        );

    \I__10584\ : LocalMux
    port map (
            O => \N__48486\,
            I => \serializer_mod_inst.un22_next_state_5\
        );

    \I__10583\ : InMux
    port map (
            O => \N__48483\,
            I => \N__48479\
        );

    \I__10582\ : InMux
    port map (
            O => \N__48482\,
            I => \N__48475\
        );

    \I__10581\ : LocalMux
    port map (
            O => \N__48479\,
            I => \N__48472\
        );

    \I__10580\ : InMux
    port map (
            O => \N__48478\,
            I => \N__48469\
        );

    \I__10579\ : LocalMux
    port map (
            O => \N__48475\,
            I => \serializer_mod_inst.counter_srZ0Z_0\
        );

    \I__10578\ : Odrv4
    port map (
            O => \N__48472\,
            I => \serializer_mod_inst.counter_srZ0Z_0\
        );

    \I__10577\ : LocalMux
    port map (
            O => \N__48469\,
            I => \serializer_mod_inst.counter_srZ0Z_0\
        );

    \I__10576\ : InMux
    port map (
            O => \N__48462\,
            I => \bfn_21_27_0_\
        );

    \I__10575\ : CascadeMux
    port map (
            O => \N__48459\,
            I => \N__48454\
        );

    \I__10574\ : InMux
    port map (
            O => \N__48458\,
            I => \N__48451\
        );

    \I__10573\ : InMux
    port map (
            O => \N__48457\,
            I => \N__48448\
        );

    \I__10572\ : InMux
    port map (
            O => \N__48454\,
            I => \N__48445\
        );

    \I__10571\ : LocalMux
    port map (
            O => \N__48451\,
            I => \serializer_mod_inst.counter_srZ0Z_1\
        );

    \I__10570\ : LocalMux
    port map (
            O => \N__48448\,
            I => \serializer_mod_inst.counter_srZ0Z_1\
        );

    \I__10569\ : LocalMux
    port map (
            O => \N__48445\,
            I => \serializer_mod_inst.counter_srZ0Z_1\
        );

    \I__10568\ : InMux
    port map (
            O => \N__48438\,
            I => \serializer_mod_inst.counter_sr_cry_0\
        );

    \I__10567\ : InMux
    port map (
            O => \N__48435\,
            I => \N__48431\
        );

    \I__10566\ : InMux
    port map (
            O => \N__48434\,
            I => \N__48427\
        );

    \I__10565\ : LocalMux
    port map (
            O => \N__48431\,
            I => \N__48424\
        );

    \I__10564\ : InMux
    port map (
            O => \N__48430\,
            I => \N__48421\
        );

    \I__10563\ : LocalMux
    port map (
            O => \N__48427\,
            I => \serializer_mod_inst.counter_srZ0Z_2\
        );

    \I__10562\ : Odrv4
    port map (
            O => \N__48424\,
            I => \serializer_mod_inst.counter_srZ0Z_2\
        );

    \I__10561\ : LocalMux
    port map (
            O => \N__48421\,
            I => \serializer_mod_inst.counter_srZ0Z_2\
        );

    \I__10560\ : InMux
    port map (
            O => \N__48414\,
            I => \serializer_mod_inst.counter_sr_cry_1\
        );

    \I__10559\ : InMux
    port map (
            O => \N__48411\,
            I => \N__48406\
        );

    \I__10558\ : InMux
    port map (
            O => \N__48410\,
            I => \N__48401\
        );

    \I__10557\ : InMux
    port map (
            O => \N__48409\,
            I => \N__48401\
        );

    \I__10556\ : LocalMux
    port map (
            O => \N__48406\,
            I => \serializer_mod_inst.counter_srZ0Z_3\
        );

    \I__10555\ : LocalMux
    port map (
            O => \N__48401\,
            I => \serializer_mod_inst.counter_srZ0Z_3\
        );

    \I__10554\ : InMux
    port map (
            O => \N__48396\,
            I => \serializer_mod_inst.counter_sr_cry_2\
        );

    \I__10553\ : InMux
    port map (
            O => \N__48393\,
            I => \N__48388\
        );

    \I__10552\ : InMux
    port map (
            O => \N__48392\,
            I => \N__48383\
        );

    \I__10551\ : InMux
    port map (
            O => \N__48391\,
            I => \N__48383\
        );

    \I__10550\ : LocalMux
    port map (
            O => \N__48388\,
            I => \serializer_mod_inst.counter_srZ0Z_4\
        );

    \I__10549\ : LocalMux
    port map (
            O => \N__48383\,
            I => \serializer_mod_inst.counter_srZ0Z_4\
        );

    \I__10548\ : InMux
    port map (
            O => \N__48378\,
            I => \serializer_mod_inst.counter_sr_cry_3\
        );

    \I__10547\ : InMux
    port map (
            O => \N__48375\,
            I => \N__48370\
        );

    \I__10546\ : InMux
    port map (
            O => \N__48374\,
            I => \N__48365\
        );

    \I__10545\ : InMux
    port map (
            O => \N__48373\,
            I => \N__48365\
        );

    \I__10544\ : LocalMux
    port map (
            O => \N__48370\,
            I => \serializer_mod_inst.counter_srZ0Z_5\
        );

    \I__10543\ : LocalMux
    port map (
            O => \N__48365\,
            I => \serializer_mod_inst.counter_srZ0Z_5\
        );

    \I__10542\ : InMux
    port map (
            O => \N__48360\,
            I => \serializer_mod_inst.counter_sr_cry_4\
        );

    \I__10541\ : InMux
    port map (
            O => \N__48357\,
            I => \N__48352\
        );

    \I__10540\ : CascadeMux
    port map (
            O => \N__48356\,
            I => \N__48349\
        );

    \I__10539\ : InMux
    port map (
            O => \N__48355\,
            I => \N__48346\
        );

    \I__10538\ : LocalMux
    port map (
            O => \N__48352\,
            I => \N__48343\
        );

    \I__10537\ : InMux
    port map (
            O => \N__48349\,
            I => \N__48340\
        );

    \I__10536\ : LocalMux
    port map (
            O => \N__48346\,
            I => \serializer_mod_inst.counter_srZ0Z_6\
        );

    \I__10535\ : Odrv4
    port map (
            O => \N__48343\,
            I => \serializer_mod_inst.counter_srZ0Z_6\
        );

    \I__10534\ : LocalMux
    port map (
            O => \N__48340\,
            I => \serializer_mod_inst.counter_srZ0Z_6\
        );

    \I__10533\ : InMux
    port map (
            O => \N__48333\,
            I => \serializer_mod_inst.counter_sr_cry_5\
        );

    \I__10532\ : CascadeMux
    port map (
            O => \N__48330\,
            I => \N__48326\
        );

    \I__10531\ : InMux
    port map (
            O => \N__48329\,
            I => \N__48322\
        );

    \I__10530\ : InMux
    port map (
            O => \N__48326\,
            I => \N__48317\
        );

    \I__10529\ : InMux
    port map (
            O => \N__48325\,
            I => \N__48317\
        );

    \I__10528\ : LocalMux
    port map (
            O => \N__48322\,
            I => \N__48314\
        );

    \I__10527\ : LocalMux
    port map (
            O => \N__48317\,
            I => \N__48311\
        );

    \I__10526\ : Span12Mux_v
    port map (
            O => \N__48314\,
            I => \N__48307\
        );

    \I__10525\ : Span4Mux_h
    port map (
            O => \N__48311\,
            I => \N__48304\
        );

    \I__10524\ : InMux
    port map (
            O => \N__48310\,
            I => \N__48301\
        );

    \I__10523\ : Odrv12
    port map (
            O => \N__48307\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0\
        );

    \I__10522\ : Odrv4
    port map (
            O => \N__48304\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0\
        );

    \I__10521\ : LocalMux
    port map (
            O => \N__48301\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0\
        );

    \I__10520\ : InMux
    port map (
            O => \N__48294\,
            I => \N__48287\
        );

    \I__10519\ : InMux
    port map (
            O => \N__48293\,
            I => \N__48284\
        );

    \I__10518\ : InMux
    port map (
            O => \N__48292\,
            I => \N__48281\
        );

    \I__10517\ : InMux
    port map (
            O => \N__48291\,
            I => \N__48278\
        );

    \I__10516\ : InMux
    port map (
            O => \N__48290\,
            I => \N__48275\
        );

    \I__10515\ : LocalMux
    port map (
            O => \N__48287\,
            I => \N__48272\
        );

    \I__10514\ : LocalMux
    port map (
            O => \N__48284\,
            I => \N__48263\
        );

    \I__10513\ : LocalMux
    port map (
            O => \N__48281\,
            I => \N__48263\
        );

    \I__10512\ : LocalMux
    port map (
            O => \N__48278\,
            I => \N__48263\
        );

    \I__10511\ : LocalMux
    port map (
            O => \N__48275\,
            I => \N__48263\
        );

    \I__10510\ : Span4Mux_v
    port map (
            O => \N__48272\,
            I => \N__48259\
        );

    \I__10509\ : Span4Mux_v
    port map (
            O => \N__48263\,
            I => \N__48253\
        );

    \I__10508\ : InMux
    port map (
            O => \N__48262\,
            I => \N__48250\
        );

    \I__10507\ : Span4Mux_h
    port map (
            O => \N__48259\,
            I => \N__48247\
        );

    \I__10506\ : InMux
    port map (
            O => \N__48258\,
            I => \N__48244\
        );

    \I__10505\ : InMux
    port map (
            O => \N__48257\,
            I => \N__48241\
        );

    \I__10504\ : InMux
    port map (
            O => \N__48256\,
            I => \N__48238\
        );

    \I__10503\ : Span4Mux_h
    port map (
            O => \N__48253\,
            I => \N__48235\
        );

    \I__10502\ : LocalMux
    port map (
            O => \N__48250\,
            I => \I2C_top_level_inst1.s_data_ireg_0\
        );

    \I__10501\ : Odrv4
    port map (
            O => \N__48247\,
            I => \I2C_top_level_inst1.s_data_ireg_0\
        );

    \I__10500\ : LocalMux
    port map (
            O => \N__48244\,
            I => \I2C_top_level_inst1.s_data_ireg_0\
        );

    \I__10499\ : LocalMux
    port map (
            O => \N__48241\,
            I => \I2C_top_level_inst1.s_data_ireg_0\
        );

    \I__10498\ : LocalMux
    port map (
            O => \N__48238\,
            I => \I2C_top_level_inst1.s_data_ireg_0\
        );

    \I__10497\ : Odrv4
    port map (
            O => \N__48235\,
            I => \I2C_top_level_inst1.s_data_ireg_0\
        );

    \I__10496\ : CascadeMux
    port map (
            O => \N__48222\,
            I => \N__48216\
        );

    \I__10495\ : CascadeMux
    port map (
            O => \N__48221\,
            I => \N__48213\
        );

    \I__10494\ : CascadeMux
    port map (
            O => \N__48220\,
            I => \N__48210\
        );

    \I__10493\ : CascadeMux
    port map (
            O => \N__48219\,
            I => \N__48206\
        );

    \I__10492\ : InMux
    port map (
            O => \N__48216\,
            I => \N__48196\
        );

    \I__10491\ : InMux
    port map (
            O => \N__48213\,
            I => \N__48196\
        );

    \I__10490\ : InMux
    port map (
            O => \N__48210\,
            I => \N__48196\
        );

    \I__10489\ : InMux
    port map (
            O => \N__48209\,
            I => \N__48196\
        );

    \I__10488\ : InMux
    port map (
            O => \N__48206\,
            I => \N__48190\
        );

    \I__10487\ : InMux
    port map (
            O => \N__48205\,
            I => \N__48190\
        );

    \I__10486\ : LocalMux
    port map (
            O => \N__48196\,
            I => \N__48187\
        );

    \I__10485\ : InMux
    port map (
            O => \N__48195\,
            I => \N__48184\
        );

    \I__10484\ : LocalMux
    port map (
            O => \N__48190\,
            I => \N__48174\
        );

    \I__10483\ : Span4Mux_h
    port map (
            O => \N__48187\,
            I => \N__48174\
        );

    \I__10482\ : LocalMux
    port map (
            O => \N__48184\,
            I => \N__48174\
        );

    \I__10481\ : InMux
    port map (
            O => \N__48183\,
            I => \N__48167\
        );

    \I__10480\ : InMux
    port map (
            O => \N__48182\,
            I => \N__48167\
        );

    \I__10479\ : InMux
    port map (
            O => \N__48181\,
            I => \N__48167\
        );

    \I__10478\ : Odrv4
    port map (
            O => \N__48174\,
            I => \I2C_top_level_inst1.s_command_0\
        );

    \I__10477\ : LocalMux
    port map (
            O => \N__48167\,
            I => \I2C_top_level_inst1.s_command_0\
        );

    \I__10476\ : InMux
    port map (
            O => \N__48162\,
            I => \N__48159\
        );

    \I__10475\ : LocalMux
    port map (
            O => \N__48159\,
            I => \N__48153\
        );

    \I__10474\ : InMux
    port map (
            O => \N__48158\,
            I => \N__48150\
        );

    \I__10473\ : InMux
    port map (
            O => \N__48157\,
            I => \N__48147\
        );

    \I__10472\ : InMux
    port map (
            O => \N__48156\,
            I => \N__48144\
        );

    \I__10471\ : Span4Mux_v
    port map (
            O => \N__48153\,
            I => \N__48141\
        );

    \I__10470\ : LocalMux
    port map (
            O => \N__48150\,
            I => \N__48133\
        );

    \I__10469\ : LocalMux
    port map (
            O => \N__48147\,
            I => \N__48133\
        );

    \I__10468\ : LocalMux
    port map (
            O => \N__48144\,
            I => \N__48133\
        );

    \I__10467\ : Span4Mux_h
    port map (
            O => \N__48141\,
            I => \N__48129\
        );

    \I__10466\ : InMux
    port map (
            O => \N__48140\,
            I => \N__48126\
        );

    \I__10465\ : Span4Mux_v
    port map (
            O => \N__48133\,
            I => \N__48123\
        );

    \I__10464\ : InMux
    port map (
            O => \N__48132\,
            I => \N__48120\
        );

    \I__10463\ : Odrv4
    port map (
            O => \N__48129\,
            I => \I2C_top_level_inst1.s_data_ireg_1\
        );

    \I__10462\ : LocalMux
    port map (
            O => \N__48126\,
            I => \I2C_top_level_inst1.s_data_ireg_1\
        );

    \I__10461\ : Odrv4
    port map (
            O => \N__48123\,
            I => \I2C_top_level_inst1.s_data_ireg_1\
        );

    \I__10460\ : LocalMux
    port map (
            O => \N__48120\,
            I => \I2C_top_level_inst1.s_data_ireg_1\
        );

    \I__10459\ : InMux
    port map (
            O => \N__48111\,
            I => \N__48108\
        );

    \I__10458\ : LocalMux
    port map (
            O => \N__48108\,
            I => \N__48102\
        );

    \I__10457\ : InMux
    port map (
            O => \N__48107\,
            I => \N__48099\
        );

    \I__10456\ : InMux
    port map (
            O => \N__48106\,
            I => \N__48096\
        );

    \I__10455\ : InMux
    port map (
            O => \N__48105\,
            I => \N__48093\
        );

    \I__10454\ : Span4Mux_v
    port map (
            O => \N__48102\,
            I => \N__48090\
        );

    \I__10453\ : LocalMux
    port map (
            O => \N__48099\,
            I => \N__48085\
        );

    \I__10452\ : LocalMux
    port map (
            O => \N__48096\,
            I => \N__48085\
        );

    \I__10451\ : LocalMux
    port map (
            O => \N__48093\,
            I => \N__48082\
        );

    \I__10450\ : Span4Mux_h
    port map (
            O => \N__48090\,
            I => \N__48077\
        );

    \I__10449\ : Span4Mux_v
    port map (
            O => \N__48085\,
            I => \N__48074\
        );

    \I__10448\ : Span4Mux_v
    port map (
            O => \N__48082\,
            I => \N__48071\
        );

    \I__10447\ : InMux
    port map (
            O => \N__48081\,
            I => \N__48066\
        );

    \I__10446\ : InMux
    port map (
            O => \N__48080\,
            I => \N__48066\
        );

    \I__10445\ : Odrv4
    port map (
            O => \N__48077\,
            I => \I2C_top_level_inst1.s_data_ireg_2\
        );

    \I__10444\ : Odrv4
    port map (
            O => \N__48074\,
            I => \I2C_top_level_inst1.s_data_ireg_2\
        );

    \I__10443\ : Odrv4
    port map (
            O => \N__48071\,
            I => \I2C_top_level_inst1.s_data_ireg_2\
        );

    \I__10442\ : LocalMux
    port map (
            O => \N__48066\,
            I => \I2C_top_level_inst1.s_data_ireg_2\
        );

    \I__10441\ : InMux
    port map (
            O => \N__48057\,
            I => \N__48053\
        );

    \I__10440\ : InMux
    port map (
            O => \N__48056\,
            I => \N__48050\
        );

    \I__10439\ : LocalMux
    port map (
            O => \N__48053\,
            I => \N__48045\
        );

    \I__10438\ : LocalMux
    port map (
            O => \N__48050\,
            I => \N__48042\
        );

    \I__10437\ : InMux
    port map (
            O => \N__48049\,
            I => \N__48039\
        );

    \I__10436\ : InMux
    port map (
            O => \N__48048\,
            I => \N__48036\
        );

    \I__10435\ : Span4Mux_v
    port map (
            O => \N__48045\,
            I => \N__48033\
        );

    \I__10434\ : Span4Mux_v
    port map (
            O => \N__48042\,
            I => \N__48029\
        );

    \I__10433\ : LocalMux
    port map (
            O => \N__48039\,
            I => \N__48024\
        );

    \I__10432\ : LocalMux
    port map (
            O => \N__48036\,
            I => \N__48024\
        );

    \I__10431\ : Span4Mux_v
    port map (
            O => \N__48033\,
            I => \N__48021\
        );

    \I__10430\ : InMux
    port map (
            O => \N__48032\,
            I => \N__48017\
        );

    \I__10429\ : Span4Mux_h
    port map (
            O => \N__48029\,
            I => \N__48014\
        );

    \I__10428\ : Span4Mux_v
    port map (
            O => \N__48024\,
            I => \N__48009\
        );

    \I__10427\ : Span4Mux_h
    port map (
            O => \N__48021\,
            I => \N__48009\
        );

    \I__10426\ : InMux
    port map (
            O => \N__48020\,
            I => \N__48006\
        );

    \I__10425\ : LocalMux
    port map (
            O => \N__48017\,
            I => \I2C_top_level_inst1.s_data_ireg_3\
        );

    \I__10424\ : Odrv4
    port map (
            O => \N__48014\,
            I => \I2C_top_level_inst1.s_data_ireg_3\
        );

    \I__10423\ : Odrv4
    port map (
            O => \N__48009\,
            I => \I2C_top_level_inst1.s_data_ireg_3\
        );

    \I__10422\ : LocalMux
    port map (
            O => \N__48006\,
            I => \I2C_top_level_inst1.s_data_ireg_3\
        );

    \I__10421\ : ClkMux
    port map (
            O => \N__47997\,
            I => \N__47937\
        );

    \I__10420\ : ClkMux
    port map (
            O => \N__47996\,
            I => \N__47937\
        );

    \I__10419\ : ClkMux
    port map (
            O => \N__47995\,
            I => \N__47937\
        );

    \I__10418\ : ClkMux
    port map (
            O => \N__47994\,
            I => \N__47937\
        );

    \I__10417\ : ClkMux
    port map (
            O => \N__47993\,
            I => \N__47937\
        );

    \I__10416\ : ClkMux
    port map (
            O => \N__47992\,
            I => \N__47937\
        );

    \I__10415\ : ClkMux
    port map (
            O => \N__47991\,
            I => \N__47937\
        );

    \I__10414\ : ClkMux
    port map (
            O => \N__47990\,
            I => \N__47937\
        );

    \I__10413\ : ClkMux
    port map (
            O => \N__47989\,
            I => \N__47937\
        );

    \I__10412\ : ClkMux
    port map (
            O => \N__47988\,
            I => \N__47937\
        );

    \I__10411\ : ClkMux
    port map (
            O => \N__47987\,
            I => \N__47937\
        );

    \I__10410\ : ClkMux
    port map (
            O => \N__47986\,
            I => \N__47937\
        );

    \I__10409\ : ClkMux
    port map (
            O => \N__47985\,
            I => \N__47937\
        );

    \I__10408\ : ClkMux
    port map (
            O => \N__47984\,
            I => \N__47937\
        );

    \I__10407\ : ClkMux
    port map (
            O => \N__47983\,
            I => \N__47937\
        );

    \I__10406\ : ClkMux
    port map (
            O => \N__47982\,
            I => \N__47937\
        );

    \I__10405\ : ClkMux
    port map (
            O => \N__47981\,
            I => \N__47937\
        );

    \I__10404\ : ClkMux
    port map (
            O => \N__47980\,
            I => \N__47937\
        );

    \I__10403\ : ClkMux
    port map (
            O => \N__47979\,
            I => \N__47937\
        );

    \I__10402\ : ClkMux
    port map (
            O => \N__47978\,
            I => \N__47937\
        );

    \I__10401\ : GlobalMux
    port map (
            O => \N__47937\,
            I => \N__47934\
        );

    \I__10400\ : gio2CtrlBuf
    port map (
            O => \N__47934\,
            I => scl_c_g
        );

    \I__10399\ : CEMux
    port map (
            O => \N__47931\,
            I => \N__47928\
        );

    \I__10398\ : LocalMux
    port map (
            O => \N__47928\,
            I => \N__47925\
        );

    \I__10397\ : Span4Mux_h
    port map (
            O => \N__47925\,
            I => \N__47922\
        );

    \I__10396\ : Span4Mux_h
    port map (
            O => \N__47922\,
            I => \N__47918\
        );

    \I__10395\ : CEMux
    port map (
            O => \N__47921\,
            I => \N__47915\
        );

    \I__10394\ : Sp12to4
    port map (
            O => \N__47918\,
            I => \N__47907\
        );

    \I__10393\ : LocalMux
    port map (
            O => \N__47915\,
            I => \N__47907\
        );

    \I__10392\ : InMux
    port map (
            O => \N__47914\,
            I => \N__47904\
        );

    \I__10391\ : InMux
    port map (
            O => \N__47913\,
            I => \N__47899\
        );

    \I__10390\ : InMux
    port map (
            O => \N__47912\,
            I => \N__47899\
        );

    \I__10389\ : Odrv12
    port map (
            O => \N__47907\,
            I => \I2C_top_level_inst1.s_load_command\
        );

    \I__10388\ : LocalMux
    port map (
            O => \N__47904\,
            I => \I2C_top_level_inst1.s_load_command\
        );

    \I__10387\ : LocalMux
    port map (
            O => \N__47899\,
            I => \I2C_top_level_inst1.s_load_command\
        );

    \I__10386\ : InMux
    port map (
            O => \N__47892\,
            I => \N__47889\
        );

    \I__10385\ : LocalMux
    port map (
            O => \N__47889\,
            I => \serializer_mod_inst.un1_counter_srlto6_3\
        );

    \I__10384\ : CascadeMux
    port map (
            O => \N__47886\,
            I => \serializer_mod_inst.un1_counter_srlto6_4_cascade_\
        );

    \I__10383\ : InMux
    port map (
            O => \N__47883\,
            I => \N__47860\
        );

    \I__10382\ : InMux
    port map (
            O => \N__47882\,
            I => \N__47833\
        );

    \I__10381\ : InMux
    port map (
            O => \N__47881\,
            I => \N__47833\
        );

    \I__10380\ : InMux
    port map (
            O => \N__47880\,
            I => \N__47833\
        );

    \I__10379\ : InMux
    port map (
            O => \N__47879\,
            I => \N__47833\
        );

    \I__10378\ : InMux
    port map (
            O => \N__47878\,
            I => \N__47828\
        );

    \I__10377\ : InMux
    port map (
            O => \N__47877\,
            I => \N__47828\
        );

    \I__10376\ : InMux
    port map (
            O => \N__47876\,
            I => \N__47823\
        );

    \I__10375\ : InMux
    port map (
            O => \N__47875\,
            I => \N__47823\
        );

    \I__10374\ : InMux
    port map (
            O => \N__47874\,
            I => \N__47820\
        );

    \I__10373\ : InMux
    port map (
            O => \N__47873\,
            I => \N__47815\
        );

    \I__10372\ : InMux
    port map (
            O => \N__47872\,
            I => \N__47815\
        );

    \I__10371\ : InMux
    port map (
            O => \N__47871\,
            I => \N__47803\
        );

    \I__10370\ : InMux
    port map (
            O => \N__47870\,
            I => \N__47803\
        );

    \I__10369\ : InMux
    port map (
            O => \N__47869\,
            I => \N__47803\
        );

    \I__10368\ : InMux
    port map (
            O => \N__47868\,
            I => \N__47798\
        );

    \I__10367\ : InMux
    port map (
            O => \N__47867\,
            I => \N__47798\
        );

    \I__10366\ : InMux
    port map (
            O => \N__47866\,
            I => \N__47795\
        );

    \I__10365\ : InMux
    port map (
            O => \N__47865\,
            I => \N__47788\
        );

    \I__10364\ : InMux
    port map (
            O => \N__47864\,
            I => \N__47788\
        );

    \I__10363\ : InMux
    port map (
            O => \N__47863\,
            I => \N__47788\
        );

    \I__10362\ : LocalMux
    port map (
            O => \N__47860\,
            I => \N__47785\
        );

    \I__10361\ : InMux
    port map (
            O => \N__47859\,
            I => \N__47778\
        );

    \I__10360\ : InMux
    port map (
            O => \N__47858\,
            I => \N__47778\
        );

    \I__10359\ : InMux
    port map (
            O => \N__47857\,
            I => \N__47778\
        );

    \I__10358\ : InMux
    port map (
            O => \N__47856\,
            I => \N__47771\
        );

    \I__10357\ : InMux
    port map (
            O => \N__47855\,
            I => \N__47771\
        );

    \I__10356\ : InMux
    port map (
            O => \N__47854\,
            I => \N__47771\
        );

    \I__10355\ : InMux
    port map (
            O => \N__47853\,
            I => \N__47764\
        );

    \I__10354\ : InMux
    port map (
            O => \N__47852\,
            I => \N__47764\
        );

    \I__10353\ : InMux
    port map (
            O => \N__47851\,
            I => \N__47764\
        );

    \I__10352\ : InMux
    port map (
            O => \N__47850\,
            I => \N__47759\
        );

    \I__10351\ : InMux
    port map (
            O => \N__47849\,
            I => \N__47759\
        );

    \I__10350\ : InMux
    port map (
            O => \N__47848\,
            I => \N__47756\
        );

    \I__10349\ : InMux
    port map (
            O => \N__47847\,
            I => \N__47743\
        );

    \I__10348\ : InMux
    port map (
            O => \N__47846\,
            I => \N__47743\
        );

    \I__10347\ : InMux
    port map (
            O => \N__47845\,
            I => \N__47743\
        );

    \I__10346\ : InMux
    port map (
            O => \N__47844\,
            I => \N__47743\
        );

    \I__10345\ : InMux
    port map (
            O => \N__47843\,
            I => \N__47743\
        );

    \I__10344\ : InMux
    port map (
            O => \N__47842\,
            I => \N__47743\
        );

    \I__10343\ : LocalMux
    port map (
            O => \N__47833\,
            I => \N__47732\
        );

    \I__10342\ : LocalMux
    port map (
            O => \N__47828\,
            I => \N__47732\
        );

    \I__10341\ : LocalMux
    port map (
            O => \N__47823\,
            I => \N__47732\
        );

    \I__10340\ : LocalMux
    port map (
            O => \N__47820\,
            I => \N__47732\
        );

    \I__10339\ : LocalMux
    port map (
            O => \N__47815\,
            I => \N__47721\
        );

    \I__10338\ : InMux
    port map (
            O => \N__47814\,
            I => \N__47716\
        );

    \I__10337\ : InMux
    port map (
            O => \N__47813\,
            I => \N__47716\
        );

    \I__10336\ : InMux
    port map (
            O => \N__47812\,
            I => \N__47711\
        );

    \I__10335\ : InMux
    port map (
            O => \N__47811\,
            I => \N__47711\
        );

    \I__10334\ : InMux
    port map (
            O => \N__47810\,
            I => \N__47708\
        );

    \I__10333\ : LocalMux
    port map (
            O => \N__47803\,
            I => \N__47703\
        );

    \I__10332\ : LocalMux
    port map (
            O => \N__47798\,
            I => \N__47696\
        );

    \I__10331\ : LocalMux
    port map (
            O => \N__47795\,
            I => \N__47696\
        );

    \I__10330\ : LocalMux
    port map (
            O => \N__47788\,
            I => \N__47696\
        );

    \I__10329\ : Span4Mux_h
    port map (
            O => \N__47785\,
            I => \N__47681\
        );

    \I__10328\ : LocalMux
    port map (
            O => \N__47778\,
            I => \N__47681\
        );

    \I__10327\ : LocalMux
    port map (
            O => \N__47771\,
            I => \N__47681\
        );

    \I__10326\ : LocalMux
    port map (
            O => \N__47764\,
            I => \N__47681\
        );

    \I__10325\ : LocalMux
    port map (
            O => \N__47759\,
            I => \N__47681\
        );

    \I__10324\ : LocalMux
    port map (
            O => \N__47756\,
            I => \N__47681\
        );

    \I__10323\ : LocalMux
    port map (
            O => \N__47743\,
            I => \N__47681\
        );

    \I__10322\ : InMux
    port map (
            O => \N__47742\,
            I => \N__47676\
        );

    \I__10321\ : InMux
    port map (
            O => \N__47741\,
            I => \N__47676\
        );

    \I__10320\ : Span4Mux_v
    port map (
            O => \N__47732\,
            I => \N__47673\
        );

    \I__10319\ : InMux
    port map (
            O => \N__47731\,
            I => \N__47664\
        );

    \I__10318\ : InMux
    port map (
            O => \N__47730\,
            I => \N__47664\
        );

    \I__10317\ : InMux
    port map (
            O => \N__47729\,
            I => \N__47664\
        );

    \I__10316\ : InMux
    port map (
            O => \N__47728\,
            I => \N__47664\
        );

    \I__10315\ : InMux
    port map (
            O => \N__47727\,
            I => \N__47655\
        );

    \I__10314\ : InMux
    port map (
            O => \N__47726\,
            I => \N__47655\
        );

    \I__10313\ : InMux
    port map (
            O => \N__47725\,
            I => \N__47655\
        );

    \I__10312\ : InMux
    port map (
            O => \N__47724\,
            I => \N__47655\
        );

    \I__10311\ : Span4Mux_h
    port map (
            O => \N__47721\,
            I => \N__47639\
        );

    \I__10310\ : LocalMux
    port map (
            O => \N__47716\,
            I => \N__47639\
        );

    \I__10309\ : LocalMux
    port map (
            O => \N__47711\,
            I => \N__47634\
        );

    \I__10308\ : LocalMux
    port map (
            O => \N__47708\,
            I => \N__47634\
        );

    \I__10307\ : InMux
    port map (
            O => \N__47707\,
            I => \N__47629\
        );

    \I__10306\ : InMux
    port map (
            O => \N__47706\,
            I => \N__47629\
        );

    \I__10305\ : Span4Mux_h
    port map (
            O => \N__47703\,
            I => \N__47620\
        );

    \I__10304\ : Span4Mux_v
    port map (
            O => \N__47696\,
            I => \N__47620\
        );

    \I__10303\ : Span4Mux_v
    port map (
            O => \N__47681\,
            I => \N__47620\
        );

    \I__10302\ : LocalMux
    port map (
            O => \N__47676\,
            I => \N__47620\
        );

    \I__10301\ : Span4Mux_h
    port map (
            O => \N__47673\,
            I => \N__47613\
        );

    \I__10300\ : LocalMux
    port map (
            O => \N__47664\,
            I => \N__47613\
        );

    \I__10299\ : LocalMux
    port map (
            O => \N__47655\,
            I => \N__47613\
        );

    \I__10298\ : InMux
    port map (
            O => \N__47654\,
            I => \N__47602\
        );

    \I__10297\ : InMux
    port map (
            O => \N__47653\,
            I => \N__47602\
        );

    \I__10296\ : InMux
    port map (
            O => \N__47652\,
            I => \N__47602\
        );

    \I__10295\ : InMux
    port map (
            O => \N__47651\,
            I => \N__47602\
        );

    \I__10294\ : InMux
    port map (
            O => \N__47650\,
            I => \N__47602\
        );

    \I__10293\ : InMux
    port map (
            O => \N__47649\,
            I => \N__47591\
        );

    \I__10292\ : InMux
    port map (
            O => \N__47648\,
            I => \N__47591\
        );

    \I__10291\ : InMux
    port map (
            O => \N__47647\,
            I => \N__47591\
        );

    \I__10290\ : InMux
    port map (
            O => \N__47646\,
            I => \N__47591\
        );

    \I__10289\ : InMux
    port map (
            O => \N__47645\,
            I => \N__47591\
        );

    \I__10288\ : InMux
    port map (
            O => \N__47644\,
            I => \N__47588\
        );

    \I__10287\ : Odrv4
    port map (
            O => \N__47639\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10286\ : Odrv12
    port map (
            O => \N__47634\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10285\ : LocalMux
    port map (
            O => \N__47629\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10284\ : Odrv4
    port map (
            O => \N__47620\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10283\ : Odrv4
    port map (
            O => \N__47613\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10282\ : LocalMux
    port map (
            O => \N__47602\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10281\ : LocalMux
    port map (
            O => \N__47591\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10280\ : LocalMux
    port map (
            O => \N__47588\,
            I => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\
        );

    \I__10279\ : CascadeMux
    port map (
            O => \N__47571\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_10_cascade_\
        );

    \I__10278\ : CascadeMux
    port map (
            O => \N__47568\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_18_cascade_\
        );

    \I__10277\ : InMux
    port map (
            O => \N__47565\,
            I => \N__47557\
        );

    \I__10276\ : InMux
    port map (
            O => \N__47564\,
            I => \N__47557\
        );

    \I__10275\ : InMux
    port map (
            O => \N__47563\,
            I => \N__47552\
        );

    \I__10274\ : InMux
    port map (
            O => \N__47562\,
            I => \N__47552\
        );

    \I__10273\ : LocalMux
    port map (
            O => \N__47557\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18\
        );

    \I__10272\ : LocalMux
    port map (
            O => \N__47552\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18\
        );

    \I__10271\ : InMux
    port map (
            O => \N__47547\,
            I => \N__47538\
        );

    \I__10270\ : InMux
    port map (
            O => \N__47546\,
            I => \N__47538\
        );

    \I__10269\ : InMux
    port map (
            O => \N__47545\,
            I => \N__47538\
        );

    \I__10268\ : LocalMux
    port map (
            O => \N__47538\,
            I => \N__47535\
        );

    \I__10267\ : Span4Mux_h
    port map (
            O => \N__47535\,
            I => \N__47532\
        );

    \I__10266\ : Span4Mux_v
    port map (
            O => \N__47532\,
            I => \N__47529\
        );

    \I__10265\ : Odrv4
    port map (
            O => \N__47529\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1605_0\
        );

    \I__10264\ : InMux
    port map (
            O => \N__47526\,
            I => \N__47523\
        );

    \I__10263\ : LocalMux
    port map (
            O => \N__47523\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0\
        );

    \I__10262\ : CascadeMux
    port map (
            O => \N__47520\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0_cascade_\
        );

    \I__10261\ : InMux
    port map (
            O => \N__47517\,
            I => \N__47514\
        );

    \I__10260\ : LocalMux
    port map (
            O => \N__47514\,
            I => \N__47511\
        );

    \I__10259\ : Span4Mux_v
    port map (
            O => \N__47511\,
            I => \N__47507\
        );

    \I__10258\ : InMux
    port map (
            O => \N__47510\,
            I => \N__47504\
        );

    \I__10257\ : Span4Mux_v
    port map (
            O => \N__47507\,
            I => \N__47501\
        );

    \I__10256\ : LocalMux
    port map (
            O => \N__47504\,
            I => \N__47498\
        );

    \I__10255\ : Odrv4
    port map (
            O => \N__47501\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0\
        );

    \I__10254\ : Odrv4
    port map (
            O => \N__47498\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0\
        );

    \I__10253\ : InMux
    port map (
            O => \N__47493\,
            I => \N__47490\
        );

    \I__10252\ : LocalMux
    port map (
            O => \N__47490\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_0_1_14\
        );

    \I__10251\ : CascadeMux
    port map (
            O => \N__47487\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_279_cascade_\
        );

    \I__10250\ : CascadeMux
    port map (
            O => \N__47484\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_0_1_7_cascade_\
        );

    \I__10249\ : CascadeMux
    port map (
            O => \N__47481\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_268_cascade_\
        );

    \I__10248\ : InMux
    port map (
            O => \N__47478\,
            I => \N__47475\
        );

    \I__10247\ : LocalMux
    port map (
            O => \N__47475\,
            I => \N__47472\
        );

    \I__10246\ : Odrv4
    port map (
            O => \N__47472\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_7_3_i_a2_0\
        );

    \I__10245\ : InMux
    port map (
            O => \N__47469\,
            I => \N__47463\
        );

    \I__10244\ : InMux
    port map (
            O => \N__47468\,
            I => \N__47463\
        );

    \I__10243\ : LocalMux
    port map (
            O => \N__47463\,
            I => \N__47460\
        );

    \I__10242\ : Span4Mux_h
    port map (
            O => \N__47460\,
            I => \N__47457\
        );

    \I__10241\ : Span4Mux_h
    port map (
            O => \N__47457\,
            I => \N__47453\
        );

    \I__10240\ : InMux
    port map (
            O => \N__47456\,
            I => \N__47450\
        );

    \I__10239\ : Odrv4
    port map (
            O => \N__47453\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0\
        );

    \I__10238\ : LocalMux
    port map (
            O => \N__47450\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0\
        );

    \I__10237\ : InMux
    port map (
            O => \N__47445\,
            I => \N__47442\
        );

    \I__10236\ : LocalMux
    port map (
            O => \N__47442\,
            I => \N__47439\
        );

    \I__10235\ : Odrv12
    port map (
            O => \N__47439\,
            I => \I2C_top_level_inst1.s_addr1_o_0\
        );

    \I__10234\ : CascadeMux
    port map (
            O => \N__47436\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0_cascade_\
        );

    \I__10233\ : InMux
    port map (
            O => \N__47433\,
            I => \N__47430\
        );

    \I__10232\ : LocalMux
    port map (
            O => \N__47430\,
            I => \N__47427\
        );

    \I__10231\ : Span4Mux_h
    port map (
            O => \N__47427\,
            I => \N__47423\
        );

    \I__10230\ : InMux
    port map (
            O => \N__47426\,
            I => \N__47420\
        );

    \I__10229\ : Odrv4
    port map (
            O => \N__47423\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1\
        );

    \I__10228\ : LocalMux
    port map (
            O => \N__47420\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1\
        );

    \I__10227\ : InMux
    port map (
            O => \N__47415\,
            I => \N__47404\
        );

    \I__10226\ : InMux
    port map (
            O => \N__47414\,
            I => \N__47404\
        );

    \I__10225\ : InMux
    port map (
            O => \N__47413\,
            I => \N__47400\
        );

    \I__10224\ : InMux
    port map (
            O => \N__47412\,
            I => \N__47391\
        );

    \I__10223\ : InMux
    port map (
            O => \N__47411\,
            I => \N__47391\
        );

    \I__10222\ : InMux
    port map (
            O => \N__47410\,
            I => \N__47391\
        );

    \I__10221\ : InMux
    port map (
            O => \N__47409\,
            I => \N__47391\
        );

    \I__10220\ : LocalMux
    port map (
            O => \N__47404\,
            I => \N__47388\
        );

    \I__10219\ : CascadeMux
    port map (
            O => \N__47403\,
            I => \N__47385\
        );

    \I__10218\ : LocalMux
    port map (
            O => \N__47400\,
            I => \N__47375\
        );

    \I__10217\ : LocalMux
    port map (
            O => \N__47391\,
            I => \N__47372\
        );

    \I__10216\ : Span4Mux_h
    port map (
            O => \N__47388\,
            I => \N__47369\
        );

    \I__10215\ : InMux
    port map (
            O => \N__47385\,
            I => \N__47366\
        );

    \I__10214\ : InMux
    port map (
            O => \N__47384\,
            I => \N__47357\
        );

    \I__10213\ : InMux
    port map (
            O => \N__47383\,
            I => \N__47357\
        );

    \I__10212\ : InMux
    port map (
            O => \N__47382\,
            I => \N__47357\
        );

    \I__10211\ : InMux
    port map (
            O => \N__47381\,
            I => \N__47357\
        );

    \I__10210\ : InMux
    port map (
            O => \N__47380\,
            I => \N__47350\
        );

    \I__10209\ : InMux
    port map (
            O => \N__47379\,
            I => \N__47350\
        );

    \I__10208\ : InMux
    port map (
            O => \N__47378\,
            I => \N__47350\
        );

    \I__10207\ : Span4Mux_h
    port map (
            O => \N__47375\,
            I => \N__47347\
        );

    \I__10206\ : Span4Mux_h
    port map (
            O => \N__47372\,
            I => \N__47344\
        );

    \I__10205\ : Sp12to4
    port map (
            O => \N__47369\,
            I => \N__47341\
        );

    \I__10204\ : LocalMux
    port map (
            O => \N__47366\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\
        );

    \I__10203\ : LocalMux
    port map (
            O => \N__47357\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\
        );

    \I__10202\ : LocalMux
    port map (
            O => \N__47350\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\
        );

    \I__10201\ : Odrv4
    port map (
            O => \N__47347\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\
        );

    \I__10200\ : Odrv4
    port map (
            O => \N__47344\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\
        );

    \I__10199\ : Odrv12
    port map (
            O => \N__47341\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\
        );

    \I__10198\ : CascadeMux
    port map (
            O => \N__47328\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_8_cascade_\
        );

    \I__10197\ : InMux
    port map (
            O => \N__47325\,
            I => \N__47322\
        );

    \I__10196\ : LocalMux
    port map (
            O => \N__47322\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_CO\
        );

    \I__10195\ : InMux
    port map (
            O => \N__47319\,
            I => \N__47316\
        );

    \I__10194\ : LocalMux
    port map (
            O => \N__47316\,
            I => \N__47313\
        );

    \I__10193\ : Span4Mux_v
    port map (
            O => \N__47313\,
            I => \N__47310\
        );

    \I__10192\ : Odrv4
    port map (
            O => \N__47310\,
            I => \I2C_top_level_inst1.s_addr0_o_1\
        );

    \I__10191\ : CascadeMux
    port map (
            O => \N__47307\,
            I => \N__47304\
        );

    \I__10190\ : InMux
    port map (
            O => \N__47304\,
            I => \N__47301\
        );

    \I__10189\ : LocalMux
    port map (
            O => \N__47301\,
            I => \N__47298\
        );

    \I__10188\ : Span4Mux_v
    port map (
            O => \N__47298\,
            I => \N__47295\
        );

    \I__10187\ : Span4Mux_h
    port map (
            O => \N__47295\,
            I => \N__47292\
        );

    \I__10186\ : Span4Mux_v
    port map (
            O => \N__47292\,
            I => \N__47289\
        );

    \I__10185\ : Odrv4
    port map (
            O => \N__47289\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1651\
        );

    \I__10184\ : InMux
    port map (
            O => \N__47286\,
            I => \N__47283\
        );

    \I__10183\ : LocalMux
    port map (
            O => \N__47283\,
            I => \N__47280\
        );

    \I__10182\ : Span4Mux_h
    port map (
            O => \N__47280\,
            I => \N__47277\
        );

    \I__10181\ : Span4Mux_h
    port map (
            O => \N__47277\,
            I => \N__47274\
        );

    \I__10180\ : Odrv4
    port map (
            O => \N__47274\,
            I => \I2C_top_level_inst1.s_addr0_o_2\
        );

    \I__10179\ : CascadeMux
    port map (
            O => \N__47271\,
            I => \N__47268\
        );

    \I__10178\ : InMux
    port map (
            O => \N__47268\,
            I => \N__47265\
        );

    \I__10177\ : LocalMux
    port map (
            O => \N__47265\,
            I => \N__47262\
        );

    \I__10176\ : Span4Mux_h
    port map (
            O => \N__47262\,
            I => \N__47259\
        );

    \I__10175\ : Sp12to4
    port map (
            O => \N__47259\,
            I => \N__47256\
        );

    \I__10174\ : Span12Mux_v
    port map (
            O => \N__47256\,
            I => \N__47253\
        );

    \I__10173\ : Odrv12
    port map (
            O => \N__47253\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1652\
        );

    \I__10172\ : CascadeMux
    port map (
            O => \N__47250\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_0_4_cascade_\
        );

    \I__10171\ : InMux
    port map (
            O => \N__47247\,
            I => \N__47240\
        );

    \I__10170\ : InMux
    port map (
            O => \N__47246\,
            I => \N__47237\
        );

    \I__10169\ : InMux
    port map (
            O => \N__47245\,
            I => \N__47232\
        );

    \I__10168\ : InMux
    port map (
            O => \N__47244\,
            I => \N__47232\
        );

    \I__10167\ : InMux
    port map (
            O => \N__47243\,
            I => \N__47229\
        );

    \I__10166\ : LocalMux
    port map (
            O => \N__47240\,
            I => \N__47222\
        );

    \I__10165\ : LocalMux
    port map (
            O => \N__47237\,
            I => \N__47222\
        );

    \I__10164\ : LocalMux
    port map (
            O => \N__47232\,
            I => \N__47222\
        );

    \I__10163\ : LocalMux
    port map (
            O => \N__47229\,
            I => \N__47219\
        );

    \I__10162\ : Span4Mux_h
    port map (
            O => \N__47222\,
            I => \N__47216\
        );

    \I__10161\ : Span4Mux_v
    port map (
            O => \N__47219\,
            I => \N__47213\
        );

    \I__10160\ : Odrv4
    port map (
            O => \N__47216\,
            I => \s_paddr_I2C_5\
        );

    \I__10159\ : Odrv4
    port map (
            O => \N__47213\,
            I => \s_paddr_I2C_5\
        );

    \I__10158\ : InMux
    port map (
            O => \N__47208\,
            I => \N__47201\
        );

    \I__10157\ : InMux
    port map (
            O => \N__47207\,
            I => \N__47201\
        );

    \I__10156\ : InMux
    port map (
            O => \N__47206\,
            I => \N__47198\
        );

    \I__10155\ : LocalMux
    port map (
            O => \N__47201\,
            I => \N__47193\
        );

    \I__10154\ : LocalMux
    port map (
            O => \N__47198\,
            I => \N__47190\
        );

    \I__10153\ : InMux
    port map (
            O => \N__47197\,
            I => \N__47187\
        );

    \I__10152\ : InMux
    port map (
            O => \N__47196\,
            I => \N__47184\
        );

    \I__10151\ : Span4Mux_v
    port map (
            O => \N__47193\,
            I => \N__47179\
        );

    \I__10150\ : Span4Mux_v
    port map (
            O => \N__47190\,
            I => \N__47179\
        );

    \I__10149\ : LocalMux
    port map (
            O => \N__47187\,
            I => \s_paddr_I2C_4\
        );

    \I__10148\ : LocalMux
    port map (
            O => \N__47184\,
            I => \s_paddr_I2C_4\
        );

    \I__10147\ : Odrv4
    port map (
            O => \N__47179\,
            I => \s_paddr_I2C_4\
        );

    \I__10146\ : InMux
    port map (
            O => \N__47172\,
            I => \N__47165\
        );

    \I__10145\ : InMux
    port map (
            O => \N__47171\,
            I => \N__47161\
        );

    \I__10144\ : InMux
    port map (
            O => \N__47170\,
            I => \N__47158\
        );

    \I__10143\ : InMux
    port map (
            O => \N__47169\,
            I => \N__47153\
        );

    \I__10142\ : InMux
    port map (
            O => \N__47168\,
            I => \N__47153\
        );

    \I__10141\ : LocalMux
    port map (
            O => \N__47165\,
            I => \N__47150\
        );

    \I__10140\ : InMux
    port map (
            O => \N__47164\,
            I => \N__47147\
        );

    \I__10139\ : LocalMux
    port map (
            O => \N__47161\,
            I => \N__47140\
        );

    \I__10138\ : LocalMux
    port map (
            O => \N__47158\,
            I => \N__47140\
        );

    \I__10137\ : LocalMux
    port map (
            O => \N__47153\,
            I => \N__47140\
        );

    \I__10136\ : Span4Mux_v
    port map (
            O => \N__47150\,
            I => \N__47137\
        );

    \I__10135\ : LocalMux
    port map (
            O => \N__47147\,
            I => \N__47134\
        );

    \I__10134\ : Span4Mux_v
    port map (
            O => \N__47140\,
            I => \N__47129\
        );

    \I__10133\ : Span4Mux_h
    port map (
            O => \N__47137\,
            I => \N__47129\
        );

    \I__10132\ : Odrv4
    port map (
            O => \N__47134\,
            I => \s_paddr_I2C_6\
        );

    \I__10131\ : Odrv4
    port map (
            O => \N__47129\,
            I => \s_paddr_I2C_6\
        );

    \I__10130\ : CascadeMux
    port map (
            O => \N__47124\,
            I => \N__47119\
        );

    \I__10129\ : CascadeMux
    port map (
            O => \N__47123\,
            I => \N__47115\
        );

    \I__10128\ : CascadeMux
    port map (
            O => \N__47122\,
            I => \N__47112\
        );

    \I__10127\ : InMux
    port map (
            O => \N__47119\,
            I => \N__47107\
        );

    \I__10126\ : InMux
    port map (
            O => \N__47118\,
            I => \N__47104\
        );

    \I__10125\ : InMux
    port map (
            O => \N__47115\,
            I => \N__47099\
        );

    \I__10124\ : InMux
    port map (
            O => \N__47112\,
            I => \N__47099\
        );

    \I__10123\ : InMux
    port map (
            O => \N__47111\,
            I => \N__47094\
        );

    \I__10122\ : InMux
    port map (
            O => \N__47110\,
            I => \N__47094\
        );

    \I__10121\ : LocalMux
    port map (
            O => \N__47107\,
            I => \N__47090\
        );

    \I__10120\ : LocalMux
    port map (
            O => \N__47104\,
            I => \N__47085\
        );

    \I__10119\ : LocalMux
    port map (
            O => \N__47099\,
            I => \N__47085\
        );

    \I__10118\ : LocalMux
    port map (
            O => \N__47094\,
            I => \N__47082\
        );

    \I__10117\ : InMux
    port map (
            O => \N__47093\,
            I => \N__47079\
        );

    \I__10116\ : Span4Mux_h
    port map (
            O => \N__47090\,
            I => \N__47076\
        );

    \I__10115\ : Span4Mux_h
    port map (
            O => \N__47085\,
            I => \N__47073\
        );

    \I__10114\ : Span4Mux_h
    port map (
            O => \N__47082\,
            I => \N__47068\
        );

    \I__10113\ : LocalMux
    port map (
            O => \N__47079\,
            I => \N__47068\
        );

    \I__10112\ : Odrv4
    port map (
            O => \N__47076\,
            I => \s_paddr_I2C_7\
        );

    \I__10111\ : Odrv4
    port map (
            O => \N__47073\,
            I => \s_paddr_I2C_7\
        );

    \I__10110\ : Odrv4
    port map (
            O => \N__47068\,
            I => \s_paddr_I2C_7\
        );

    \I__10109\ : InMux
    port map (
            O => \N__47061\,
            I => \N__47058\
        );

    \I__10108\ : LocalMux
    port map (
            O => \N__47058\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_2\
        );

    \I__10107\ : InMux
    port map (
            O => \N__47055\,
            I => \N__47052\
        );

    \I__10106\ : LocalMux
    port map (
            O => \N__47052\,
            I => \N__47049\
        );

    \I__10105\ : Span4Mux_v
    port map (
            O => \N__47049\,
            I => \N__47046\
        );

    \I__10104\ : Odrv4
    port map (
            O => \N__47046\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_5\
        );

    \I__10103\ : InMux
    port map (
            O => \N__47043\,
            I => \N__47038\
        );

    \I__10102\ : InMux
    port map (
            O => \N__47042\,
            I => \N__47034\
        );

    \I__10101\ : InMux
    port map (
            O => \N__47041\,
            I => \N__47031\
        );

    \I__10100\ : LocalMux
    port map (
            O => \N__47038\,
            I => \N__47028\
        );

    \I__10099\ : InMux
    port map (
            O => \N__47037\,
            I => \N__47025\
        );

    \I__10098\ : LocalMux
    port map (
            O => \N__47034\,
            I => \N__47018\
        );

    \I__10097\ : LocalMux
    port map (
            O => \N__47031\,
            I => \N__47018\
        );

    \I__10096\ : Span4Mux_v
    port map (
            O => \N__47028\,
            I => \N__47018\
        );

    \I__10095\ : LocalMux
    port map (
            O => \N__47025\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10\
        );

    \I__10094\ : Odrv4
    port map (
            O => \N__47018\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10\
        );

    \I__10093\ : InMux
    port map (
            O => \N__47013\,
            I => \N__47009\
        );

    \I__10092\ : InMux
    port map (
            O => \N__47012\,
            I => \N__47004\
        );

    \I__10091\ : LocalMux
    port map (
            O => \N__47009\,
            I => \N__47001\
        );

    \I__10090\ : InMux
    port map (
            O => \N__47008\,
            I => \N__46998\
        );

    \I__10089\ : InMux
    port map (
            O => \N__47007\,
            I => \N__46995\
        );

    \I__10088\ : LocalMux
    port map (
            O => \N__47004\,
            I => \N__46992\
        );

    \I__10087\ : Span4Mux_h
    port map (
            O => \N__47001\,
            I => \N__46989\
        );

    \I__10086\ : LocalMux
    port map (
            O => \N__46998\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9\
        );

    \I__10085\ : LocalMux
    port map (
            O => \N__46995\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9\
        );

    \I__10084\ : Odrv4
    port map (
            O => \N__46992\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9\
        );

    \I__10083\ : Odrv4
    port map (
            O => \N__46989\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9\
        );

    \I__10082\ : InMux
    port map (
            O => \N__46980\,
            I => \N__46977\
        );

    \I__10081\ : LocalMux
    port map (
            O => \N__46977\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_3\
        );

    \I__10080\ : InMux
    port map (
            O => \N__46974\,
            I => \N__46971\
        );

    \I__10079\ : LocalMux
    port map (
            O => \N__46971\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_2_2\
        );

    \I__10078\ : CascadeMux
    port map (
            O => \N__46968\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0_cascade_\
        );

    \I__10077\ : CascadeMux
    port map (
            O => \N__46965\,
            I => \N__46962\
        );

    \I__10076\ : InMux
    port map (
            O => \N__46962\,
            I => \N__46959\
        );

    \I__10075\ : LocalMux
    port map (
            O => \N__46959\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0\
        );

    \I__10074\ : InMux
    port map (
            O => \N__46956\,
            I => \N__46953\
        );

    \I__10073\ : LocalMux
    port map (
            O => \N__46953\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_1_0\
        );

    \I__10072\ : CascadeMux
    port map (
            O => \N__46950\,
            I => \N__46947\
        );

    \I__10071\ : InMux
    port map (
            O => \N__46947\,
            I => \N__46943\
        );

    \I__10070\ : InMux
    port map (
            O => \N__46946\,
            I => \N__46939\
        );

    \I__10069\ : LocalMux
    port map (
            O => \N__46943\,
            I => \N__46935\
        );

    \I__10068\ : InMux
    port map (
            O => \N__46942\,
            I => \N__46932\
        );

    \I__10067\ : LocalMux
    port map (
            O => \N__46939\,
            I => \N__46929\
        );

    \I__10066\ : InMux
    port map (
            O => \N__46938\,
            I => \N__46926\
        );

    \I__10065\ : Span4Mux_h
    port map (
            O => \N__46935\,
            I => \N__46923\
        );

    \I__10064\ : LocalMux
    port map (
            O => \N__46932\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11\
        );

    \I__10063\ : Odrv4
    port map (
            O => \N__46929\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11\
        );

    \I__10062\ : LocalMux
    port map (
            O => \N__46926\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11\
        );

    \I__10061\ : Odrv4
    port map (
            O => \N__46923\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11\
        );

    \I__10060\ : CascadeMux
    port map (
            O => \N__46914\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0_cascade_\
        );

    \I__10059\ : InMux
    port map (
            O => \N__46911\,
            I => \N__46904\
        );

    \I__10058\ : CascadeMux
    port map (
            O => \N__46910\,
            I => \N__46901\
        );

    \I__10057\ : CascadeMux
    port map (
            O => \N__46909\,
            I => \N__46897\
        );

    \I__10056\ : CascadeMux
    port map (
            O => \N__46908\,
            I => \N__46893\
        );

    \I__10055\ : InMux
    port map (
            O => \N__46907\,
            I => \N__46888\
        );

    \I__10054\ : LocalMux
    port map (
            O => \N__46904\,
            I => \N__46885\
        );

    \I__10053\ : InMux
    port map (
            O => \N__46901\,
            I => \N__46876\
        );

    \I__10052\ : InMux
    port map (
            O => \N__46900\,
            I => \N__46876\
        );

    \I__10051\ : InMux
    port map (
            O => \N__46897\,
            I => \N__46876\
        );

    \I__10050\ : InMux
    port map (
            O => \N__46896\,
            I => \N__46876\
        );

    \I__10049\ : InMux
    port map (
            O => \N__46893\,
            I => \N__46869\
        );

    \I__10048\ : InMux
    port map (
            O => \N__46892\,
            I => \N__46869\
        );

    \I__10047\ : InMux
    port map (
            O => \N__46891\,
            I => \N__46869\
        );

    \I__10046\ : LocalMux
    port map (
            O => \N__46888\,
            I => \N__46866\
        );

    \I__10045\ : Span4Mux_v
    port map (
            O => \N__46885\,
            I => \N__46863\
        );

    \I__10044\ : LocalMux
    port map (
            O => \N__46876\,
            I => \N__46860\
        );

    \I__10043\ : LocalMux
    port map (
            O => \N__46869\,
            I => \N__46857\
        );

    \I__10042\ : Span4Mux_v
    port map (
            O => \N__46866\,
            I => \N__46854\
        );

    \I__10041\ : Span4Mux_h
    port map (
            O => \N__46863\,
            I => \N__46849\
        );

    \I__10040\ : Span4Mux_v
    port map (
            O => \N__46860\,
            I => \N__46849\
        );

    \I__10039\ : Span4Mux_h
    port map (
            O => \N__46857\,
            I => \N__46846\
        );

    \I__10038\ : Sp12to4
    port map (
            O => \N__46854\,
            I => \N__46843\
        );

    \I__10037\ : Sp12to4
    port map (
            O => \N__46849\,
            I => \N__46840\
        );

    \I__10036\ : Span4Mux_v
    port map (
            O => \N__46846\,
            I => \N__46837\
        );

    \I__10035\ : Span12Mux_h
    port map (
            O => \N__46843\,
            I => \N__46832\
        );

    \I__10034\ : Span12Mux_h
    port map (
            O => \N__46840\,
            I => \N__46832\
        );

    \I__10033\ : Span4Mux_v
    port map (
            O => \N__46837\,
            I => \N__46829\
        );

    \I__10032\ : Odrv12
    port map (
            O => \N__46832\,
            I => \s_paddr_I2C_2\
        );

    \I__10031\ : Odrv4
    port map (
            O => \N__46829\,
            I => \s_paddr_I2C_2\
        );

    \I__10030\ : InMux
    port map (
            O => \N__46824\,
            I => \N__46821\
        );

    \I__10029\ : LocalMux
    port map (
            O => \N__46821\,
            I => \N__46818\
        );

    \I__10028\ : Span4Mux_v
    port map (
            O => \N__46818\,
            I => \N__46814\
        );

    \I__10027\ : InMux
    port map (
            O => \N__46817\,
            I => \N__46808\
        );

    \I__10026\ : Span4Mux_h
    port map (
            O => \N__46814\,
            I => \N__46804\
        );

    \I__10025\ : InMux
    port map (
            O => \N__46813\,
            I => \N__46799\
        );

    \I__10024\ : InMux
    port map (
            O => \N__46812\,
            I => \N__46799\
        );

    \I__10023\ : InMux
    port map (
            O => \N__46811\,
            I => \N__46796\
        );

    \I__10022\ : LocalMux
    port map (
            O => \N__46808\,
            I => \N__46793\
        );

    \I__10021\ : InMux
    port map (
            O => \N__46807\,
            I => \N__46790\
        );

    \I__10020\ : Sp12to4
    port map (
            O => \N__46804\,
            I => \N__46787\
        );

    \I__10019\ : LocalMux
    port map (
            O => \N__46799\,
            I => \N__46782\
        );

    \I__10018\ : LocalMux
    port map (
            O => \N__46796\,
            I => \N__46782\
        );

    \I__10017\ : Span4Mux_v
    port map (
            O => \N__46793\,
            I => \N__46779\
        );

    \I__10016\ : LocalMux
    port map (
            O => \N__46790\,
            I => \N__46772\
        );

    \I__10015\ : Span12Mux_v
    port map (
            O => \N__46787\,
            I => \N__46772\
        );

    \I__10014\ : Span12Mux_h
    port map (
            O => \N__46782\,
            I => \N__46772\
        );

    \I__10013\ : Span4Mux_v
    port map (
            O => \N__46779\,
            I => \N__46769\
        );

    \I__10012\ : Odrv12
    port map (
            O => \N__46772\,
            I => \s_paddr_I2C_1\
        );

    \I__10011\ : Odrv4
    port map (
            O => \N__46769\,
            I => \s_paddr_I2C_1\
        );

    \I__10010\ : InMux
    port map (
            O => \N__46764\,
            I => \N__46757\
        );

    \I__10009\ : CascadeMux
    port map (
            O => \N__46763\,
            I => \N__46753\
        );

    \I__10008\ : InMux
    port map (
            O => \N__46762\,
            I => \N__46746\
        );

    \I__10007\ : InMux
    port map (
            O => \N__46761\,
            I => \N__46746\
        );

    \I__10006\ : InMux
    port map (
            O => \N__46760\,
            I => \N__46746\
        );

    \I__10005\ : LocalMux
    port map (
            O => \N__46757\,
            I => \N__46743\
        );

    \I__10004\ : InMux
    port map (
            O => \N__46756\,
            I => \N__46740\
        );

    \I__10003\ : InMux
    port map (
            O => \N__46753\,
            I => \N__46737\
        );

    \I__10002\ : LocalMux
    port map (
            O => \N__46746\,
            I => \N__46732\
        );

    \I__10001\ : Span4Mux_v
    port map (
            O => \N__46743\,
            I => \N__46732\
        );

    \I__10000\ : LocalMux
    port map (
            O => \N__46740\,
            I => \s_paddr_I2C_0\
        );

    \I__9999\ : LocalMux
    port map (
            O => \N__46737\,
            I => \s_paddr_I2C_0\
        );

    \I__9998\ : Odrv4
    port map (
            O => \N__46732\,
            I => \s_paddr_I2C_0\
        );

    \I__9997\ : InMux
    port map (
            O => \N__46725\,
            I => \N__46722\
        );

    \I__9996\ : LocalMux
    port map (
            O => \N__46722\,
            I => \N__46719\
        );

    \I__9995\ : Span4Mux_v
    port map (
            O => \N__46719\,
            I => \N__46716\
        );

    \I__9994\ : Span4Mux_h
    port map (
            O => \N__46716\,
            I => \N__46713\
        );

    \I__9993\ : Odrv4
    port map (
            O => \N__46713\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_10\
        );

    \I__9992\ : InMux
    port map (
            O => \N__46710\,
            I => \N__46707\
        );

    \I__9991\ : LocalMux
    port map (
            O => \N__46707\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_10\
        );

    \I__9990\ : CascadeMux
    port map (
            O => \N__46704\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7DZ0Z7_cascade_\
        );

    \I__9989\ : InMux
    port map (
            O => \N__46701\,
            I => \N__46698\
        );

    \I__9988\ : LocalMux
    port map (
            O => \N__46698\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10\
        );

    \I__9987\ : InMux
    port map (
            O => \N__46695\,
            I => \N__46692\
        );

    \I__9986\ : LocalMux
    port map (
            O => \N__46692\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_9\
        );

    \I__9985\ : CascadeMux
    port map (
            O => \N__46689\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10_cascade_\
        );

    \I__9984\ : InMux
    port map (
            O => \N__46686\,
            I => \N__46683\
        );

    \I__9983\ : LocalMux
    port map (
            O => \N__46683\,
            I => \N__46680\
        );

    \I__9982\ : Span4Mux_h
    port map (
            O => \N__46680\,
            I => \N__46677\
        );

    \I__9981\ : Span4Mux_v
    port map (
            O => \N__46677\,
            I => \N__46674\
        );

    \I__9980\ : Odrv4
    port map (
            O => \N__46674\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_10\
        );

    \I__9979\ : InMux
    port map (
            O => \N__46671\,
            I => \N__46668\
        );

    \I__9978\ : LocalMux
    port map (
            O => \N__46668\,
            I => \N__46664\
        );

    \I__9977\ : CascadeMux
    port map (
            O => \N__46667\,
            I => \N__46661\
        );

    \I__9976\ : Span4Mux_v
    port map (
            O => \N__46664\,
            I => \N__46657\
        );

    \I__9975\ : InMux
    port map (
            O => \N__46661\,
            I => \N__46654\
        );

    \I__9974\ : InMux
    port map (
            O => \N__46660\,
            I => \N__46651\
        );

    \I__9973\ : Span4Mux_h
    port map (
            O => \N__46657\,
            I => \N__46644\
        );

    \I__9972\ : LocalMux
    port map (
            O => \N__46654\,
            I => \N__46644\
        );

    \I__9971\ : LocalMux
    port map (
            O => \N__46651\,
            I => \N__46644\
        );

    \I__9970\ : Odrv4
    port map (
            O => \N__46644\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_9
        );

    \I__9969\ : InMux
    port map (
            O => \N__46641\,
            I => \N__46638\
        );

    \I__9968\ : LocalMux
    port map (
            O => \N__46638\,
            I => \N__46635\
        );

    \I__9967\ : Span4Mux_h
    port map (
            O => \N__46635\,
            I => \N__46631\
        );

    \I__9966\ : CascadeMux
    port map (
            O => \N__46634\,
            I => \N__46628\
        );

    \I__9965\ : Span4Mux_h
    port map (
            O => \N__46631\,
            I => \N__46624\
        );

    \I__9964\ : InMux
    port map (
            O => \N__46628\,
            I => \N__46619\
        );

    \I__9963\ : InMux
    port map (
            O => \N__46627\,
            I => \N__46619\
        );

    \I__9962\ : Odrv4
    port map (
            O => \N__46624\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_9
        );

    \I__9961\ : LocalMux
    port map (
            O => \N__46619\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_9
        );

    \I__9960\ : InMux
    port map (
            O => \N__46614\,
            I => \N__46611\
        );

    \I__9959\ : LocalMux
    port map (
            O => \N__46611\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_9\
        );

    \I__9958\ : CascadeMux
    port map (
            O => \N__46608\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i_cascade_\
        );

    \I__9957\ : InMux
    port map (
            O => \N__46605\,
            I => \N__46602\
        );

    \I__9956\ : LocalMux
    port map (
            O => \N__46602\,
            I => \N__46599\
        );

    \I__9955\ : Sp12to4
    port map (
            O => \N__46599\,
            I => \N__46594\
        );

    \I__9954\ : InMux
    port map (
            O => \N__46598\,
            I => \N__46589\
        );

    \I__9953\ : InMux
    port map (
            O => \N__46597\,
            I => \N__46589\
        );

    \I__9952\ : Span12Mux_v
    port map (
            O => \N__46594\,
            I => \N__46586\
        );

    \I__9951\ : LocalMux
    port map (
            O => \N__46589\,
            I => \N__46583\
        );

    \I__9950\ : Odrv12
    port map (
            O => \N__46586\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_15
        );

    \I__9949\ : Odrv4
    port map (
            O => \N__46583\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_15
        );

    \I__9948\ : InMux
    port map (
            O => \N__46578\,
            I => \N__46575\
        );

    \I__9947\ : LocalMux
    port map (
            O => \N__46575\,
            I => \N__46572\
        );

    \I__9946\ : Span4Mux_v
    port map (
            O => \N__46572\,
            I => \N__46569\
        );

    \I__9945\ : Span4Mux_v
    port map (
            O => \N__46569\,
            I => \N__46566\
        );

    \I__9944\ : Odrv4
    port map (
            O => \N__46566\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_24\
        );

    \I__9943\ : InMux
    port map (
            O => \N__46563\,
            I => \N__46560\
        );

    \I__9942\ : LocalMux
    port map (
            O => \N__46560\,
            I => \N__46557\
        );

    \I__9941\ : Span4Mux_v
    port map (
            O => \N__46557\,
            I => \N__46553\
        );

    \I__9940\ : CascadeMux
    port map (
            O => \N__46556\,
            I => \N__46549\
        );

    \I__9939\ : Span4Mux_v
    port map (
            O => \N__46553\,
            I => \N__46546\
        );

    \I__9938\ : InMux
    port map (
            O => \N__46552\,
            I => \N__46541\
        );

    \I__9937\ : InMux
    port map (
            O => \N__46549\,
            I => \N__46541\
        );

    \I__9936\ : Span4Mux_h
    port map (
            O => \N__46546\,
            I => \N__46538\
        );

    \I__9935\ : LocalMux
    port map (
            O => \N__46541\,
            I => \N__46535\
        );

    \I__9934\ : Odrv4
    port map (
            O => \N__46538\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_17
        );

    \I__9933\ : Odrv12
    port map (
            O => \N__46535\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_17
        );

    \I__9932\ : InMux
    port map (
            O => \N__46530\,
            I => \N__46527\
        );

    \I__9931\ : LocalMux
    port map (
            O => \N__46527\,
            I => \N__46520\
        );

    \I__9930\ : InMux
    port map (
            O => \N__46526\,
            I => \N__46517\
        );

    \I__9929\ : InMux
    port map (
            O => \N__46525\,
            I => \N__46514\
        );

    \I__9928\ : InMux
    port map (
            O => \N__46524\,
            I => \N__46511\
        );

    \I__9927\ : InMux
    port map (
            O => \N__46523\,
            I => \N__46508\
        );

    \I__9926\ : Span4Mux_v
    port map (
            O => \N__46520\,
            I => \N__46502\
        );

    \I__9925\ : LocalMux
    port map (
            O => \N__46517\,
            I => \N__46502\
        );

    \I__9924\ : LocalMux
    port map (
            O => \N__46514\,
            I => \N__46497\
        );

    \I__9923\ : LocalMux
    port map (
            O => \N__46511\,
            I => \N__46494\
        );

    \I__9922\ : LocalMux
    port map (
            O => \N__46508\,
            I => \N__46491\
        );

    \I__9921\ : CascadeMux
    port map (
            O => \N__46507\,
            I => \N__46488\
        );

    \I__9920\ : Span4Mux_h
    port map (
            O => \N__46502\,
            I => \N__46485\
        );

    \I__9919\ : InMux
    port map (
            O => \N__46501\,
            I => \N__46482\
        );

    \I__9918\ : InMux
    port map (
            O => \N__46500\,
            I => \N__46479\
        );

    \I__9917\ : Span4Mux_v
    port map (
            O => \N__46497\,
            I => \N__46476\
        );

    \I__9916\ : Span4Mux_v
    port map (
            O => \N__46494\,
            I => \N__46471\
        );

    \I__9915\ : Span4Mux_h
    port map (
            O => \N__46491\,
            I => \N__46471\
        );

    \I__9914\ : InMux
    port map (
            O => \N__46488\,
            I => \N__46468\
        );

    \I__9913\ : Span4Mux_h
    port map (
            O => \N__46485\,
            I => \N__46465\
        );

    \I__9912\ : LocalMux
    port map (
            O => \N__46482\,
            I => \N__46462\
        );

    \I__9911\ : LocalMux
    port map (
            O => \N__46479\,
            I => \N__46458\
        );

    \I__9910\ : Span4Mux_v
    port map (
            O => \N__46476\,
            I => \N__46453\
        );

    \I__9909\ : Span4Mux_h
    port map (
            O => \N__46471\,
            I => \N__46453\
        );

    \I__9908\ : LocalMux
    port map (
            O => \N__46468\,
            I => \N__46450\
        );

    \I__9907\ : Span4Mux_h
    port map (
            O => \N__46465\,
            I => \N__46447\
        );

    \I__9906\ : Span4Mux_v
    port map (
            O => \N__46462\,
            I => \N__46444\
        );

    \I__9905\ : InMux
    port map (
            O => \N__46461\,
            I => \N__46441\
        );

    \I__9904\ : Span12Mux_v
    port map (
            O => \N__46458\,
            I => \N__46438\
        );

    \I__9903\ : Span4Mux_h
    port map (
            O => \N__46453\,
            I => \N__46435\
        );

    \I__9902\ : Span4Mux_h
    port map (
            O => \N__46450\,
            I => \N__46428\
        );

    \I__9901\ : Span4Mux_h
    port map (
            O => \N__46447\,
            I => \N__46428\
        );

    \I__9900\ : Span4Mux_h
    port map (
            O => \N__46444\,
            I => \N__46428\
        );

    \I__9899\ : LocalMux
    port map (
            O => \N__46441\,
            I => \I2C_top_level_inst1_s_data_oreg_9\
        );

    \I__9898\ : Odrv12
    port map (
            O => \N__46438\,
            I => \I2C_top_level_inst1_s_data_oreg_9\
        );

    \I__9897\ : Odrv4
    port map (
            O => \N__46435\,
            I => \I2C_top_level_inst1_s_data_oreg_9\
        );

    \I__9896\ : Odrv4
    port map (
            O => \N__46428\,
            I => \I2C_top_level_inst1_s_data_oreg_9\
        );

    \I__9895\ : CascadeMux
    port map (
            O => \N__46419\,
            I => \N__46416\
        );

    \I__9894\ : InMux
    port map (
            O => \N__46416\,
            I => \N__46413\
        );

    \I__9893\ : LocalMux
    port map (
            O => \N__46413\,
            I => \N__46410\
        );

    \I__9892\ : Span4Mux_v
    port map (
            O => \N__46410\,
            I => \N__46407\
        );

    \I__9891\ : Odrv4
    port map (
            O => \N__46407\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_9\
        );

    \I__9890\ : CascadeMux
    port map (
            O => \N__46404\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSLZ0Z7_cascade_\
        );

    \I__9889\ : InMux
    port map (
            O => \N__46401\,
            I => \N__46398\
        );

    \I__9888\ : LocalMux
    port map (
            O => \N__46398\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9\
        );

    \I__9887\ : CascadeMux
    port map (
            O => \N__46395\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9_cascade_\
        );

    \I__9886\ : InMux
    port map (
            O => \N__46392\,
            I => \N__46389\
        );

    \I__9885\ : LocalMux
    port map (
            O => \N__46389\,
            I => \N__46386\
        );

    \I__9884\ : Span4Mux_h
    port map (
            O => \N__46386\,
            I => \N__46383\
        );

    \I__9883\ : Odrv4
    port map (
            O => \N__46383\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_8\
        );

    \I__9882\ : InMux
    port map (
            O => \N__46380\,
            I => \N__46377\
        );

    \I__9881\ : LocalMux
    port map (
            O => \N__46377\,
            I => \N__46373\
        );

    \I__9880\ : InMux
    port map (
            O => \N__46376\,
            I => \N__46370\
        );

    \I__9879\ : Span4Mux_v
    port map (
            O => \N__46373\,
            I => \N__46366\
        );

    \I__9878\ : LocalMux
    port map (
            O => \N__46370\,
            I => \N__46363\
        );

    \I__9877\ : InMux
    port map (
            O => \N__46369\,
            I => \N__46360\
        );

    \I__9876\ : Span4Mux_h
    port map (
            O => \N__46366\,
            I => \N__46355\
        );

    \I__9875\ : Span4Mux_v
    port map (
            O => \N__46363\,
            I => \N__46355\
        );

    \I__9874\ : LocalMux
    port map (
            O => \N__46360\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_11
        );

    \I__9873\ : Odrv4
    port map (
            O => \N__46355\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_11
        );

    \I__9872\ : InMux
    port map (
            O => \N__46350\,
            I => \N__46347\
        );

    \I__9871\ : LocalMux
    port map (
            O => \N__46347\,
            I => \N__46343\
        );

    \I__9870\ : InMux
    port map (
            O => \N__46346\,
            I => \N__46340\
        );

    \I__9869\ : Span4Mux_v
    port map (
            O => \N__46343\,
            I => \N__46336\
        );

    \I__9868\ : LocalMux
    port map (
            O => \N__46340\,
            I => \N__46333\
        );

    \I__9867\ : InMux
    port map (
            O => \N__46339\,
            I => \N__46330\
        );

    \I__9866\ : Span4Mux_h
    port map (
            O => \N__46336\,
            I => \N__46327\
        );

    \I__9865\ : Span4Mux_v
    port map (
            O => \N__46333\,
            I => \N__46322\
        );

    \I__9864\ : LocalMux
    port map (
            O => \N__46330\,
            I => \N__46322\
        );

    \I__9863\ : Odrv4
    port map (
            O => \N__46327\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_12
        );

    \I__9862\ : Odrv4
    port map (
            O => \N__46322\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_12
        );

    \I__9861\ : InMux
    port map (
            O => \N__46317\,
            I => \N__46314\
        );

    \I__9860\ : LocalMux
    port map (
            O => \N__46314\,
            I => \N__46311\
        );

    \I__9859\ : Span4Mux_h
    port map (
            O => \N__46311\,
            I => \N__46308\
        );

    \I__9858\ : Span4Mux_h
    port map (
            O => \N__46308\,
            I => \N__46303\
        );

    \I__9857\ : InMux
    port map (
            O => \N__46307\,
            I => \N__46298\
        );

    \I__9856\ : InMux
    port map (
            O => \N__46306\,
            I => \N__46298\
        );

    \I__9855\ : Odrv4
    port map (
            O => \N__46303\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_21
        );

    \I__9854\ : LocalMux
    port map (
            O => \N__46298\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_21
        );

    \I__9853\ : CascadeMux
    port map (
            O => \N__46293\,
            I => \N__46290\
        );

    \I__9852\ : InMux
    port map (
            O => \N__46290\,
            I => \N__46287\
        );

    \I__9851\ : LocalMux
    port map (
            O => \N__46287\,
            I => \N__46284\
        );

    \I__9850\ : Span4Mux_h
    port map (
            O => \N__46284\,
            I => \N__46281\
        );

    \I__9849\ : Span4Mux_h
    port map (
            O => \N__46281\,
            I => \N__46278\
        );

    \I__9848\ : Span4Mux_h
    port map (
            O => \N__46278\,
            I => \N__46275\
        );

    \I__9847\ : Odrv4
    port map (
            O => \N__46275\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_30\
        );

    \I__9846\ : InMux
    port map (
            O => \N__46272\,
            I => \N__46267\
        );

    \I__9845\ : InMux
    port map (
            O => \N__46271\,
            I => \N__46264\
        );

    \I__9844\ : InMux
    port map (
            O => \N__46270\,
            I => \N__46261\
        );

    \I__9843\ : LocalMux
    port map (
            O => \N__46267\,
            I => \N__46258\
        );

    \I__9842\ : LocalMux
    port map (
            O => \N__46264\,
            I => \N__46255\
        );

    \I__9841\ : LocalMux
    port map (
            O => \N__46261\,
            I => \N__46252\
        );

    \I__9840\ : Span4Mux_v
    port map (
            O => \N__46258\,
            I => \N__46249\
        );

    \I__9839\ : Span4Mux_h
    port map (
            O => \N__46255\,
            I => \N__46246\
        );

    \I__9838\ : Span4Mux_h
    port map (
            O => \N__46252\,
            I => \N__46243\
        );

    \I__9837\ : Span4Mux_h
    port map (
            O => \N__46249\,
            I => \N__46240\
        );

    \I__9836\ : Span4Mux_h
    port map (
            O => \N__46246\,
            I => \N__46237\
        );

    \I__9835\ : Span4Mux_h
    port map (
            O => \N__46243\,
            I => \N__46234\
        );

    \I__9834\ : Odrv4
    port map (
            O => \N__46240\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_13
        );

    \I__9833\ : Odrv4
    port map (
            O => \N__46237\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_13
        );

    \I__9832\ : Odrv4
    port map (
            O => \N__46234\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_13
        );

    \I__9831\ : CascadeMux
    port map (
            O => \N__46227\,
            I => \N__46224\
        );

    \I__9830\ : InMux
    port map (
            O => \N__46224\,
            I => \N__46221\
        );

    \I__9829\ : LocalMux
    port map (
            O => \N__46221\,
            I => \N__46218\
        );

    \I__9828\ : Span12Mux_v
    port map (
            O => \N__46218\,
            I => \N__46215\
        );

    \I__9827\ : Odrv12
    port map (
            O => \N__46215\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_31\
        );

    \I__9826\ : InMux
    port map (
            O => \N__46212\,
            I => \N__46208\
        );

    \I__9825\ : InMux
    port map (
            O => \N__46211\,
            I => \N__46205\
        );

    \I__9824\ : LocalMux
    port map (
            O => \N__46208\,
            I => \N__46202\
        );

    \I__9823\ : LocalMux
    port map (
            O => \N__46205\,
            I => \N__46199\
        );

    \I__9822\ : Span4Mux_h
    port map (
            O => \N__46202\,
            I => \N__46195\
        );

    \I__9821\ : Span4Mux_h
    port map (
            O => \N__46199\,
            I => \N__46192\
        );

    \I__9820\ : InMux
    port map (
            O => \N__46198\,
            I => \N__46189\
        );

    \I__9819\ : Span4Mux_h
    port map (
            O => \N__46195\,
            I => \N__46186\
        );

    \I__9818\ : Span4Mux_h
    port map (
            O => \N__46192\,
            I => \N__46183\
        );

    \I__9817\ : LocalMux
    port map (
            O => \N__46189\,
            I => \N__46180\
        );

    \I__9816\ : Odrv4
    port map (
            O => \N__46186\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_15
        );

    \I__9815\ : Odrv4
    port map (
            O => \N__46183\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_15
        );

    \I__9814\ : Odrv12
    port map (
            O => \N__46180\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_15
        );

    \I__9813\ : InMux
    port map (
            O => \N__46173\,
            I => \N__46169\
        );

    \I__9812\ : CascadeMux
    port map (
            O => \N__46172\,
            I => \N__46166\
        );

    \I__9811\ : LocalMux
    port map (
            O => \N__46169\,
            I => \N__46163\
        );

    \I__9810\ : InMux
    port map (
            O => \N__46166\,
            I => \N__46160\
        );

    \I__9809\ : Span4Mux_v
    port map (
            O => \N__46163\,
            I => \N__46154\
        );

    \I__9808\ : LocalMux
    port map (
            O => \N__46160\,
            I => \N__46154\
        );

    \I__9807\ : CascadeMux
    port map (
            O => \N__46159\,
            I => \N__46151\
        );

    \I__9806\ : Span4Mux_v
    port map (
            O => \N__46154\,
            I => \N__46148\
        );

    \I__9805\ : InMux
    port map (
            O => \N__46151\,
            I => \N__46145\
        );

    \I__9804\ : Span4Mux_h
    port map (
            O => \N__46148\,
            I => \N__46142\
        );

    \I__9803\ : LocalMux
    port map (
            O => \N__46145\,
            I => \N__46137\
        );

    \I__9802\ : Span4Mux_h
    port map (
            O => \N__46142\,
            I => \N__46137\
        );

    \I__9801\ : Odrv4
    port map (
            O => \N__46137\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_13
        );

    \I__9800\ : InMux
    port map (
            O => \N__46134\,
            I => \N__46131\
        );

    \I__9799\ : LocalMux
    port map (
            O => \N__46131\,
            I => \N__46128\
        );

    \I__9798\ : Span4Mux_h
    port map (
            O => \N__46128\,
            I => \N__46125\
        );

    \I__9797\ : Span4Mux_h
    port map (
            O => \N__46125\,
            I => \N__46122\
        );

    \I__9796\ : Span4Mux_h
    port map (
            O => \N__46122\,
            I => \N__46119\
        );

    \I__9795\ : Odrv4
    port map (
            O => \N__46119\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_31\
        );

    \I__9794\ : InMux
    port map (
            O => \N__46116\,
            I => \N__46112\
        );

    \I__9793\ : InMux
    port map (
            O => \N__46115\,
            I => \N__46109\
        );

    \I__9792\ : LocalMux
    port map (
            O => \N__46112\,
            I => \N__46106\
        );

    \I__9791\ : LocalMux
    port map (
            O => \N__46109\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11\
        );

    \I__9790\ : Odrv4
    port map (
            O => \N__46106\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11\
        );

    \I__9789\ : InMux
    port map (
            O => \N__46101\,
            I => \N__46098\
        );

    \I__9788\ : LocalMux
    port map (
            O => \N__46098\,
            I => \N__46095\
        );

    \I__9787\ : Span4Mux_h
    port map (
            O => \N__46095\,
            I => \N__46092\
        );

    \I__9786\ : Odrv4
    port map (
            O => \N__46092\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_11\
        );

    \I__9785\ : CascadeMux
    port map (
            O => \N__46089\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_21_cascade_\
        );

    \I__9784\ : InMux
    port map (
            O => \N__46086\,
            I => \N__46083\
        );

    \I__9783\ : LocalMux
    port map (
            O => \N__46083\,
            I => \N__46080\
        );

    \I__9782\ : Span4Mux_h
    port map (
            O => \N__46080\,
            I => \N__46077\
        );

    \I__9781\ : Odrv4
    port map (
            O => \N__46077\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LHZ0Z5\
        );

    \I__9780\ : InMux
    port map (
            O => \N__46074\,
            I => \N__46071\
        );

    \I__9779\ : LocalMux
    port map (
            O => \N__46071\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_21\
        );

    \I__9778\ : CascadeMux
    port map (
            O => \N__46068\,
            I => \N__46065\
        );

    \I__9777\ : InMux
    port map (
            O => \N__46065\,
            I => \N__46061\
        );

    \I__9776\ : InMux
    port map (
            O => \N__46064\,
            I => \N__46047\
        );

    \I__9775\ : LocalMux
    port map (
            O => \N__46061\,
            I => \N__46038\
        );

    \I__9774\ : InMux
    port map (
            O => \N__46060\,
            I => \N__46035\
        );

    \I__9773\ : InMux
    port map (
            O => \N__46059\,
            I => \N__46032\
        );

    \I__9772\ : InMux
    port map (
            O => \N__46058\,
            I => \N__46027\
        );

    \I__9771\ : InMux
    port map (
            O => \N__46057\,
            I => \N__46027\
        );

    \I__9770\ : InMux
    port map (
            O => \N__46056\,
            I => \N__46014\
        );

    \I__9769\ : InMux
    port map (
            O => \N__46055\,
            I => \N__46014\
        );

    \I__9768\ : InMux
    port map (
            O => \N__46054\,
            I => \N__46014\
        );

    \I__9767\ : InMux
    port map (
            O => \N__46053\,
            I => \N__46014\
        );

    \I__9766\ : InMux
    port map (
            O => \N__46052\,
            I => \N__46014\
        );

    \I__9765\ : InMux
    port map (
            O => \N__46051\,
            I => \N__46014\
        );

    \I__9764\ : InMux
    port map (
            O => \N__46050\,
            I => \N__46010\
        );

    \I__9763\ : LocalMux
    port map (
            O => \N__46047\,
            I => \N__46007\
        );

    \I__9762\ : InMux
    port map (
            O => \N__46046\,
            I => \N__45996\
        );

    \I__9761\ : InMux
    port map (
            O => \N__46045\,
            I => \N__45996\
        );

    \I__9760\ : InMux
    port map (
            O => \N__46044\,
            I => \N__45996\
        );

    \I__9759\ : InMux
    port map (
            O => \N__46043\,
            I => \N__45996\
        );

    \I__9758\ : InMux
    port map (
            O => \N__46042\,
            I => \N__45996\
        );

    \I__9757\ : CascadeMux
    port map (
            O => \N__46041\,
            I => \N__45993\
        );

    \I__9756\ : Span4Mux_h
    port map (
            O => \N__46038\,
            I => \N__45984\
        );

    \I__9755\ : LocalMux
    port map (
            O => \N__46035\,
            I => \N__45984\
        );

    \I__9754\ : LocalMux
    port map (
            O => \N__46032\,
            I => \N__45977\
        );

    \I__9753\ : LocalMux
    port map (
            O => \N__46027\,
            I => \N__45977\
        );

    \I__9752\ : LocalMux
    port map (
            O => \N__46014\,
            I => \N__45977\
        );

    \I__9751\ : InMux
    port map (
            O => \N__46013\,
            I => \N__45974\
        );

    \I__9750\ : LocalMux
    port map (
            O => \N__46010\,
            I => \N__45967\
        );

    \I__9749\ : Span4Mux_v
    port map (
            O => \N__46007\,
            I => \N__45967\
        );

    \I__9748\ : LocalMux
    port map (
            O => \N__45996\,
            I => \N__45967\
        );

    \I__9747\ : InMux
    port map (
            O => \N__45993\,
            I => \N__45962\
        );

    \I__9746\ : InMux
    port map (
            O => \N__45992\,
            I => \N__45962\
        );

    \I__9745\ : InMux
    port map (
            O => \N__45991\,
            I => \N__45959\
        );

    \I__9744\ : InMux
    port map (
            O => \N__45990\,
            I => \N__45954\
        );

    \I__9743\ : InMux
    port map (
            O => \N__45989\,
            I => \N__45954\
        );

    \I__9742\ : Span4Mux_h
    port map (
            O => \N__45984\,
            I => \N__45949\
        );

    \I__9741\ : Span4Mux_v
    port map (
            O => \N__45977\,
            I => \N__45949\
        );

    \I__9740\ : LocalMux
    port map (
            O => \N__45974\,
            I => \N__45944\
        );

    \I__9739\ : Span4Mux_h
    port map (
            O => \N__45967\,
            I => \N__45944\
        );

    \I__9738\ : LocalMux
    port map (
            O => \N__45962\,
            I => \N__45941\
        );

    \I__9737\ : LocalMux
    port map (
            O => \N__45959\,
            I => \N__45934\
        );

    \I__9736\ : LocalMux
    port map (
            O => \N__45954\,
            I => \N__45934\
        );

    \I__9735\ : Span4Mux_h
    port map (
            O => \N__45949\,
            I => \N__45934\
        );

    \I__9734\ : Span4Mux_h
    port map (
            O => \N__45944\,
            I => \N__45931\
        );

    \I__9733\ : Span4Mux_v
    port map (
            O => \N__45941\,
            I => \N__45926\
        );

    \I__9732\ : Span4Mux_h
    port map (
            O => \N__45934\,
            I => \N__45926\
        );

    \I__9731\ : Odrv4
    port map (
            O => \N__45931\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0\
        );

    \I__9730\ : Odrv4
    port map (
            O => \N__45926\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0\
        );

    \I__9729\ : CascadeMux
    port map (
            O => \N__45921\,
            I => \N__45916\
        );

    \I__9728\ : CascadeMux
    port map (
            O => \N__45920\,
            I => \N__45912\
        );

    \I__9727\ : CascadeMux
    port map (
            O => \N__45919\,
            I => \N__45909\
        );

    \I__9726\ : InMux
    port map (
            O => \N__45916\,
            I => \N__45899\
        );

    \I__9725\ : CascadeMux
    port map (
            O => \N__45915\,
            I => \N__45896\
        );

    \I__9724\ : InMux
    port map (
            O => \N__45912\,
            I => \N__45879\
        );

    \I__9723\ : InMux
    port map (
            O => \N__45909\,
            I => \N__45879\
        );

    \I__9722\ : InMux
    port map (
            O => \N__45908\,
            I => \N__45879\
        );

    \I__9721\ : InMux
    port map (
            O => \N__45907\,
            I => \N__45879\
        );

    \I__9720\ : InMux
    port map (
            O => \N__45906\,
            I => \N__45879\
        );

    \I__9719\ : InMux
    port map (
            O => \N__45905\,
            I => \N__45879\
        );

    \I__9718\ : InMux
    port map (
            O => \N__45904\,
            I => \N__45879\
        );

    \I__9717\ : InMux
    port map (
            O => \N__45903\,
            I => \N__45879\
        );

    \I__9716\ : InMux
    port map (
            O => \N__45902\,
            I => \N__45876\
        );

    \I__9715\ : LocalMux
    port map (
            O => \N__45899\,
            I => \N__45863\
        );

    \I__9714\ : InMux
    port map (
            O => \N__45896\,
            I => \N__45860\
        );

    \I__9713\ : LocalMux
    port map (
            O => \N__45879\,
            I => \N__45857\
        );

    \I__9712\ : LocalMux
    port map (
            O => \N__45876\,
            I => \N__45854\
        );

    \I__9711\ : InMux
    port map (
            O => \N__45875\,
            I => \N__45843\
        );

    \I__9710\ : InMux
    port map (
            O => \N__45874\,
            I => \N__45843\
        );

    \I__9709\ : InMux
    port map (
            O => \N__45873\,
            I => \N__45843\
        );

    \I__9708\ : InMux
    port map (
            O => \N__45872\,
            I => \N__45843\
        );

    \I__9707\ : InMux
    port map (
            O => \N__45871\,
            I => \N__45843\
        );

    \I__9706\ : CascadeMux
    port map (
            O => \N__45870\,
            I => \N__45839\
        );

    \I__9705\ : InMux
    port map (
            O => \N__45869\,
            I => \N__45836\
        );

    \I__9704\ : CascadeMux
    port map (
            O => \N__45868\,
            I => \N__45833\
        );

    \I__9703\ : InMux
    port map (
            O => \N__45867\,
            I => \N__45826\
        );

    \I__9702\ : InMux
    port map (
            O => \N__45866\,
            I => \N__45826\
        );

    \I__9701\ : Span4Mux_v
    port map (
            O => \N__45863\,
            I => \N__45819\
        );

    \I__9700\ : LocalMux
    port map (
            O => \N__45860\,
            I => \N__45819\
        );

    \I__9699\ : Span4Mux_v
    port map (
            O => \N__45857\,
            I => \N__45819\
        );

    \I__9698\ : Span4Mux_v
    port map (
            O => \N__45854\,
            I => \N__45814\
        );

    \I__9697\ : LocalMux
    port map (
            O => \N__45843\,
            I => \N__45814\
        );

    \I__9696\ : InMux
    port map (
            O => \N__45842\,
            I => \N__45811\
        );

    \I__9695\ : InMux
    port map (
            O => \N__45839\,
            I => \N__45808\
        );

    \I__9694\ : LocalMux
    port map (
            O => \N__45836\,
            I => \N__45805\
        );

    \I__9693\ : InMux
    port map (
            O => \N__45833\,
            I => \N__45798\
        );

    \I__9692\ : InMux
    port map (
            O => \N__45832\,
            I => \N__45798\
        );

    \I__9691\ : InMux
    port map (
            O => \N__45831\,
            I => \N__45798\
        );

    \I__9690\ : LocalMux
    port map (
            O => \N__45826\,
            I => \N__45795\
        );

    \I__9689\ : Span4Mux_h
    port map (
            O => \N__45819\,
            I => \N__45788\
        );

    \I__9688\ : Span4Mux_h
    port map (
            O => \N__45814\,
            I => \N__45788\
        );

    \I__9687\ : LocalMux
    port map (
            O => \N__45811\,
            I => \N__45788\
        );

    \I__9686\ : LocalMux
    port map (
            O => \N__45808\,
            I => \N__45781\
        );

    \I__9685\ : Sp12to4
    port map (
            O => \N__45805\,
            I => \N__45781\
        );

    \I__9684\ : LocalMux
    port map (
            O => \N__45798\,
            I => \N__45781\
        );

    \I__9683\ : Span4Mux_v
    port map (
            O => \N__45795\,
            I => \N__45776\
        );

    \I__9682\ : Span4Mux_h
    port map (
            O => \N__45788\,
            I => \N__45776\
        );

    \I__9681\ : Span12Mux_h
    port map (
            O => \N__45781\,
            I => \N__45773\
        );

    \I__9680\ : Odrv4
    port map (
            O => \N__45776\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271\
        );

    \I__9679\ : Odrv12
    port map (
            O => \N__45773\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271\
        );

    \I__9678\ : CascadeMux
    port map (
            O => \N__45768\,
            I => \N__45765\
        );

    \I__9677\ : InMux
    port map (
            O => \N__45765\,
            I => \N__45760\
        );

    \I__9676\ : InMux
    port map (
            O => \N__45764\,
            I => \N__45755\
        );

    \I__9675\ : InMux
    port map (
            O => \N__45763\,
            I => \N__45755\
        );

    \I__9674\ : LocalMux
    port map (
            O => \N__45760\,
            I => \N__45752\
        );

    \I__9673\ : LocalMux
    port map (
            O => \N__45755\,
            I => \N__45749\
        );

    \I__9672\ : Odrv4
    port map (
            O => \N__45752\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_21
        );

    \I__9671\ : Odrv4
    port map (
            O => \N__45749\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_21
        );

    \I__9670\ : InMux
    port map (
            O => \N__45744\,
            I => \N__45739\
        );

    \I__9669\ : CascadeMux
    port map (
            O => \N__45743\,
            I => \N__45736\
        );

    \I__9668\ : InMux
    port map (
            O => \N__45742\,
            I => \N__45733\
        );

    \I__9667\ : LocalMux
    port map (
            O => \N__45739\,
            I => \N__45730\
        );

    \I__9666\ : InMux
    port map (
            O => \N__45736\,
            I => \N__45727\
        );

    \I__9665\ : LocalMux
    port map (
            O => \N__45733\,
            I => \N__45724\
        );

    \I__9664\ : Span4Mux_h
    port map (
            O => \N__45730\,
            I => \N__45719\
        );

    \I__9663\ : LocalMux
    port map (
            O => \N__45727\,
            I => \N__45719\
        );

    \I__9662\ : Span4Mux_v
    port map (
            O => \N__45724\,
            I => \N__45714\
        );

    \I__9661\ : Span4Mux_v
    port map (
            O => \N__45719\,
            I => \N__45714\
        );

    \I__9660\ : Odrv4
    port map (
            O => \N__45714\,
            I => cemf_module_64ch_ctrl_inst1_data_config_21
        );

    \I__9659\ : CascadeMux
    port map (
            O => \N__45711\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_21_cascade_\
        );

    \I__9658\ : InMux
    port map (
            O => \N__45708\,
            I => \N__45705\
        );

    \I__9657\ : LocalMux
    port map (
            O => \N__45705\,
            I => \N__45702\
        );

    \I__9656\ : Odrv12
    port map (
            O => \N__45702\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDDZ0Z7\
        );

    \I__9655\ : InMux
    port map (
            O => \N__45699\,
            I => \N__45696\
        );

    \I__9654\ : LocalMux
    port map (
            O => \N__45696\,
            I => \N__45693\
        );

    \I__9653\ : Span4Mux_v
    port map (
            O => \N__45693\,
            I => \N__45688\
        );

    \I__9652\ : InMux
    port map (
            O => \N__45692\,
            I => \N__45683\
        );

    \I__9651\ : InMux
    port map (
            O => \N__45691\,
            I => \N__45683\
        );

    \I__9650\ : Odrv4
    port map (
            O => \N__45688\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_21
        );

    \I__9649\ : LocalMux
    port map (
            O => \N__45683\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_21
        );

    \I__9648\ : InMux
    port map (
            O => \N__45678\,
            I => \N__45675\
        );

    \I__9647\ : LocalMux
    port map (
            O => \N__45675\,
            I => \N__45671\
        );

    \I__9646\ : CascadeMux
    port map (
            O => \N__45674\,
            I => \N__45667\
        );

    \I__9645\ : Span4Mux_h
    port map (
            O => \N__45671\,
            I => \N__45664\
        );

    \I__9644\ : InMux
    port map (
            O => \N__45670\,
            I => \N__45661\
        );

    \I__9643\ : InMux
    port map (
            O => \N__45667\,
            I => \N__45658\
        );

    \I__9642\ : Odrv4
    port map (
            O => \N__45664\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_21
        );

    \I__9641\ : LocalMux
    port map (
            O => \N__45661\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_21
        );

    \I__9640\ : LocalMux
    port map (
            O => \N__45658\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_21
        );

    \I__9639\ : InMux
    port map (
            O => \N__45651\,
            I => \N__45648\
        );

    \I__9638\ : LocalMux
    port map (
            O => \N__45648\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_21\
        );

    \I__9637\ : CascadeMux
    port map (
            O => \N__45645\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_17_cascade_\
        );

    \I__9636\ : CascadeMux
    port map (
            O => \N__45642\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029DZ0Z7_cascade_\
        );

    \I__9635\ : InMux
    port map (
            O => \N__45639\,
            I => \N__45636\
        );

    \I__9634\ : LocalMux
    port map (
            O => \N__45636\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17\
        );

    \I__9633\ : CascadeMux
    port map (
            O => \N__45633\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17_cascade_\
        );

    \I__9632\ : InMux
    port map (
            O => \N__45630\,
            I => \N__45627\
        );

    \I__9631\ : LocalMux
    port map (
            O => \N__45627\,
            I => \N__45624\
        );

    \I__9630\ : Sp12to4
    port map (
            O => \N__45624\,
            I => \N__45621\
        );

    \I__9629\ : Odrv12
    port map (
            O => \N__45621\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_16\
        );

    \I__9628\ : CascadeMux
    port map (
            O => \N__45618\,
            I => \N__45614\
        );

    \I__9627\ : InMux
    port map (
            O => \N__45617\,
            I => \N__45610\
        );

    \I__9626\ : InMux
    port map (
            O => \N__45614\,
            I => \N__45605\
        );

    \I__9625\ : InMux
    port map (
            O => \N__45613\,
            I => \N__45605\
        );

    \I__9624\ : LocalMux
    port map (
            O => \N__45610\,
            I => \N__45602\
        );

    \I__9623\ : LocalMux
    port map (
            O => \N__45605\,
            I => \N__45599\
        );

    \I__9622\ : Odrv12
    port map (
            O => \N__45602\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_17
        );

    \I__9621\ : Odrv4
    port map (
            O => \N__45599\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_17
        );

    \I__9620\ : InMux
    port map (
            O => \N__45594\,
            I => \N__45591\
        );

    \I__9619\ : LocalMux
    port map (
            O => \N__45591\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_17\
        );

    \I__9618\ : InMux
    port map (
            O => \N__45588\,
            I => \N__45585\
        );

    \I__9617\ : LocalMux
    port map (
            O => \N__45585\,
            I => \N__45582\
        );

    \I__9616\ : Span4Mux_h
    port map (
            O => \N__45582\,
            I => \N__45579\
        );

    \I__9615\ : Sp12to4
    port map (
            O => \N__45579\,
            I => \N__45576\
        );

    \I__9614\ : Odrv12
    port map (
            O => \N__45576\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_3Z0Z_26\
        );

    \I__9613\ : CEMux
    port map (
            O => \N__45573\,
            I => \N__45552\
        );

    \I__9612\ : CEMux
    port map (
            O => \N__45572\,
            I => \N__45552\
        );

    \I__9611\ : CEMux
    port map (
            O => \N__45571\,
            I => \N__45552\
        );

    \I__9610\ : CEMux
    port map (
            O => \N__45570\,
            I => \N__45552\
        );

    \I__9609\ : CEMux
    port map (
            O => \N__45569\,
            I => \N__45552\
        );

    \I__9608\ : CEMux
    port map (
            O => \N__45568\,
            I => \N__45552\
        );

    \I__9607\ : CEMux
    port map (
            O => \N__45567\,
            I => \N__45552\
        );

    \I__9606\ : GlobalMux
    port map (
            O => \N__45552\,
            I => \N__45549\
        );

    \I__9605\ : gio2CtrlBuf
    port map (
            O => \N__45549\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g\
        );

    \I__9604\ : InMux
    port map (
            O => \N__45546\,
            I => \N__45543\
        );

    \I__9603\ : LocalMux
    port map (
            O => \N__45543\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_15\
        );

    \I__9602\ : InMux
    port map (
            O => \N__45540\,
            I => \N__45537\
        );

    \I__9601\ : LocalMux
    port map (
            O => \N__45537\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_16\
        );

    \I__9600\ : InMux
    port map (
            O => \N__45534\,
            I => \N__45531\
        );

    \I__9599\ : LocalMux
    port map (
            O => \N__45531\,
            I => \N__45526\
        );

    \I__9598\ : InMux
    port map (
            O => \N__45530\,
            I => \N__45523\
        );

    \I__9597\ : InMux
    port map (
            O => \N__45529\,
            I => \N__45520\
        );

    \I__9596\ : Odrv12
    port map (
            O => \N__45526\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_7
        );

    \I__9595\ : LocalMux
    port map (
            O => \N__45523\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_7
        );

    \I__9594\ : LocalMux
    port map (
            O => \N__45520\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_7
        );

    \I__9593\ : InMux
    port map (
            O => \N__45513\,
            I => \N__45510\
        );

    \I__9592\ : LocalMux
    port map (
            O => \N__45510\,
            I => \N__45507\
        );

    \I__9591\ : Span12Mux_v
    port map (
            O => \N__45507\,
            I => \N__45504\
        );

    \I__9590\ : Odrv12
    port map (
            O => \N__45504\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_7\
        );

    \I__9589\ : CascadeMux
    port map (
            O => \N__45501\,
            I => \serializer_mod_inst.un22_next_state_1_cascade_\
        );

    \I__9588\ : InMux
    port map (
            O => \N__45498\,
            I => \N__45495\
        );

    \I__9587\ : LocalMux
    port map (
            O => \N__45495\,
            I => \N__45492\
        );

    \I__9586\ : Span4Mux_h
    port map (
            O => \N__45492\,
            I => \N__45489\
        );

    \I__9585\ : Odrv4
    port map (
            O => \N__45489\,
            I => \serializer_mod_inst.un22_next_state\
        );

    \I__9584\ : InMux
    port map (
            O => \N__45486\,
            I => \N__45482\
        );

    \I__9583\ : InMux
    port map (
            O => \N__45485\,
            I => \N__45479\
        );

    \I__9582\ : LocalMux
    port map (
            O => \N__45482\,
            I => \N__45476\
        );

    \I__9581\ : LocalMux
    port map (
            O => \N__45479\,
            I => \N__45473\
        );

    \I__9580\ : Span4Mux_v
    port map (
            O => \N__45476\,
            I => \N__45470\
        );

    \I__9579\ : Span4Mux_v
    port map (
            O => \N__45473\,
            I => \N__45466\
        );

    \I__9578\ : Span4Mux_v
    port map (
            O => \N__45470\,
            I => \N__45438\
        );

    \I__9577\ : InMux
    port map (
            O => \N__45469\,
            I => \N__45435\
        );

    \I__9576\ : Span4Mux_v
    port map (
            O => \N__45466\,
            I => \N__45432\
        );

    \I__9575\ : CascadeMux
    port map (
            O => \N__45465\,
            I => \N__45429\
        );

    \I__9574\ : CascadeMux
    port map (
            O => \N__45464\,
            I => \N__45423\
        );

    \I__9573\ : CascadeMux
    port map (
            O => \N__45463\,
            I => \N__45419\
        );

    \I__9572\ : CascadeMux
    port map (
            O => \N__45462\,
            I => \N__45412\
        );

    \I__9571\ : InMux
    port map (
            O => \N__45461\,
            I => \N__45397\
        );

    \I__9570\ : InMux
    port map (
            O => \N__45460\,
            I => \N__45397\
        );

    \I__9569\ : InMux
    port map (
            O => \N__45459\,
            I => \N__45392\
        );

    \I__9568\ : InMux
    port map (
            O => \N__45458\,
            I => \N__45392\
        );

    \I__9567\ : InMux
    port map (
            O => \N__45457\,
            I => \N__45385\
        );

    \I__9566\ : InMux
    port map (
            O => \N__45456\,
            I => \N__45382\
        );

    \I__9565\ : InMux
    port map (
            O => \N__45455\,
            I => \N__45373\
        );

    \I__9564\ : InMux
    port map (
            O => \N__45454\,
            I => \N__45373\
        );

    \I__9563\ : InMux
    port map (
            O => \N__45453\,
            I => \N__45373\
        );

    \I__9562\ : InMux
    port map (
            O => \N__45452\,
            I => \N__45373\
        );

    \I__9561\ : InMux
    port map (
            O => \N__45451\,
            I => \N__45364\
        );

    \I__9560\ : InMux
    port map (
            O => \N__45450\,
            I => \N__45364\
        );

    \I__9559\ : InMux
    port map (
            O => \N__45449\,
            I => \N__45364\
        );

    \I__9558\ : InMux
    port map (
            O => \N__45448\,
            I => \N__45364\
        );

    \I__9557\ : InMux
    port map (
            O => \N__45447\,
            I => \N__45361\
        );

    \I__9556\ : InMux
    port map (
            O => \N__45446\,
            I => \N__45354\
        );

    \I__9555\ : InMux
    port map (
            O => \N__45445\,
            I => \N__45349\
        );

    \I__9554\ : InMux
    port map (
            O => \N__45444\,
            I => \N__45349\
        );

    \I__9553\ : InMux
    port map (
            O => \N__45443\,
            I => \N__45346\
        );

    \I__9552\ : InMux
    port map (
            O => \N__45442\,
            I => \N__45341\
        );

    \I__9551\ : InMux
    port map (
            O => \N__45441\,
            I => \N__45341\
        );

    \I__9550\ : Span4Mux_h
    port map (
            O => \N__45438\,
            I => \N__45336\
        );

    \I__9549\ : LocalMux
    port map (
            O => \N__45435\,
            I => \N__45336\
        );

    \I__9548\ : Span4Mux_v
    port map (
            O => \N__45432\,
            I => \N__45333\
        );

    \I__9547\ : InMux
    port map (
            O => \N__45429\,
            I => \N__45326\
        );

    \I__9546\ : InMux
    port map (
            O => \N__45428\,
            I => \N__45326\
        );

    \I__9545\ : InMux
    port map (
            O => \N__45427\,
            I => \N__45326\
        );

    \I__9544\ : InMux
    port map (
            O => \N__45426\,
            I => \N__45319\
        );

    \I__9543\ : InMux
    port map (
            O => \N__45423\,
            I => \N__45319\
        );

    \I__9542\ : InMux
    port map (
            O => \N__45422\,
            I => \N__45319\
        );

    \I__9541\ : InMux
    port map (
            O => \N__45419\,
            I => \N__45310\
        );

    \I__9540\ : InMux
    port map (
            O => \N__45418\,
            I => \N__45310\
        );

    \I__9539\ : InMux
    port map (
            O => \N__45417\,
            I => \N__45310\
        );

    \I__9538\ : InMux
    port map (
            O => \N__45416\,
            I => \N__45310\
        );

    \I__9537\ : InMux
    port map (
            O => \N__45415\,
            I => \N__45303\
        );

    \I__9536\ : InMux
    port map (
            O => \N__45412\,
            I => \N__45303\
        );

    \I__9535\ : InMux
    port map (
            O => \N__45411\,
            I => \N__45303\
        );

    \I__9534\ : InMux
    port map (
            O => \N__45410\,
            I => \N__45294\
        );

    \I__9533\ : InMux
    port map (
            O => \N__45409\,
            I => \N__45294\
        );

    \I__9532\ : InMux
    port map (
            O => \N__45408\,
            I => \N__45294\
        );

    \I__9531\ : InMux
    port map (
            O => \N__45407\,
            I => \N__45294\
        );

    \I__9530\ : InMux
    port map (
            O => \N__45406\,
            I => \N__45285\
        );

    \I__9529\ : InMux
    port map (
            O => \N__45405\,
            I => \N__45285\
        );

    \I__9528\ : InMux
    port map (
            O => \N__45404\,
            I => \N__45285\
        );

    \I__9527\ : InMux
    port map (
            O => \N__45403\,
            I => \N__45285\
        );

    \I__9526\ : InMux
    port map (
            O => \N__45402\,
            I => \N__45282\
        );

    \I__9525\ : LocalMux
    port map (
            O => \N__45397\,
            I => \N__45277\
        );

    \I__9524\ : LocalMux
    port map (
            O => \N__45392\,
            I => \N__45277\
        );

    \I__9523\ : InMux
    port map (
            O => \N__45391\,
            I => \N__45274\
        );

    \I__9522\ : InMux
    port map (
            O => \N__45390\,
            I => \N__45271\
        );

    \I__9521\ : InMux
    port map (
            O => \N__45389\,
            I => \N__45266\
        );

    \I__9520\ : InMux
    port map (
            O => \N__45388\,
            I => \N__45266\
        );

    \I__9519\ : LocalMux
    port map (
            O => \N__45385\,
            I => \N__45263\
        );

    \I__9518\ : LocalMux
    port map (
            O => \N__45382\,
            I => \N__45254\
        );

    \I__9517\ : LocalMux
    port map (
            O => \N__45373\,
            I => \N__45254\
        );

    \I__9516\ : LocalMux
    port map (
            O => \N__45364\,
            I => \N__45254\
        );

    \I__9515\ : LocalMux
    port map (
            O => \N__45361\,
            I => \N__45254\
        );

    \I__9514\ : InMux
    port map (
            O => \N__45360\,
            I => \N__45251\
        );

    \I__9513\ : InMux
    port map (
            O => \N__45359\,
            I => \N__45248\
        );

    \I__9512\ : CascadeMux
    port map (
            O => \N__45358\,
            I => \N__45236\
        );

    \I__9511\ : CascadeMux
    port map (
            O => \N__45357\,
            I => \N__45233\
        );

    \I__9510\ : LocalMux
    port map (
            O => \N__45354\,
            I => \N__45229\
        );

    \I__9509\ : LocalMux
    port map (
            O => \N__45349\,
            I => \N__45222\
        );

    \I__9508\ : LocalMux
    port map (
            O => \N__45346\,
            I => \N__45222\
        );

    \I__9507\ : LocalMux
    port map (
            O => \N__45341\,
            I => \N__45222\
        );

    \I__9506\ : Span4Mux_h
    port map (
            O => \N__45336\,
            I => \N__45205\
        );

    \I__9505\ : Span4Mux_h
    port map (
            O => \N__45333\,
            I => \N__45205\
        );

    \I__9504\ : LocalMux
    port map (
            O => \N__45326\,
            I => \N__45205\
        );

    \I__9503\ : LocalMux
    port map (
            O => \N__45319\,
            I => \N__45205\
        );

    \I__9502\ : LocalMux
    port map (
            O => \N__45310\,
            I => \N__45205\
        );

    \I__9501\ : LocalMux
    port map (
            O => \N__45303\,
            I => \N__45205\
        );

    \I__9500\ : LocalMux
    port map (
            O => \N__45294\,
            I => \N__45205\
        );

    \I__9499\ : LocalMux
    port map (
            O => \N__45285\,
            I => \N__45205\
        );

    \I__9498\ : LocalMux
    port map (
            O => \N__45282\,
            I => \N__45202\
        );

    \I__9497\ : Span4Mux_v
    port map (
            O => \N__45277\,
            I => \N__45194\
        );

    \I__9496\ : LocalMux
    port map (
            O => \N__45274\,
            I => \N__45194\
        );

    \I__9495\ : LocalMux
    port map (
            O => \N__45271\,
            I => \N__45194\
        );

    \I__9494\ : LocalMux
    port map (
            O => \N__45266\,
            I => \N__45191\
        );

    \I__9493\ : Span4Mux_v
    port map (
            O => \N__45263\,
            I => \N__45182\
        );

    \I__9492\ : Span4Mux_v
    port map (
            O => \N__45254\,
            I => \N__45182\
        );

    \I__9491\ : LocalMux
    port map (
            O => \N__45251\,
            I => \N__45182\
        );

    \I__9490\ : LocalMux
    port map (
            O => \N__45248\,
            I => \N__45182\
        );

    \I__9489\ : InMux
    port map (
            O => \N__45247\,
            I => \N__45179\
        );

    \I__9488\ : InMux
    port map (
            O => \N__45246\,
            I => \N__45169\
        );

    \I__9487\ : InMux
    port map (
            O => \N__45245\,
            I => \N__45169\
        );

    \I__9486\ : InMux
    port map (
            O => \N__45244\,
            I => \N__45162\
        );

    \I__9485\ : InMux
    port map (
            O => \N__45243\,
            I => \N__45162\
        );

    \I__9484\ : InMux
    port map (
            O => \N__45242\,
            I => \N__45162\
        );

    \I__9483\ : InMux
    port map (
            O => \N__45241\,
            I => \N__45155\
        );

    \I__9482\ : InMux
    port map (
            O => \N__45240\,
            I => \N__45155\
        );

    \I__9481\ : InMux
    port map (
            O => \N__45239\,
            I => \N__45155\
        );

    \I__9480\ : InMux
    port map (
            O => \N__45236\,
            I => \N__45148\
        );

    \I__9479\ : InMux
    port map (
            O => \N__45233\,
            I => \N__45148\
        );

    \I__9478\ : InMux
    port map (
            O => \N__45232\,
            I => \N__45148\
        );

    \I__9477\ : Span4Mux_v
    port map (
            O => \N__45229\,
            I => \N__45139\
        );

    \I__9476\ : Span4Mux_v
    port map (
            O => \N__45222\,
            I => \N__45139\
        );

    \I__9475\ : Span4Mux_v
    port map (
            O => \N__45205\,
            I => \N__45139\
        );

    \I__9474\ : Span4Mux_v
    port map (
            O => \N__45202\,
            I => \N__45139\
        );

    \I__9473\ : InMux
    port map (
            O => \N__45201\,
            I => \N__45136\
        );

    \I__9472\ : Span4Mux_h
    port map (
            O => \N__45194\,
            I => \N__45127\
        );

    \I__9471\ : Span4Mux_v
    port map (
            O => \N__45191\,
            I => \N__45127\
        );

    \I__9470\ : Span4Mux_h
    port map (
            O => \N__45182\,
            I => \N__45127\
        );

    \I__9469\ : LocalMux
    port map (
            O => \N__45179\,
            I => \N__45127\
        );

    \I__9468\ : InMux
    port map (
            O => \N__45178\,
            I => \N__45120\
        );

    \I__9467\ : InMux
    port map (
            O => \N__45177\,
            I => \N__45120\
        );

    \I__9466\ : InMux
    port map (
            O => \N__45176\,
            I => \N__45120\
        );

    \I__9465\ : InMux
    port map (
            O => \N__45175\,
            I => \N__45117\
        );

    \I__9464\ : InMux
    port map (
            O => \N__45174\,
            I => \N__45114\
        );

    \I__9463\ : LocalMux
    port map (
            O => \N__45169\,
            I => \N__45101\
        );

    \I__9462\ : LocalMux
    port map (
            O => \N__45162\,
            I => \N__45101\
        );

    \I__9461\ : LocalMux
    port map (
            O => \N__45155\,
            I => \N__45101\
        );

    \I__9460\ : LocalMux
    port map (
            O => \N__45148\,
            I => \N__45101\
        );

    \I__9459\ : Sp12to4
    port map (
            O => \N__45139\,
            I => \N__45101\
        );

    \I__9458\ : LocalMux
    port map (
            O => \N__45136\,
            I => \N__45101\
        );

    \I__9457\ : Odrv4
    port map (
            O => \N__45127\,
            I => \serializer_mod_inst.current_stateZ0Z_1\
        );

    \I__9456\ : LocalMux
    port map (
            O => \N__45120\,
            I => \serializer_mod_inst.current_stateZ0Z_1\
        );

    \I__9455\ : LocalMux
    port map (
            O => \N__45117\,
            I => \serializer_mod_inst.current_stateZ0Z_1\
        );

    \I__9454\ : LocalMux
    port map (
            O => \N__45114\,
            I => \serializer_mod_inst.current_stateZ0Z_1\
        );

    \I__9453\ : Odrv12
    port map (
            O => \N__45101\,
            I => \serializer_mod_inst.current_stateZ0Z_1\
        );

    \I__9452\ : InMux
    port map (
            O => \N__45090\,
            I => \N__45061\
        );

    \I__9451\ : InMux
    port map (
            O => \N__45089\,
            I => \N__45054\
        );

    \I__9450\ : InMux
    port map (
            O => \N__45088\,
            I => \N__45036\
        );

    \I__9449\ : InMux
    port map (
            O => \N__45087\,
            I => \N__45023\
        );

    \I__9448\ : InMux
    port map (
            O => \N__45086\,
            I => \N__45020\
        );

    \I__9447\ : InMux
    port map (
            O => \N__45085\,
            I => \N__45013\
        );

    \I__9446\ : InMux
    port map (
            O => \N__45084\,
            I => \N__45013\
        );

    \I__9445\ : InMux
    port map (
            O => \N__45083\,
            I => \N__45013\
        );

    \I__9444\ : InMux
    port map (
            O => \N__45082\,
            I => \N__45010\
        );

    \I__9443\ : InMux
    port map (
            O => \N__45081\,
            I => \N__44999\
        );

    \I__9442\ : InMux
    port map (
            O => \N__45080\,
            I => \N__44999\
        );

    \I__9441\ : InMux
    port map (
            O => \N__45079\,
            I => \N__44999\
        );

    \I__9440\ : InMux
    port map (
            O => \N__45078\,
            I => \N__44999\
        );

    \I__9439\ : InMux
    port map (
            O => \N__45077\,
            I => \N__44999\
        );

    \I__9438\ : InMux
    port map (
            O => \N__45076\,
            I => \N__44992\
        );

    \I__9437\ : InMux
    port map (
            O => \N__45075\,
            I => \N__44992\
        );

    \I__9436\ : InMux
    port map (
            O => \N__45074\,
            I => \N__44992\
        );

    \I__9435\ : InMux
    port map (
            O => \N__45073\,
            I => \N__44983\
        );

    \I__9434\ : InMux
    port map (
            O => \N__45072\,
            I => \N__44983\
        );

    \I__9433\ : InMux
    port map (
            O => \N__45071\,
            I => \N__44983\
        );

    \I__9432\ : InMux
    port map (
            O => \N__45070\,
            I => \N__44983\
        );

    \I__9431\ : InMux
    port map (
            O => \N__45069\,
            I => \N__44974\
        );

    \I__9430\ : InMux
    port map (
            O => \N__45068\,
            I => \N__44974\
        );

    \I__9429\ : InMux
    port map (
            O => \N__45067\,
            I => \N__44974\
        );

    \I__9428\ : InMux
    port map (
            O => \N__45066\,
            I => \N__44974\
        );

    \I__9427\ : InMux
    port map (
            O => \N__45065\,
            I => \N__44971\
        );

    \I__9426\ : InMux
    port map (
            O => \N__45064\,
            I => \N__44968\
        );

    \I__9425\ : LocalMux
    port map (
            O => \N__45061\,
            I => \N__44965\
        );

    \I__9424\ : InMux
    port map (
            O => \N__45060\,
            I => \N__44961\
        );

    \I__9423\ : InMux
    port map (
            O => \N__45059\,
            I => \N__44956\
        );

    \I__9422\ : InMux
    port map (
            O => \N__45058\,
            I => \N__44956\
        );

    \I__9421\ : InMux
    port map (
            O => \N__45057\,
            I => \N__44953\
        );

    \I__9420\ : LocalMux
    port map (
            O => \N__45054\,
            I => \N__44950\
        );

    \I__9419\ : InMux
    port map (
            O => \N__45053\,
            I => \N__44943\
        );

    \I__9418\ : InMux
    port map (
            O => \N__45052\,
            I => \N__44943\
        );

    \I__9417\ : InMux
    port map (
            O => \N__45051\,
            I => \N__44936\
        );

    \I__9416\ : InMux
    port map (
            O => \N__45050\,
            I => \N__44936\
        );

    \I__9415\ : InMux
    port map (
            O => \N__45049\,
            I => \N__44936\
        );

    \I__9414\ : InMux
    port map (
            O => \N__45048\,
            I => \N__44931\
        );

    \I__9413\ : InMux
    port map (
            O => \N__45047\,
            I => \N__44931\
        );

    \I__9412\ : InMux
    port map (
            O => \N__45046\,
            I => \N__44926\
        );

    \I__9411\ : InMux
    port map (
            O => \N__45045\,
            I => \N__44923\
        );

    \I__9410\ : InMux
    port map (
            O => \N__45044\,
            I => \N__44914\
        );

    \I__9409\ : InMux
    port map (
            O => \N__45043\,
            I => \N__44914\
        );

    \I__9408\ : InMux
    port map (
            O => \N__45042\,
            I => \N__44914\
        );

    \I__9407\ : InMux
    port map (
            O => \N__45041\,
            I => \N__44914\
        );

    \I__9406\ : InMux
    port map (
            O => \N__45040\,
            I => \N__44909\
        );

    \I__9405\ : InMux
    port map (
            O => \N__45039\,
            I => \N__44909\
        );

    \I__9404\ : LocalMux
    port map (
            O => \N__45036\,
            I => \N__44906\
        );

    \I__9403\ : InMux
    port map (
            O => \N__45035\,
            I => \N__44903\
        );

    \I__9402\ : InMux
    port map (
            O => \N__45034\,
            I => \N__44889\
        );

    \I__9401\ : InMux
    port map (
            O => \N__45033\,
            I => \N__44889\
        );

    \I__9400\ : InMux
    port map (
            O => \N__45032\,
            I => \N__44882\
        );

    \I__9399\ : InMux
    port map (
            O => \N__45031\,
            I => \N__44882\
        );

    \I__9398\ : InMux
    port map (
            O => \N__45030\,
            I => \N__44882\
        );

    \I__9397\ : InMux
    port map (
            O => \N__45029\,
            I => \N__44873\
        );

    \I__9396\ : InMux
    port map (
            O => \N__45028\,
            I => \N__44873\
        );

    \I__9395\ : InMux
    port map (
            O => \N__45027\,
            I => \N__44873\
        );

    \I__9394\ : InMux
    port map (
            O => \N__45026\,
            I => \N__44873\
        );

    \I__9393\ : LocalMux
    port map (
            O => \N__45023\,
            I => \N__44870\
        );

    \I__9392\ : LocalMux
    port map (
            O => \N__45020\,
            I => \N__44853\
        );

    \I__9391\ : LocalMux
    port map (
            O => \N__45013\,
            I => \N__44853\
        );

    \I__9390\ : LocalMux
    port map (
            O => \N__45010\,
            I => \N__44853\
        );

    \I__9389\ : LocalMux
    port map (
            O => \N__44999\,
            I => \N__44853\
        );

    \I__9388\ : LocalMux
    port map (
            O => \N__44992\,
            I => \N__44853\
        );

    \I__9387\ : LocalMux
    port map (
            O => \N__44983\,
            I => \N__44853\
        );

    \I__9386\ : LocalMux
    port map (
            O => \N__44974\,
            I => \N__44853\
        );

    \I__9385\ : LocalMux
    port map (
            O => \N__44971\,
            I => \N__44853\
        );

    \I__9384\ : LocalMux
    port map (
            O => \N__44968\,
            I => \N__44850\
        );

    \I__9383\ : Span4Mux_v
    port map (
            O => \N__44965\,
            I => \N__44847\
        );

    \I__9382\ : InMux
    port map (
            O => \N__44964\,
            I => \N__44844\
        );

    \I__9381\ : LocalMux
    port map (
            O => \N__44961\,
            I => \N__44835\
        );

    \I__9380\ : LocalMux
    port map (
            O => \N__44956\,
            I => \N__44835\
        );

    \I__9379\ : LocalMux
    port map (
            O => \N__44953\,
            I => \N__44835\
        );

    \I__9378\ : Span4Mux_h
    port map (
            O => \N__44950\,
            I => \N__44835\
        );

    \I__9377\ : InMux
    port map (
            O => \N__44949\,
            I => \N__44832\
        );

    \I__9376\ : InMux
    port map (
            O => \N__44948\,
            I => \N__44829\
        );

    \I__9375\ : LocalMux
    port map (
            O => \N__44943\,
            I => \N__44822\
        );

    \I__9374\ : LocalMux
    port map (
            O => \N__44936\,
            I => \N__44822\
        );

    \I__9373\ : LocalMux
    port map (
            O => \N__44931\,
            I => \N__44822\
        );

    \I__9372\ : InMux
    port map (
            O => \N__44930\,
            I => \N__44817\
        );

    \I__9371\ : InMux
    port map (
            O => \N__44929\,
            I => \N__44817\
        );

    \I__9370\ : LocalMux
    port map (
            O => \N__44926\,
            I => \N__44804\
        );

    \I__9369\ : LocalMux
    port map (
            O => \N__44923\,
            I => \N__44804\
        );

    \I__9368\ : LocalMux
    port map (
            O => \N__44914\,
            I => \N__44804\
        );

    \I__9367\ : LocalMux
    port map (
            O => \N__44909\,
            I => \N__44804\
        );

    \I__9366\ : Span4Mux_v
    port map (
            O => \N__44906\,
            I => \N__44804\
        );

    \I__9365\ : LocalMux
    port map (
            O => \N__44903\,
            I => \N__44804\
        );

    \I__9364\ : InMux
    port map (
            O => \N__44902\,
            I => \N__44801\
        );

    \I__9363\ : InMux
    port map (
            O => \N__44901\,
            I => \N__44796\
        );

    \I__9362\ : InMux
    port map (
            O => \N__44900\,
            I => \N__44796\
        );

    \I__9361\ : InMux
    port map (
            O => \N__44899\,
            I => \N__44793\
        );

    \I__9360\ : InMux
    port map (
            O => \N__44898\,
            I => \N__44788\
        );

    \I__9359\ : InMux
    port map (
            O => \N__44897\,
            I => \N__44788\
        );

    \I__9358\ : InMux
    port map (
            O => \N__44896\,
            I => \N__44781\
        );

    \I__9357\ : InMux
    port map (
            O => \N__44895\,
            I => \N__44781\
        );

    \I__9356\ : InMux
    port map (
            O => \N__44894\,
            I => \N__44781\
        );

    \I__9355\ : LocalMux
    port map (
            O => \N__44889\,
            I => \N__44776\
        );

    \I__9354\ : LocalMux
    port map (
            O => \N__44882\,
            I => \N__44776\
        );

    \I__9353\ : LocalMux
    port map (
            O => \N__44873\,
            I => \N__44771\
        );

    \I__9352\ : Span12Mux_h
    port map (
            O => \N__44870\,
            I => \N__44771\
        );

    \I__9351\ : Span4Mux_v
    port map (
            O => \N__44853\,
            I => \N__44766\
        );

    \I__9350\ : Span4Mux_v
    port map (
            O => \N__44850\,
            I => \N__44766\
        );

    \I__9349\ : Span4Mux_v
    port map (
            O => \N__44847\,
            I => \N__44763\
        );

    \I__9348\ : LocalMux
    port map (
            O => \N__44844\,
            I => \N__44758\
        );

    \I__9347\ : Span4Mux_v
    port map (
            O => \N__44835\,
            I => \N__44758\
        );

    \I__9346\ : LocalMux
    port map (
            O => \N__44832\,
            I => \N__44751\
        );

    \I__9345\ : LocalMux
    port map (
            O => \N__44829\,
            I => \N__44751\
        );

    \I__9344\ : Span4Mux_v
    port map (
            O => \N__44822\,
            I => \N__44751\
        );

    \I__9343\ : LocalMux
    port map (
            O => \N__44817\,
            I => \N__44746\
        );

    \I__9342\ : Span4Mux_v
    port map (
            O => \N__44804\,
            I => \N__44746\
        );

    \I__9341\ : LocalMux
    port map (
            O => \N__44801\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9340\ : LocalMux
    port map (
            O => \N__44796\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9339\ : LocalMux
    port map (
            O => \N__44793\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9338\ : LocalMux
    port map (
            O => \N__44788\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9337\ : LocalMux
    port map (
            O => \N__44781\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9336\ : Odrv4
    port map (
            O => \N__44776\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9335\ : Odrv12
    port map (
            O => \N__44771\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9334\ : Odrv4
    port map (
            O => \N__44766\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9333\ : Odrv4
    port map (
            O => \N__44763\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9332\ : Odrv4
    port map (
            O => \N__44758\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9331\ : Odrv4
    port map (
            O => \N__44751\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9330\ : Odrv4
    port map (
            O => \N__44746\,
            I => \serializer_mod_inst.current_stateZ0Z_0\
        );

    \I__9329\ : CascadeMux
    port map (
            O => \N__44721\,
            I => \N__44718\
        );

    \I__9328\ : InMux
    port map (
            O => \N__44718\,
            I => \N__44715\
        );

    \I__9327\ : LocalMux
    port map (
            O => \N__44715\,
            I => \N__44712\
        );

    \I__9326\ : Span4Mux_h
    port map (
            O => \N__44712\,
            I => \N__44709\
        );

    \I__9325\ : Odrv4
    port map (
            O => \N__44709\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_0\
        );

    \I__9324\ : InMux
    port map (
            O => \N__44706\,
            I => \N__44703\
        );

    \I__9323\ : LocalMux
    port map (
            O => \N__44703\,
            I => \N__44700\
        );

    \I__9322\ : Span4Mux_h
    port map (
            O => \N__44700\,
            I => \N__44697\
        );

    \I__9321\ : Span4Mux_h
    port map (
            O => \N__44697\,
            I => \N__44694\
        );

    \I__9320\ : Odrv4
    port map (
            O => \N__44694\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_0\
        );

    \I__9319\ : InMux
    port map (
            O => \N__44691\,
            I => \N__44688\
        );

    \I__9318\ : LocalMux
    port map (
            O => \N__44688\,
            I => \N__44685\
        );

    \I__9317\ : Span12Mux_v
    port map (
            O => \N__44685\,
            I => \N__44682\
        );

    \I__9316\ : Span12Mux_h
    port map (
            O => \N__44682\,
            I => \N__44679\
        );

    \I__9315\ : Odrv12
    port map (
            O => \N__44679\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_0
        );

    \I__9314\ : InMux
    port map (
            O => \N__44676\,
            I => \N__44672\
        );

    \I__9313\ : InMux
    port map (
            O => \N__44675\,
            I => \N__44669\
        );

    \I__9312\ : LocalMux
    port map (
            O => \N__44672\,
            I => \N__44666\
        );

    \I__9311\ : LocalMux
    port map (
            O => \N__44669\,
            I => \N__44654\
        );

    \I__9310\ : Span4Mux_h
    port map (
            O => \N__44666\,
            I => \N__44651\
        );

    \I__9309\ : CascadeMux
    port map (
            O => \N__44665\,
            I => \N__44648\
        );

    \I__9308\ : InMux
    port map (
            O => \N__44664\,
            I => \N__44644\
        );

    \I__9307\ : InMux
    port map (
            O => \N__44663\,
            I => \N__44641\
        );

    \I__9306\ : CascadeMux
    port map (
            O => \N__44662\,
            I => \N__44636\
        );

    \I__9305\ : InMux
    port map (
            O => \N__44661\,
            I => \N__44632\
        );

    \I__9304\ : CascadeMux
    port map (
            O => \N__44660\,
            I => \N__44629\
        );

    \I__9303\ : CascadeMux
    port map (
            O => \N__44659\,
            I => \N__44625\
        );

    \I__9302\ : InMux
    port map (
            O => \N__44658\,
            I => \N__44621\
        );

    \I__9301\ : InMux
    port map (
            O => \N__44657\,
            I => \N__44618\
        );

    \I__9300\ : Span4Mux_h
    port map (
            O => \N__44654\,
            I => \N__44609\
        );

    \I__9299\ : Span4Mux_h
    port map (
            O => \N__44651\,
            I => \N__44609\
        );

    \I__9298\ : InMux
    port map (
            O => \N__44648\,
            I => \N__44606\
        );

    \I__9297\ : CascadeMux
    port map (
            O => \N__44647\,
            I => \N__44603\
        );

    \I__9296\ : LocalMux
    port map (
            O => \N__44644\,
            I => \N__44598\
        );

    \I__9295\ : LocalMux
    port map (
            O => \N__44641\,
            I => \N__44598\
        );

    \I__9294\ : InMux
    port map (
            O => \N__44640\,
            I => \N__44593\
        );

    \I__9293\ : InMux
    port map (
            O => \N__44639\,
            I => \N__44593\
        );

    \I__9292\ : InMux
    port map (
            O => \N__44636\,
            I => \N__44585\
        );

    \I__9291\ : InMux
    port map (
            O => \N__44635\,
            I => \N__44585\
        );

    \I__9290\ : LocalMux
    port map (
            O => \N__44632\,
            I => \N__44582\
        );

    \I__9289\ : InMux
    port map (
            O => \N__44629\,
            I => \N__44577\
        );

    \I__9288\ : InMux
    port map (
            O => \N__44628\,
            I => \N__44577\
        );

    \I__9287\ : InMux
    port map (
            O => \N__44625\,
            I => \N__44572\
        );

    \I__9286\ : InMux
    port map (
            O => \N__44624\,
            I => \N__44572\
        );

    \I__9285\ : LocalMux
    port map (
            O => \N__44621\,
            I => \N__44567\
        );

    \I__9284\ : LocalMux
    port map (
            O => \N__44618\,
            I => \N__44567\
        );

    \I__9283\ : InMux
    port map (
            O => \N__44617\,
            I => \N__44564\
        );

    \I__9282\ : InMux
    port map (
            O => \N__44616\,
            I => \N__44557\
        );

    \I__9281\ : InMux
    port map (
            O => \N__44615\,
            I => \N__44557\
        );

    \I__9280\ : InMux
    port map (
            O => \N__44614\,
            I => \N__44557\
        );

    \I__9279\ : Span4Mux_h
    port map (
            O => \N__44609\,
            I => \N__44552\
        );

    \I__9278\ : LocalMux
    port map (
            O => \N__44606\,
            I => \N__44552\
        );

    \I__9277\ : InMux
    port map (
            O => \N__44603\,
            I => \N__44549\
        );

    \I__9276\ : Sp12to4
    port map (
            O => \N__44598\,
            I => \N__44542\
        );

    \I__9275\ : LocalMux
    port map (
            O => \N__44593\,
            I => \N__44542\
        );

    \I__9274\ : CascadeMux
    port map (
            O => \N__44592\,
            I => \N__44538\
        );

    \I__9273\ : CascadeMux
    port map (
            O => \N__44591\,
            I => \N__44535\
        );

    \I__9272\ : InMux
    port map (
            O => \N__44590\,
            I => \N__44530\
        );

    \I__9271\ : LocalMux
    port map (
            O => \N__44585\,
            I => \N__44527\
        );

    \I__9270\ : Span4Mux_v
    port map (
            O => \N__44582\,
            I => \N__44518\
        );

    \I__9269\ : LocalMux
    port map (
            O => \N__44577\,
            I => \N__44518\
        );

    \I__9268\ : LocalMux
    port map (
            O => \N__44572\,
            I => \N__44518\
        );

    \I__9267\ : Span4Mux_h
    port map (
            O => \N__44567\,
            I => \N__44518\
        );

    \I__9266\ : LocalMux
    port map (
            O => \N__44564\,
            I => \N__44515\
        );

    \I__9265\ : LocalMux
    port map (
            O => \N__44557\,
            I => \N__44510\
        );

    \I__9264\ : Span4Mux_h
    port map (
            O => \N__44552\,
            I => \N__44510\
        );

    \I__9263\ : LocalMux
    port map (
            O => \N__44549\,
            I => \N__44505\
        );

    \I__9262\ : InMux
    port map (
            O => \N__44548\,
            I => \N__44500\
        );

    \I__9261\ : InMux
    port map (
            O => \N__44547\,
            I => \N__44500\
        );

    \I__9260\ : Span12Mux_s11_v
    port map (
            O => \N__44542\,
            I => \N__44497\
        );

    \I__9259\ : InMux
    port map (
            O => \N__44541\,
            I => \N__44486\
        );

    \I__9258\ : InMux
    port map (
            O => \N__44538\,
            I => \N__44486\
        );

    \I__9257\ : InMux
    port map (
            O => \N__44535\,
            I => \N__44486\
        );

    \I__9256\ : InMux
    port map (
            O => \N__44534\,
            I => \N__44486\
        );

    \I__9255\ : InMux
    port map (
            O => \N__44533\,
            I => \N__44486\
        );

    \I__9254\ : LocalMux
    port map (
            O => \N__44530\,
            I => \N__44479\
        );

    \I__9253\ : Span4Mux_v
    port map (
            O => \N__44527\,
            I => \N__44479\
        );

    \I__9252\ : Span4Mux_h
    port map (
            O => \N__44518\,
            I => \N__44479\
        );

    \I__9251\ : Span4Mux_v
    port map (
            O => \N__44515\,
            I => \N__44474\
        );

    \I__9250\ : Span4Mux_v
    port map (
            O => \N__44510\,
            I => \N__44474\
        );

    \I__9249\ : InMux
    port map (
            O => \N__44509\,
            I => \N__44469\
        );

    \I__9248\ : InMux
    port map (
            O => \N__44508\,
            I => \N__44469\
        );

    \I__9247\ : Odrv12
    port map (
            O => \N__44505\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9246\ : LocalMux
    port map (
            O => \N__44500\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9245\ : Odrv12
    port map (
            O => \N__44497\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9244\ : LocalMux
    port map (
            O => \N__44486\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9243\ : Odrv4
    port map (
            O => \N__44479\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9242\ : Odrv4
    port map (
            O => \N__44474\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9241\ : LocalMux
    port map (
            O => \N__44469\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\
        );

    \I__9240\ : CascadeMux
    port map (
            O => \N__44454\,
            I => \N__44451\
        );

    \I__9239\ : InMux
    port map (
            O => \N__44451\,
            I => \N__44448\
        );

    \I__9238\ : LocalMux
    port map (
            O => \N__44448\,
            I => \N__44445\
        );

    \I__9237\ : Span4Mux_h
    port map (
            O => \N__44445\,
            I => \N__44442\
        );

    \I__9236\ : Sp12to4
    port map (
            O => \N__44442\,
            I => \N__44439\
        );

    \I__9235\ : Span12Mux_v
    port map (
            O => \N__44439\,
            I => \N__44436\
        );

    \I__9234\ : Odrv12
    port map (
            O => \N__44436\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_0\
        );

    \I__9233\ : InMux
    port map (
            O => \N__44433\,
            I => \N__44428\
        );

    \I__9232\ : InMux
    port map (
            O => \N__44432\,
            I => \N__44422\
        );

    \I__9231\ : InMux
    port map (
            O => \N__44431\,
            I => \N__44422\
        );

    \I__9230\ : LocalMux
    port map (
            O => \N__44428\,
            I => \N__44419\
        );

    \I__9229\ : InMux
    port map (
            O => \N__44427\,
            I => \N__44415\
        );

    \I__9228\ : LocalMux
    port map (
            O => \N__44422\,
            I => \N__44410\
        );

    \I__9227\ : Span4Mux_h
    port map (
            O => \N__44419\,
            I => \N__44403\
        );

    \I__9226\ : InMux
    port map (
            O => \N__44418\,
            I => \N__44400\
        );

    \I__9225\ : LocalMux
    port map (
            O => \N__44415\,
            I => \N__44397\
        );

    \I__9224\ : InMux
    port map (
            O => \N__44414\,
            I => \N__44394\
        );

    \I__9223\ : InMux
    port map (
            O => \N__44413\,
            I => \N__44391\
        );

    \I__9222\ : Span4Mux_h
    port map (
            O => \N__44410\,
            I => \N__44388\
        );

    \I__9221\ : InMux
    port map (
            O => \N__44409\,
            I => \N__44383\
        );

    \I__9220\ : InMux
    port map (
            O => \N__44408\,
            I => \N__44383\
        );

    \I__9219\ : InMux
    port map (
            O => \N__44407\,
            I => \N__44378\
        );

    \I__9218\ : InMux
    port map (
            O => \N__44406\,
            I => \N__44378\
        );

    \I__9217\ : Span4Mux_h
    port map (
            O => \N__44403\,
            I => \N__44373\
        );

    \I__9216\ : LocalMux
    port map (
            O => \N__44400\,
            I => \N__44373\
        );

    \I__9215\ : Span4Mux_h
    port map (
            O => \N__44397\,
            I => \N__44360\
        );

    \I__9214\ : LocalMux
    port map (
            O => \N__44394\,
            I => \N__44360\
        );

    \I__9213\ : LocalMux
    port map (
            O => \N__44391\,
            I => \N__44360\
        );

    \I__9212\ : Span4Mux_h
    port map (
            O => \N__44388\,
            I => \N__44355\
        );

    \I__9211\ : LocalMux
    port map (
            O => \N__44383\,
            I => \N__44355\
        );

    \I__9210\ : LocalMux
    port map (
            O => \N__44378\,
            I => \N__44350\
        );

    \I__9209\ : Span4Mux_h
    port map (
            O => \N__44373\,
            I => \N__44350\
        );

    \I__9208\ : InMux
    port map (
            O => \N__44372\,
            I => \N__44343\
        );

    \I__9207\ : InMux
    port map (
            O => \N__44371\,
            I => \N__44343\
        );

    \I__9206\ : InMux
    port map (
            O => \N__44370\,
            I => \N__44343\
        );

    \I__9205\ : InMux
    port map (
            O => \N__44369\,
            I => \N__44340\
        );

    \I__9204\ : InMux
    port map (
            O => \N__44368\,
            I => \N__44335\
        );

    \I__9203\ : InMux
    port map (
            O => \N__44367\,
            I => \N__44335\
        );

    \I__9202\ : Span4Mux_h
    port map (
            O => \N__44360\,
            I => \N__44323\
        );

    \I__9201\ : Span4Mux_h
    port map (
            O => \N__44355\,
            I => \N__44320\
        );

    \I__9200\ : Span4Mux_v
    port map (
            O => \N__44350\,
            I => \N__44315\
        );

    \I__9199\ : LocalMux
    port map (
            O => \N__44343\,
            I => \N__44315\
        );

    \I__9198\ : LocalMux
    port map (
            O => \N__44340\,
            I => \N__44310\
        );

    \I__9197\ : LocalMux
    port map (
            O => \N__44335\,
            I => \N__44310\
        );

    \I__9196\ : InMux
    port map (
            O => \N__44334\,
            I => \N__44305\
        );

    \I__9195\ : InMux
    port map (
            O => \N__44333\,
            I => \N__44305\
        );

    \I__9194\ : InMux
    port map (
            O => \N__44332\,
            I => \N__44300\
        );

    \I__9193\ : InMux
    port map (
            O => \N__44331\,
            I => \N__44300\
        );

    \I__9192\ : InMux
    port map (
            O => \N__44330\,
            I => \N__44289\
        );

    \I__9191\ : InMux
    port map (
            O => \N__44329\,
            I => \N__44289\
        );

    \I__9190\ : InMux
    port map (
            O => \N__44328\,
            I => \N__44289\
        );

    \I__9189\ : InMux
    port map (
            O => \N__44327\,
            I => \N__44289\
        );

    \I__9188\ : InMux
    port map (
            O => \N__44326\,
            I => \N__44289\
        );

    \I__9187\ : Odrv4
    port map (
            O => \N__44323\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9186\ : Odrv4
    port map (
            O => \N__44320\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9185\ : Odrv4
    port map (
            O => \N__44315\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9184\ : Odrv12
    port map (
            O => \N__44310\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9183\ : LocalMux
    port map (
            O => \N__44305\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9182\ : LocalMux
    port map (
            O => \N__44300\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9181\ : LocalMux
    port map (
            O => \N__44289\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\
        );

    \I__9180\ : InMux
    port map (
            O => \N__44274\,
            I => \N__44271\
        );

    \I__9179\ : LocalMux
    port map (
            O => \N__44271\,
            I => \N__44268\
        );

    \I__9178\ : Span4Mux_h
    port map (
            O => \N__44268\,
            I => \N__44265\
        );

    \I__9177\ : Span4Mux_v
    port map (
            O => \N__44265\,
            I => \N__44262\
        );

    \I__9176\ : Span4Mux_h
    port map (
            O => \N__44262\,
            I => \N__44259\
        );

    \I__9175\ : Span4Mux_h
    port map (
            O => \N__44259\,
            I => \N__44256\
        );

    \I__9174\ : Odrv4
    port map (
            O => \N__44256\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_940\
        );

    \I__9173\ : CascadeMux
    port map (
            O => \N__44253\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_cascade_\
        );

    \I__9172\ : InMux
    port map (
            O => \N__44250\,
            I => \N__44247\
        );

    \I__9171\ : LocalMux
    port map (
            O => \N__44247\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_0\
        );

    \I__9170\ : InMux
    port map (
            O => \N__44244\,
            I => \N__44241\
        );

    \I__9169\ : LocalMux
    port map (
            O => \N__44241\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_0\
        );

    \I__9168\ : CascadeMux
    port map (
            O => \N__44238\,
            I => \N__44235\
        );

    \I__9167\ : InMux
    port map (
            O => \N__44235\,
            I => \N__44232\
        );

    \I__9166\ : LocalMux
    port map (
            O => \N__44232\,
            I => \N__44229\
        );

    \I__9165\ : Span4Mux_v
    port map (
            O => \N__44229\,
            I => \N__44226\
        );

    \I__9164\ : Span4Mux_h
    port map (
            O => \N__44226\,
            I => \N__44223\
        );

    \I__9163\ : Odrv4
    port map (
            O => \N__44223\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_25\
        );

    \I__9162\ : InMux
    port map (
            O => \N__44220\,
            I => \N__44217\
        );

    \I__9161\ : LocalMux
    port map (
            O => \N__44217\,
            I => \serializer_mod_inst.shift_regZ0Z_29\
        );

    \I__9160\ : InMux
    port map (
            O => \N__44214\,
            I => \N__44211\
        );

    \I__9159\ : LocalMux
    port map (
            O => \N__44211\,
            I => \N__44208\
        );

    \I__9158\ : Odrv12
    port map (
            O => \N__44208\,
            I => \serializer_mod_inst.shift_regZ0Z_30\
        );

    \I__9157\ : InMux
    port map (
            O => \N__44205\,
            I => \N__44202\
        );

    \I__9156\ : LocalMux
    port map (
            O => \N__44202\,
            I => \serializer_mod_inst.shift_regZ0Z_62\
        );

    \I__9155\ : InMux
    port map (
            O => \N__44199\,
            I => \N__44196\
        );

    \I__9154\ : LocalMux
    port map (
            O => \N__44196\,
            I => \serializer_mod_inst.shift_regZ0Z_63\
        );

    \I__9153\ : InMux
    port map (
            O => \N__44193\,
            I => \N__44190\
        );

    \I__9152\ : LocalMux
    port map (
            O => \N__44190\,
            I => \serializer_mod_inst.shift_regZ0Z_58\
        );

    \I__9151\ : InMux
    port map (
            O => \N__44187\,
            I => \N__44184\
        );

    \I__9150\ : LocalMux
    port map (
            O => \N__44184\,
            I => \serializer_mod_inst.shift_regZ0Z_59\
        );

    \I__9149\ : InMux
    port map (
            O => \N__44181\,
            I => \N__44178\
        );

    \I__9148\ : LocalMux
    port map (
            O => \N__44178\,
            I => \serializer_mod_inst.shift_regZ0Z_60\
        );

    \I__9147\ : InMux
    port map (
            O => \N__44175\,
            I => \N__44172\
        );

    \I__9146\ : LocalMux
    port map (
            O => \N__44172\,
            I => \serializer_mod_inst.shift_regZ0Z_61\
        );

    \I__9145\ : InMux
    port map (
            O => \N__44169\,
            I => \N__44166\
        );

    \I__9144\ : LocalMux
    port map (
            O => \N__44166\,
            I => \N__44163\
        );

    \I__9143\ : Span4Mux_h
    port map (
            O => \N__44163\,
            I => \N__44160\
        );

    \I__9142\ : Odrv4
    port map (
            O => \N__44160\,
            I => \serializer_mod_inst.shift_regZ0Z_56\
        );

    \I__9141\ : InMux
    port map (
            O => \N__44157\,
            I => \N__44154\
        );

    \I__9140\ : LocalMux
    port map (
            O => \N__44154\,
            I => \serializer_mod_inst.shift_regZ0Z_57\
        );

    \I__9139\ : CascadeMux
    port map (
            O => \N__44151\,
            I => \N__44148\
        );

    \I__9138\ : InMux
    port map (
            O => \N__44148\,
            I => \N__44145\
        );

    \I__9137\ : LocalMux
    port map (
            O => \N__44145\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_3\
        );

    \I__9136\ : InMux
    port map (
            O => \N__44142\,
            I => \N__44135\
        );

    \I__9135\ : InMux
    port map (
            O => \N__44141\,
            I => \N__44135\
        );

    \I__9134\ : InMux
    port map (
            O => \N__44140\,
            I => \N__44132\
        );

    \I__9133\ : LocalMux
    port map (
            O => \N__44135\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0\
        );

    \I__9132\ : LocalMux
    port map (
            O => \N__44132\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0\
        );

    \I__9131\ : CascadeMux
    port map (
            O => \N__44127\,
            I => \N__44124\
        );

    \I__9130\ : InMux
    port map (
            O => \N__44124\,
            I => \N__44121\
        );

    \I__9129\ : LocalMux
    port map (
            O => \N__44121\,
            I => \N__44118\
        );

    \I__9128\ : Sp12to4
    port map (
            O => \N__44118\,
            I => \N__44115\
        );

    \I__9127\ : Span12Mux_s8_h
    port map (
            O => \N__44115\,
            I => \N__44112\
        );

    \I__9126\ : Span12Mux_v
    port map (
            O => \N__44112\,
            I => \N__44109\
        );

    \I__9125\ : Odrv12
    port map (
            O => \N__44109\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_1\
        );

    \I__9124\ : CEMux
    port map (
            O => \N__44106\,
            I => \N__44102\
        );

    \I__9123\ : CEMux
    port map (
            O => \N__44105\,
            I => \N__44099\
        );

    \I__9122\ : LocalMux
    port map (
            O => \N__44102\,
            I => \N__44096\
        );

    \I__9121\ : LocalMux
    port map (
            O => \N__44099\,
            I => \N__44093\
        );

    \I__9120\ : Span4Mux_h
    port map (
            O => \N__44096\,
            I => \N__44089\
        );

    \I__9119\ : Span4Mux_v
    port map (
            O => \N__44093\,
            I => \N__44085\
        );

    \I__9118\ : CEMux
    port map (
            O => \N__44092\,
            I => \N__44082\
        );

    \I__9117\ : Span4Mux_v
    port map (
            O => \N__44089\,
            I => \N__44079\
        );

    \I__9116\ : CEMux
    port map (
            O => \N__44088\,
            I => \N__44076\
        );

    \I__9115\ : Span4Mux_h
    port map (
            O => \N__44085\,
            I => \N__44071\
        );

    \I__9114\ : LocalMux
    port map (
            O => \N__44082\,
            I => \N__44071\
        );

    \I__9113\ : Span4Mux_v
    port map (
            O => \N__44079\,
            I => \N__44068\
        );

    \I__9112\ : LocalMux
    port map (
            O => \N__44076\,
            I => \N__44065\
        );

    \I__9111\ : Span4Mux_h
    port map (
            O => \N__44071\,
            I => \N__44062\
        );

    \I__9110\ : Span4Mux_v
    port map (
            O => \N__44068\,
            I => \N__44058\
        );

    \I__9109\ : Span4Mux_v
    port map (
            O => \N__44065\,
            I => \N__44055\
        );

    \I__9108\ : Sp12to4
    port map (
            O => \N__44062\,
            I => \N__44052\
        );

    \I__9107\ : CEMux
    port map (
            O => \N__44061\,
            I => \N__44049\
        );

    \I__9106\ : Span4Mux_h
    port map (
            O => \N__44058\,
            I => \N__44046\
        );

    \I__9105\ : Span4Mux_h
    port map (
            O => \N__44055\,
            I => \N__44043\
        );

    \I__9104\ : Span12Mux_v
    port map (
            O => \N__44052\,
            I => \N__44040\
        );

    \I__9103\ : LocalMux
    port map (
            O => \N__44049\,
            I => \N__44035\
        );

    \I__9102\ : Span4Mux_h
    port map (
            O => \N__44046\,
            I => \N__44035\
        );

    \I__9101\ : Sp12to4
    port map (
            O => \N__44043\,
            I => \N__44030\
        );

    \I__9100\ : Span12Mux_h
    port map (
            O => \N__44040\,
            I => \N__44030\
        );

    \I__9099\ : Odrv4
    port map (
            O => \N__44035\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0\
        );

    \I__9098\ : Odrv12
    port map (
            O => \N__44030\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0\
        );

    \I__9097\ : InMux
    port map (
            O => \N__44025\,
            I => \N__44022\
        );

    \I__9096\ : LocalMux
    port map (
            O => \N__44022\,
            I => \serializer_mod_inst.shift_regZ0Z_64\
        );

    \I__9095\ : InMux
    port map (
            O => \N__44019\,
            I => \N__44016\
        );

    \I__9094\ : LocalMux
    port map (
            O => \N__44016\,
            I => \N__44013\
        );

    \I__9093\ : Span4Mux_h
    port map (
            O => \N__44013\,
            I => \N__44010\
        );

    \I__9092\ : Odrv4
    port map (
            O => \N__44010\,
            I => \serializer_mod_inst.shift_regZ0Z_65\
        );

    \I__9091\ : InMux
    port map (
            O => \N__44007\,
            I => \N__44004\
        );

    \I__9090\ : LocalMux
    port map (
            O => \N__44004\,
            I => \N__44000\
        );

    \I__9089\ : InMux
    port map (
            O => \N__44003\,
            I => \N__43997\
        );

    \I__9088\ : Span4Mux_h
    port map (
            O => \N__44000\,
            I => \N__43994\
        );

    \I__9087\ : LocalMux
    port map (
            O => \N__43997\,
            I => \N__43991\
        );

    \I__9086\ : Span4Mux_v
    port map (
            O => \N__43994\,
            I => \N__43988\
        );

    \I__9085\ : Span4Mux_h
    port map (
            O => \N__43991\,
            I => \N__43985\
        );

    \I__9084\ : Span4Mux_v
    port map (
            O => \N__43988\,
            I => \N__43982\
        );

    \I__9083\ : Span4Mux_v
    port map (
            O => \N__43985\,
            I => \N__43979\
        );

    \I__9082\ : Odrv4
    port map (
            O => \N__43982\,
            I => \serializer_mod_inst.shift_regZ0Z_128\
        );

    \I__9081\ : Odrv4
    port map (
            O => \N__43979\,
            I => \serializer_mod_inst.shift_regZ0Z_128\
        );

    \I__9080\ : InMux
    port map (
            O => \N__43974\,
            I => \N__43971\
        );

    \I__9079\ : LocalMux
    port map (
            O => \N__43971\,
            I => \serializer_mod_inst.shift_regZ0Z_126\
        );

    \I__9078\ : InMux
    port map (
            O => \N__43968\,
            I => \N__43965\
        );

    \I__9077\ : LocalMux
    port map (
            O => \N__43965\,
            I => \serializer_mod_inst.shift_regZ0Z_127\
        );

    \I__9076\ : InMux
    port map (
            O => \N__43962\,
            I => \N__43959\
        );

    \I__9075\ : LocalMux
    port map (
            O => \N__43959\,
            I => \serializer_mod_inst.shift_regZ0Z_28\
        );

    \I__9074\ : InMux
    port map (
            O => \N__43956\,
            I => \N__43951\
        );

    \I__9073\ : InMux
    port map (
            O => \N__43955\,
            I => \N__43948\
        );

    \I__9072\ : InMux
    port map (
            O => \N__43954\,
            I => \N__43945\
        );

    \I__9071\ : LocalMux
    port map (
            O => \N__43951\,
            I => \N__43942\
        );

    \I__9070\ : LocalMux
    port map (
            O => \N__43948\,
            I => \N__43939\
        );

    \I__9069\ : LocalMux
    port map (
            O => \N__43945\,
            I => \N__43933\
        );

    \I__9068\ : Span4Mux_v
    port map (
            O => \N__43942\,
            I => \N__43933\
        );

    \I__9067\ : Span4Mux_h
    port map (
            O => \N__43939\,
            I => \N__43928\
        );

    \I__9066\ : InMux
    port map (
            O => \N__43938\,
            I => \N__43925\
        );

    \I__9065\ : Sp12to4
    port map (
            O => \N__43933\,
            I => \N__43922\
        );

    \I__9064\ : InMux
    port map (
            O => \N__43932\,
            I => \N__43917\
        );

    \I__9063\ : InMux
    port map (
            O => \N__43931\,
            I => \N__43917\
        );

    \I__9062\ : Span4Mux_h
    port map (
            O => \N__43928\,
            I => \N__43914\
        );

    \I__9061\ : LocalMux
    port map (
            O => \N__43925\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13\
        );

    \I__9060\ : Odrv12
    port map (
            O => \N__43922\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13\
        );

    \I__9059\ : LocalMux
    port map (
            O => \N__43917\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13\
        );

    \I__9058\ : Odrv4
    port map (
            O => \N__43914\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13\
        );

    \I__9057\ : InMux
    port map (
            O => \N__43905\,
            I => \N__43898\
        );

    \I__9056\ : InMux
    port map (
            O => \N__43904\,
            I => \N__43891\
        );

    \I__9055\ : InMux
    port map (
            O => \N__43903\,
            I => \N__43891\
        );

    \I__9054\ : InMux
    port map (
            O => \N__43902\,
            I => \N__43891\
        );

    \I__9053\ : CascadeMux
    port map (
            O => \N__43901\,
            I => \N__43888\
        );

    \I__9052\ : LocalMux
    port map (
            O => \N__43898\,
            I => \N__43882\
        );

    \I__9051\ : LocalMux
    port map (
            O => \N__43891\,
            I => \N__43879\
        );

    \I__9050\ : InMux
    port map (
            O => \N__43888\,
            I => \N__43874\
        );

    \I__9049\ : InMux
    port map (
            O => \N__43887\,
            I => \N__43874\
        );

    \I__9048\ : InMux
    port map (
            O => \N__43886\,
            I => \N__43869\
        );

    \I__9047\ : InMux
    port map (
            O => \N__43885\,
            I => \N__43869\
        );

    \I__9046\ : Span4Mux_v
    port map (
            O => \N__43882\,
            I => \N__43866\
        );

    \I__9045\ : Odrv4
    port map (
            O => \N__43879\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3\
        );

    \I__9044\ : LocalMux
    port map (
            O => \N__43874\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3\
        );

    \I__9043\ : LocalMux
    port map (
            O => \N__43869\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3\
        );

    \I__9042\ : Odrv4
    port map (
            O => \N__43866\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3\
        );

    \I__9041\ : InMux
    port map (
            O => \N__43857\,
            I => \N__43854\
        );

    \I__9040\ : LocalMux
    port map (
            O => \N__43854\,
            I => \N__43849\
        );

    \I__9039\ : InMux
    port map (
            O => \N__43853\,
            I => \N__43844\
        );

    \I__9038\ : InMux
    port map (
            O => \N__43852\,
            I => \N__43844\
        );

    \I__9037\ : Span4Mux_v
    port map (
            O => \N__43849\,
            I => \N__43841\
        );

    \I__9036\ : LocalMux
    port map (
            O => \N__43844\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_300_6\
        );

    \I__9035\ : Odrv4
    port map (
            O => \N__43841\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_300_6\
        );

    \I__9034\ : InMux
    port map (
            O => \N__43836\,
            I => \N__43833\
        );

    \I__9033\ : LocalMux
    port map (
            O => \N__43833\,
            I => \N__43830\
        );

    \I__9032\ : Span4Mux_v
    port map (
            O => \N__43830\,
            I => \N__43825\
        );

    \I__9031\ : InMux
    port map (
            O => \N__43829\,
            I => \N__43822\
        );

    \I__9030\ : InMux
    port map (
            O => \N__43828\,
            I => \N__43819\
        );

    \I__9029\ : Span4Mux_h
    port map (
            O => \N__43825\,
            I => \N__43814\
        );

    \I__9028\ : LocalMux
    port map (
            O => \N__43822\,
            I => \N__43814\
        );

    \I__9027\ : LocalMux
    port map (
            O => \N__43819\,
            I => \N__43810\
        );

    \I__9026\ : Span4Mux_h
    port map (
            O => \N__43814\,
            I => \N__43807\
        );

    \I__9025\ : InMux
    port map (
            O => \N__43813\,
            I => \N__43804\
        );

    \I__9024\ : Span4Mux_v
    port map (
            O => \N__43810\,
            I => \N__43799\
        );

    \I__9023\ : Span4Mux_v
    port map (
            O => \N__43807\,
            I => \N__43799\
        );

    \I__9022\ : LocalMux
    port map (
            O => \N__43804\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2\
        );

    \I__9021\ : Odrv4
    port map (
            O => \N__43799\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2\
        );

    \I__9020\ : InMux
    port map (
            O => \N__43794\,
            I => \N__43791\
        );

    \I__9019\ : LocalMux
    port map (
            O => \N__43791\,
            I => \N__43786\
        );

    \I__9018\ : InMux
    port map (
            O => \N__43790\,
            I => \N__43781\
        );

    \I__9017\ : InMux
    port map (
            O => \N__43789\,
            I => \N__43781\
        );

    \I__9016\ : Span4Mux_h
    port map (
            O => \N__43786\,
            I => \N__43778\
        );

    \I__9015\ : LocalMux
    port map (
            O => \N__43781\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1425_1\
        );

    \I__9014\ : Odrv4
    port map (
            O => \N__43778\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1425_1\
        );

    \I__9013\ : InMux
    port map (
            O => \N__43773\,
            I => \N__43770\
        );

    \I__9012\ : LocalMux
    port map (
            O => \N__43770\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_0\
        );

    \I__9011\ : InMux
    port map (
            O => \N__43767\,
            I => \N__43764\
        );

    \I__9010\ : LocalMux
    port map (
            O => \N__43764\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_1\
        );

    \I__9009\ : InMux
    port map (
            O => \N__43761\,
            I => \N__43758\
        );

    \I__9008\ : LocalMux
    port map (
            O => \N__43758\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_0\
        );

    \I__9007\ : InMux
    port map (
            O => \N__43755\,
            I => \N__43752\
        );

    \I__9006\ : LocalMux
    port map (
            O => \N__43752\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_1\
        );

    \I__9005\ : CascadeMux
    port map (
            O => \N__43749\,
            I => \N__43743\
        );

    \I__9004\ : CascadeMux
    port map (
            O => \N__43748\,
            I => \N__43740\
        );

    \I__9003\ : InMux
    port map (
            O => \N__43747\,
            I => \N__43734\
        );

    \I__9002\ : InMux
    port map (
            O => \N__43746\,
            I => \N__43734\
        );

    \I__9001\ : InMux
    port map (
            O => \N__43743\,
            I => \N__43728\
        );

    \I__9000\ : InMux
    port map (
            O => \N__43740\,
            I => \N__43728\
        );

    \I__8999\ : CEMux
    port map (
            O => \N__43739\,
            I => \N__43725\
        );

    \I__8998\ : LocalMux
    port map (
            O => \N__43734\,
            I => \N__43722\
        );

    \I__8997\ : CascadeMux
    port map (
            O => \N__43733\,
            I => \N__43717\
        );

    \I__8996\ : LocalMux
    port map (
            O => \N__43728\,
            I => \N__43712\
        );

    \I__8995\ : LocalMux
    port map (
            O => \N__43725\,
            I => \N__43712\
        );

    \I__8994\ : Span4Mux_h
    port map (
            O => \N__43722\,
            I => \N__43709\
        );

    \I__8993\ : InMux
    port map (
            O => \N__43721\,
            I => \N__43704\
        );

    \I__8992\ : InMux
    port map (
            O => \N__43720\,
            I => \N__43704\
        );

    \I__8991\ : InMux
    port map (
            O => \N__43717\,
            I => \N__43701\
        );

    \I__8990\ : Span4Mux_h
    port map (
            O => \N__43712\,
            I => \N__43698\
        );

    \I__8989\ : Span4Mux_h
    port map (
            O => \N__43709\,
            I => \N__43695\
        );

    \I__8988\ : LocalMux
    port map (
            O => \N__43704\,
            I => \I2C_top_level_inst1.s_load_addr0\
        );

    \I__8987\ : LocalMux
    port map (
            O => \N__43701\,
            I => \I2C_top_level_inst1.s_load_addr0\
        );

    \I__8986\ : Odrv4
    port map (
            O => \N__43698\,
            I => \I2C_top_level_inst1.s_load_addr0\
        );

    \I__8985\ : Odrv4
    port map (
            O => \N__43695\,
            I => \I2C_top_level_inst1.s_load_addr0\
        );

    \I__8984\ : CascadeMux
    port map (
            O => \N__43686\,
            I => \N__43683\
        );

    \I__8983\ : InMux
    port map (
            O => \N__43683\,
            I => \N__43680\
        );

    \I__8982\ : LocalMux
    port map (
            O => \N__43680\,
            I => \N__43677\
        );

    \I__8981\ : Span4Mux_h
    port map (
            O => \N__43677\,
            I => \N__43674\
        );

    \I__8980\ : Odrv4
    port map (
            O => \N__43674\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_6_0_0\
        );

    \I__8979\ : InMux
    port map (
            O => \N__43671\,
            I => \N__43666\
        );

    \I__8978\ : InMux
    port map (
            O => \N__43670\,
            I => \N__43659\
        );

    \I__8977\ : InMux
    port map (
            O => \N__43669\,
            I => \N__43659\
        );

    \I__8976\ : LocalMux
    port map (
            O => \N__43666\,
            I => \N__43656\
        );

    \I__8975\ : InMux
    port map (
            O => \N__43665\,
            I => \N__43651\
        );

    \I__8974\ : InMux
    port map (
            O => \N__43664\,
            I => \N__43651\
        );

    \I__8973\ : LocalMux
    port map (
            O => \N__43659\,
            I => \N__43648\
        );

    \I__8972\ : Span4Mux_h
    port map (
            O => \N__43656\,
            I => \N__43645\
        );

    \I__8971\ : LocalMux
    port map (
            O => \N__43651\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0\
        );

    \I__8970\ : Odrv12
    port map (
            O => \N__43648\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0\
        );

    \I__8969\ : Odrv4
    port map (
            O => \N__43645\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0\
        );

    \I__8968\ : CascadeMux
    port map (
            O => \N__43638\,
            I => \N__43635\
        );

    \I__8967\ : InMux
    port map (
            O => \N__43635\,
            I => \N__43632\
        );

    \I__8966\ : LocalMux
    port map (
            O => \N__43632\,
            I => \N__43629\
        );

    \I__8965\ : Odrv12
    port map (
            O => \N__43629\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1378\
        );

    \I__8964\ : CascadeMux
    port map (
            O => \N__43626\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_1676_cascade_\
        );

    \I__8963\ : InMux
    port map (
            O => \N__43623\,
            I => \N__43620\
        );

    \I__8962\ : LocalMux
    port map (
            O => \N__43620\,
            I => \N__43616\
        );

    \I__8961\ : InMux
    port map (
            O => \N__43619\,
            I => \N__43613\
        );

    \I__8960\ : Span4Mux_h
    port map (
            O => \N__43616\,
            I => \N__43609\
        );

    \I__8959\ : LocalMux
    port map (
            O => \N__43613\,
            I => \N__43606\
        );

    \I__8958\ : CascadeMux
    port map (
            O => \N__43612\,
            I => \N__43603\
        );

    \I__8957\ : Span4Mux_v
    port map (
            O => \N__43609\,
            I => \N__43600\
        );

    \I__8956\ : Span4Mux_h
    port map (
            O => \N__43606\,
            I => \N__43597\
        );

    \I__8955\ : InMux
    port map (
            O => \N__43603\,
            I => \N__43594\
        );

    \I__8954\ : Odrv4
    port map (
            O => \N__43600\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21\
        );

    \I__8953\ : Odrv4
    port map (
            O => \N__43597\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21\
        );

    \I__8952\ : LocalMux
    port map (
            O => \N__43594\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21\
        );

    \I__8951\ : CascadeMux
    port map (
            O => \N__43587\,
            I => \c_state_RNIEVJ7_22_cascade_\
        );

    \I__8950\ : InMux
    port map (
            O => \N__43584\,
            I => \N__43566\
        );

    \I__8949\ : CascadeMux
    port map (
            O => \N__43583\,
            I => \N__43563\
        );

    \I__8948\ : CascadeMux
    port map (
            O => \N__43582\,
            I => \N__43556\
        );

    \I__8947\ : CascadeMux
    port map (
            O => \N__43581\,
            I => \N__43553\
        );

    \I__8946\ : CascadeMux
    port map (
            O => \N__43580\,
            I => \N__43550\
        );

    \I__8945\ : CascadeMux
    port map (
            O => \N__43579\,
            I => \N__43546\
        );

    \I__8944\ : CascadeMux
    port map (
            O => \N__43578\,
            I => \N__43542\
        );

    \I__8943\ : InMux
    port map (
            O => \N__43577\,
            I => \N__43537\
        );

    \I__8942\ : CascadeMux
    port map (
            O => \N__43576\,
            I => \N__43534\
        );

    \I__8941\ : CascadeMux
    port map (
            O => \N__43575\,
            I => \N__43530\
        );

    \I__8940\ : CascadeMux
    port map (
            O => \N__43574\,
            I => \N__43526\
        );

    \I__8939\ : CascadeMux
    port map (
            O => \N__43573\,
            I => \N__43523\
        );

    \I__8938\ : CascadeMux
    port map (
            O => \N__43572\,
            I => \N__43520\
        );

    \I__8937\ : CascadeMux
    port map (
            O => \N__43571\,
            I => \N__43515\
        );

    \I__8936\ : InMux
    port map (
            O => \N__43570\,
            I => \N__43508\
        );

    \I__8935\ : CascadeMux
    port map (
            O => \N__43569\,
            I => \N__43505\
        );

    \I__8934\ : LocalMux
    port map (
            O => \N__43566\,
            I => \N__43502\
        );

    \I__8933\ : InMux
    port map (
            O => \N__43563\,
            I => \N__43499\
        );

    \I__8932\ : CascadeMux
    port map (
            O => \N__43562\,
            I => \N__43496\
        );

    \I__8931\ : CascadeMux
    port map (
            O => \N__43561\,
            I => \N__43493\
        );

    \I__8930\ : CascadeMux
    port map (
            O => \N__43560\,
            I => \N__43488\
        );

    \I__8929\ : CascadeMux
    port map (
            O => \N__43559\,
            I => \N__43484\
        );

    \I__8928\ : InMux
    port map (
            O => \N__43556\,
            I => \N__43481\
        );

    \I__8927\ : InMux
    port map (
            O => \N__43553\,
            I => \N__43478\
        );

    \I__8926\ : InMux
    port map (
            O => \N__43550\,
            I => \N__43463\
        );

    \I__8925\ : InMux
    port map (
            O => \N__43549\,
            I => \N__43463\
        );

    \I__8924\ : InMux
    port map (
            O => \N__43546\,
            I => \N__43463\
        );

    \I__8923\ : InMux
    port map (
            O => \N__43545\,
            I => \N__43463\
        );

    \I__8922\ : InMux
    port map (
            O => \N__43542\,
            I => \N__43463\
        );

    \I__8921\ : InMux
    port map (
            O => \N__43541\,
            I => \N__43463\
        );

    \I__8920\ : InMux
    port map (
            O => \N__43540\,
            I => \N__43463\
        );

    \I__8919\ : LocalMux
    port map (
            O => \N__43537\,
            I => \N__43460\
        );

    \I__8918\ : InMux
    port map (
            O => \N__43534\,
            I => \N__43455\
        );

    \I__8917\ : InMux
    port map (
            O => \N__43533\,
            I => \N__43455\
        );

    \I__8916\ : InMux
    port map (
            O => \N__43530\,
            I => \N__43452\
        );

    \I__8915\ : InMux
    port map (
            O => \N__43529\,
            I => \N__43437\
        );

    \I__8914\ : InMux
    port map (
            O => \N__43526\,
            I => \N__43437\
        );

    \I__8913\ : InMux
    port map (
            O => \N__43523\,
            I => \N__43437\
        );

    \I__8912\ : InMux
    port map (
            O => \N__43520\,
            I => \N__43437\
        );

    \I__8911\ : InMux
    port map (
            O => \N__43519\,
            I => \N__43437\
        );

    \I__8910\ : InMux
    port map (
            O => \N__43518\,
            I => \N__43437\
        );

    \I__8909\ : InMux
    port map (
            O => \N__43515\,
            I => \N__43437\
        );

    \I__8908\ : CascadeMux
    port map (
            O => \N__43514\,
            I => \N__43432\
        );

    \I__8907\ : InMux
    port map (
            O => \N__43513\,
            I => \N__43428\
        );

    \I__8906\ : InMux
    port map (
            O => \N__43512\,
            I => \N__43423\
        );

    \I__8905\ : InMux
    port map (
            O => \N__43511\,
            I => \N__43423\
        );

    \I__8904\ : LocalMux
    port map (
            O => \N__43508\,
            I => \N__43420\
        );

    \I__8903\ : InMux
    port map (
            O => \N__43505\,
            I => \N__43417\
        );

    \I__8902\ : Span4Mux_h
    port map (
            O => \N__43502\,
            I => \N__43412\
        );

    \I__8901\ : LocalMux
    port map (
            O => \N__43499\,
            I => \N__43412\
        );

    \I__8900\ : InMux
    port map (
            O => \N__43496\,
            I => \N__43397\
        );

    \I__8899\ : InMux
    port map (
            O => \N__43493\,
            I => \N__43397\
        );

    \I__8898\ : InMux
    port map (
            O => \N__43492\,
            I => \N__43397\
        );

    \I__8897\ : InMux
    port map (
            O => \N__43491\,
            I => \N__43397\
        );

    \I__8896\ : InMux
    port map (
            O => \N__43488\,
            I => \N__43397\
        );

    \I__8895\ : InMux
    port map (
            O => \N__43487\,
            I => \N__43397\
        );

    \I__8894\ : InMux
    port map (
            O => \N__43484\,
            I => \N__43397\
        );

    \I__8893\ : LocalMux
    port map (
            O => \N__43481\,
            I => \N__43392\
        );

    \I__8892\ : LocalMux
    port map (
            O => \N__43478\,
            I => \N__43392\
        );

    \I__8891\ : LocalMux
    port map (
            O => \N__43463\,
            I => \N__43389\
        );

    \I__8890\ : Span4Mux_h
    port map (
            O => \N__43460\,
            I => \N__43384\
        );

    \I__8889\ : LocalMux
    port map (
            O => \N__43455\,
            I => \N__43384\
        );

    \I__8888\ : LocalMux
    port map (
            O => \N__43452\,
            I => \N__43381\
        );

    \I__8887\ : LocalMux
    port map (
            O => \N__43437\,
            I => \N__43378\
        );

    \I__8886\ : InMux
    port map (
            O => \N__43436\,
            I => \N__43371\
        );

    \I__8885\ : InMux
    port map (
            O => \N__43435\,
            I => \N__43371\
        );

    \I__8884\ : InMux
    port map (
            O => \N__43432\,
            I => \N__43371\
        );

    \I__8883\ : CascadeMux
    port map (
            O => \N__43431\,
            I => \N__43367\
        );

    \I__8882\ : LocalMux
    port map (
            O => \N__43428\,
            I => \N__43362\
        );

    \I__8881\ : LocalMux
    port map (
            O => \N__43423\,
            I => \N__43359\
        );

    \I__8880\ : Span4Mux_v
    port map (
            O => \N__43420\,
            I => \N__43356\
        );

    \I__8879\ : LocalMux
    port map (
            O => \N__43417\,
            I => \N__43351\
        );

    \I__8878\ : Span4Mux_v
    port map (
            O => \N__43412\,
            I => \N__43351\
        );

    \I__8877\ : LocalMux
    port map (
            O => \N__43397\,
            I => \N__43342\
        );

    \I__8876\ : Span4Mux_v
    port map (
            O => \N__43392\,
            I => \N__43342\
        );

    \I__8875\ : Span4Mux_v
    port map (
            O => \N__43389\,
            I => \N__43342\
        );

    \I__8874\ : Span4Mux_v
    port map (
            O => \N__43384\,
            I => \N__43342\
        );

    \I__8873\ : Span4Mux_h
    port map (
            O => \N__43381\,
            I => \N__43335\
        );

    \I__8872\ : Span4Mux_v
    port map (
            O => \N__43378\,
            I => \N__43335\
        );

    \I__8871\ : LocalMux
    port map (
            O => \N__43371\,
            I => \N__43335\
        );

    \I__8870\ : InMux
    port map (
            O => \N__43370\,
            I => \N__43330\
        );

    \I__8869\ : InMux
    port map (
            O => \N__43367\,
            I => \N__43330\
        );

    \I__8868\ : InMux
    port map (
            O => \N__43366\,
            I => \N__43325\
        );

    \I__8867\ : InMux
    port map (
            O => \N__43365\,
            I => \N__43325\
        );

    \I__8866\ : Span12Mux_v
    port map (
            O => \N__43362\,
            I => \N__43322\
        );

    \I__8865\ : Span4Mux_v
    port map (
            O => \N__43359\,
            I => \N__43315\
        );

    \I__8864\ : Span4Mux_h
    port map (
            O => \N__43356\,
            I => \N__43315\
        );

    \I__8863\ : Span4Mux_v
    port map (
            O => \N__43351\,
            I => \N__43315\
        );

    \I__8862\ : Span4Mux_h
    port map (
            O => \N__43342\,
            I => \N__43310\
        );

    \I__8861\ : Span4Mux_v
    port map (
            O => \N__43335\,
            I => \N__43310\
        );

    \I__8860\ : LocalMux
    port map (
            O => \N__43330\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\
        );

    \I__8859\ : LocalMux
    port map (
            O => \N__43325\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\
        );

    \I__8858\ : Odrv12
    port map (
            O => \N__43322\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\
        );

    \I__8857\ : Odrv4
    port map (
            O => \N__43315\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\
        );

    \I__8856\ : Odrv4
    port map (
            O => \N__43310\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\
        );

    \I__8855\ : CascadeMux
    port map (
            O => \N__43299\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_77_cascade_\
        );

    \I__8854\ : IoInMux
    port map (
            O => \N__43296\,
            I => \N__43293\
        );

    \I__8853\ : LocalMux
    port map (
            O => \N__43293\,
            I => \N__43290\
        );

    \I__8852\ : Span4Mux_s1_h
    port map (
            O => \N__43290\,
            I => \N__43287\
        );

    \I__8851\ : Span4Mux_v
    port map (
            O => \N__43287\,
            I => \N__43284\
        );

    \I__8850\ : Span4Mux_h
    port map (
            O => \N__43284\,
            I => \N__43281\
        );

    \I__8849\ : Span4Mux_h
    port map (
            O => \N__43281\,
            I => \N__43278\
        );

    \I__8848\ : Odrv4
    port map (
            O => \N__43278\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0\
        );

    \I__8847\ : InMux
    port map (
            O => \N__43275\,
            I => \N__43272\
        );

    \I__8846\ : LocalMux
    port map (
            O => \N__43272\,
            I => \N__43269\
        );

    \I__8845\ : Span4Mux_v
    port map (
            O => \N__43269\,
            I => \N__43265\
        );

    \I__8844\ : InMux
    port map (
            O => \N__43268\,
            I => \N__43262\
        );

    \I__8843\ : Odrv4
    port map (
            O => \N__43265\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13\
        );

    \I__8842\ : LocalMux
    port map (
            O => \N__43262\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13\
        );

    \I__8841\ : InMux
    port map (
            O => \N__43257\,
            I => \N__43254\
        );

    \I__8840\ : LocalMux
    port map (
            O => \N__43254\,
            I => \N__43251\
        );

    \I__8839\ : Span4Mux_v
    port map (
            O => \N__43251\,
            I => \N__43248\
        );

    \I__8838\ : Odrv4
    port map (
            O => \N__43248\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_13\
        );

    \I__8837\ : InMux
    port map (
            O => \N__43245\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12\
        );

    \I__8836\ : InMux
    port map (
            O => \N__43242\,
            I => \N__43239\
        );

    \I__8835\ : LocalMux
    port map (
            O => \N__43239\,
            I => \N__43236\
        );

    \I__8834\ : Span4Mux_v
    port map (
            O => \N__43236\,
            I => \N__43232\
        );

    \I__8833\ : InMux
    port map (
            O => \N__43235\,
            I => \N__43229\
        );

    \I__8832\ : Odrv4
    port map (
            O => \N__43232\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14\
        );

    \I__8831\ : LocalMux
    port map (
            O => \N__43229\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14\
        );

    \I__8830\ : InMux
    port map (
            O => \N__43224\,
            I => \N__43221\
        );

    \I__8829\ : LocalMux
    port map (
            O => \N__43221\,
            I => \N__43218\
        );

    \I__8828\ : Span4Mux_h
    port map (
            O => \N__43218\,
            I => \N__43215\
        );

    \I__8827\ : Odrv4
    port map (
            O => \N__43215\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_14\
        );

    \I__8826\ : InMux
    port map (
            O => \N__43212\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13\
        );

    \I__8825\ : InMux
    port map (
            O => \N__43209\,
            I => \N__43206\
        );

    \I__8824\ : LocalMux
    port map (
            O => \N__43206\,
            I => \N__43202\
        );

    \I__8823\ : CascadeMux
    port map (
            O => \N__43205\,
            I => \N__43199\
        );

    \I__8822\ : Span4Mux_h
    port map (
            O => \N__43202\,
            I => \N__43196\
        );

    \I__8821\ : InMux
    port map (
            O => \N__43199\,
            I => \N__43193\
        );

    \I__8820\ : Odrv4
    port map (
            O => \N__43196\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15\
        );

    \I__8819\ : LocalMux
    port map (
            O => \N__43193\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15\
        );

    \I__8818\ : InMux
    port map (
            O => \N__43188\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_14\
        );

    \I__8817\ : InMux
    port map (
            O => \N__43185\,
            I => \N__43182\
        );

    \I__8816\ : LocalMux
    port map (
            O => \N__43182\,
            I => \N__43179\
        );

    \I__8815\ : Span4Mux_h
    port map (
            O => \N__43179\,
            I => \N__43176\
        );

    \I__8814\ : Odrv4
    port map (
            O => \N__43176\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_15\
        );

    \I__8813\ : InMux
    port map (
            O => \N__43173\,
            I => \N__43170\
        );

    \I__8812\ : LocalMux
    port map (
            O => \N__43170\,
            I => \N__43167\
        );

    \I__8811\ : Span4Mux_h
    port map (
            O => \N__43167\,
            I => \N__43164\
        );

    \I__8810\ : Span4Mux_v
    port map (
            O => \N__43164\,
            I => \N__43161\
        );

    \I__8809\ : Odrv4
    port map (
            O => \N__43161\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_103_0\
        );

    \I__8808\ : InMux
    port map (
            O => \N__43158\,
            I => \N__43155\
        );

    \I__8807\ : LocalMux
    port map (
            O => \N__43155\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_1\
        );

    \I__8806\ : InMux
    port map (
            O => \N__43152\,
            I => \N__43149\
        );

    \I__8805\ : LocalMux
    port map (
            O => \N__43149\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_0\
        );

    \I__8804\ : InMux
    port map (
            O => \N__43146\,
            I => \N__43143\
        );

    \I__8803\ : LocalMux
    port map (
            O => \N__43143\,
            I => \N__43139\
        );

    \I__8802\ : CascadeMux
    port map (
            O => \N__43142\,
            I => \N__43136\
        );

    \I__8801\ : Span4Mux_h
    port map (
            O => \N__43139\,
            I => \N__43131\
        );

    \I__8800\ : InMux
    port map (
            O => \N__43136\,
            I => \N__43124\
        );

    \I__8799\ : InMux
    port map (
            O => \N__43135\,
            I => \N__43124\
        );

    \I__8798\ : InMux
    port map (
            O => \N__43134\,
            I => \N__43124\
        );

    \I__8797\ : Odrv4
    port map (
            O => \N__43131\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5\
        );

    \I__8796\ : LocalMux
    port map (
            O => \N__43124\,
            I => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5\
        );

    \I__8795\ : CascadeMux
    port map (
            O => \N__43119\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_291_cascade_\
        );

    \I__8794\ : InMux
    port map (
            O => \N__43116\,
            I => \N__43113\
        );

    \I__8793\ : LocalMux
    port map (
            O => \N__43113\,
            I => \N__43110\
        );

    \I__8792\ : Span4Mux_h
    port map (
            O => \N__43110\,
            I => \N__43107\
        );

    \I__8791\ : Odrv4
    port map (
            O => \N__43107\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_5\
        );

    \I__8790\ : InMux
    port map (
            O => \N__43104\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4\
        );

    \I__8789\ : InMux
    port map (
            O => \N__43101\,
            I => \N__43098\
        );

    \I__8788\ : LocalMux
    port map (
            O => \N__43098\,
            I => \N__43095\
        );

    \I__8787\ : Span4Mux_h
    port map (
            O => \N__43095\,
            I => \N__43092\
        );

    \I__8786\ : Odrv4
    port map (
            O => \N__43092\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_6\
        );

    \I__8785\ : InMux
    port map (
            O => \N__43089\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5\
        );

    \I__8784\ : InMux
    port map (
            O => \N__43086\,
            I => \N__43083\
        );

    \I__8783\ : LocalMux
    port map (
            O => \N__43083\,
            I => \N__43080\
        );

    \I__8782\ : Span4Mux_h
    port map (
            O => \N__43080\,
            I => \N__43077\
        );

    \I__8781\ : Odrv4
    port map (
            O => \N__43077\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_7\
        );

    \I__8780\ : InMux
    port map (
            O => \N__43074\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6\
        );

    \I__8779\ : InMux
    port map (
            O => \N__43071\,
            I => \bfn_20_18_0_\
        );

    \I__8778\ : InMux
    port map (
            O => \N__43068\,
            I => \N__43065\
        );

    \I__8777\ : LocalMux
    port map (
            O => \N__43065\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_9\
        );

    \I__8776\ : InMux
    port map (
            O => \N__43062\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8\
        );

    \I__8775\ : InMux
    port map (
            O => \N__43059\,
            I => \N__43056\
        );

    \I__8774\ : LocalMux
    port map (
            O => \N__43056\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_10\
        );

    \I__8773\ : InMux
    port map (
            O => \N__43053\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9\
        );

    \I__8772\ : InMux
    port map (
            O => \N__43050\,
            I => \N__43047\
        );

    \I__8771\ : LocalMux
    port map (
            O => \N__43047\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_11\
        );

    \I__8770\ : InMux
    port map (
            O => \N__43044\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10\
        );

    \I__8769\ : InMux
    port map (
            O => \N__43041\,
            I => \N__43038\
        );

    \I__8768\ : LocalMux
    port map (
            O => \N__43038\,
            I => \N__43035\
        );

    \I__8767\ : Span4Mux_h
    port map (
            O => \N__43035\,
            I => \N__43031\
        );

    \I__8766\ : InMux
    port map (
            O => \N__43034\,
            I => \N__43028\
        );

    \I__8765\ : Odrv4
    port map (
            O => \N__43031\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12\
        );

    \I__8764\ : LocalMux
    port map (
            O => \N__43028\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12\
        );

    \I__8763\ : InMux
    port map (
            O => \N__43023\,
            I => \N__43020\
        );

    \I__8762\ : LocalMux
    port map (
            O => \N__43020\,
            I => \N__43017\
        );

    \I__8761\ : Span4Mux_v
    port map (
            O => \N__43017\,
            I => \N__43014\
        );

    \I__8760\ : Span4Mux_h
    port map (
            O => \N__43014\,
            I => \N__43011\
        );

    \I__8759\ : Odrv4
    port map (
            O => \N__43011\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_12\
        );

    \I__8758\ : InMux
    port map (
            O => \N__43008\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11\
        );

    \I__8757\ : InMux
    port map (
            O => \N__43005\,
            I => \N__43000\
        );

    \I__8756\ : CascadeMux
    port map (
            O => \N__43004\,
            I => \N__42997\
        );

    \I__8755\ : CascadeMux
    port map (
            O => \N__43003\,
            I => \N__42994\
        );

    \I__8754\ : LocalMux
    port map (
            O => \N__43000\,
            I => \N__42991\
        );

    \I__8753\ : InMux
    port map (
            O => \N__42997\,
            I => \N__42986\
        );

    \I__8752\ : InMux
    port map (
            O => \N__42994\,
            I => \N__42986\
        );

    \I__8751\ : Span12Mux_h
    port map (
            O => \N__42991\,
            I => \N__42983\
        );

    \I__8750\ : LocalMux
    port map (
            O => \N__42986\,
            I => \N__42980\
        );

    \I__8749\ : Odrv12
    port map (
            O => \N__42983\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_2
        );

    \I__8748\ : Odrv4
    port map (
            O => \N__42980\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_2
        );

    \I__8747\ : InMux
    port map (
            O => \N__42975\,
            I => \N__42972\
        );

    \I__8746\ : LocalMux
    port map (
            O => \N__42972\,
            I => \N__42969\
        );

    \I__8745\ : Span4Mux_v
    port map (
            O => \N__42969\,
            I => \N__42966\
        );

    \I__8744\ : Span4Mux_v
    port map (
            O => \N__42966\,
            I => \N__42961\
        );

    \I__8743\ : InMux
    port map (
            O => \N__42965\,
            I => \N__42956\
        );

    \I__8742\ : InMux
    port map (
            O => \N__42964\,
            I => \N__42956\
        );

    \I__8741\ : Odrv4
    port map (
            O => \N__42961\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_2
        );

    \I__8740\ : LocalMux
    port map (
            O => \N__42956\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_2
        );

    \I__8739\ : InMux
    port map (
            O => \N__42951\,
            I => \N__42948\
        );

    \I__8738\ : LocalMux
    port map (
            O => \N__42948\,
            I => \N__42945\
        );

    \I__8737\ : Span4Mux_h
    port map (
            O => \N__42945\,
            I => \N__42941\
        );

    \I__8736\ : CascadeMux
    port map (
            O => \N__42944\,
            I => \N__42937\
        );

    \I__8735\ : Span4Mux_v
    port map (
            O => \N__42941\,
            I => \N__42934\
        );

    \I__8734\ : InMux
    port map (
            O => \N__42940\,
            I => \N__42931\
        );

    \I__8733\ : InMux
    port map (
            O => \N__42937\,
            I => \N__42928\
        );

    \I__8732\ : Odrv4
    port map (
            O => \N__42934\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_11
        );

    \I__8731\ : LocalMux
    port map (
            O => \N__42931\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_11
        );

    \I__8730\ : LocalMux
    port map (
            O => \N__42928\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_11
        );

    \I__8729\ : InMux
    port map (
            O => \N__42921\,
            I => \N__42918\
        );

    \I__8728\ : LocalMux
    port map (
            O => \N__42918\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_11\
        );

    \I__8727\ : InMux
    port map (
            O => \N__42915\,
            I => \N__42912\
        );

    \I__8726\ : LocalMux
    port map (
            O => \N__42912\,
            I => \N__42909\
        );

    \I__8725\ : Span4Mux_v
    port map (
            O => \N__42909\,
            I => \N__42906\
        );

    \I__8724\ : Span4Mux_h
    port map (
            O => \N__42906\,
            I => \N__42901\
        );

    \I__8723\ : InMux
    port map (
            O => \N__42905\,
            I => \N__42898\
        );

    \I__8722\ : InMux
    port map (
            O => \N__42904\,
            I => \N__42895\
        );

    \I__8721\ : Odrv4
    port map (
            O => \N__42901\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_11
        );

    \I__8720\ : LocalMux
    port map (
            O => \N__42898\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_11
        );

    \I__8719\ : LocalMux
    port map (
            O => \N__42895\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_11
        );

    \I__8718\ : InMux
    port map (
            O => \N__42888\,
            I => \N__42885\
        );

    \I__8717\ : LocalMux
    port map (
            O => \N__42885\,
            I => \N__42882\
        );

    \I__8716\ : Span4Mux_h
    port map (
            O => \N__42882\,
            I => \N__42879\
        );

    \I__8715\ : Span4Mux_v
    port map (
            O => \N__42879\,
            I => \N__42876\
        );

    \I__8714\ : Odrv4
    port map (
            O => \N__42876\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_1\
        );

    \I__8713\ : InMux
    port map (
            O => \N__42873\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0\
        );

    \I__8712\ : InMux
    port map (
            O => \N__42870\,
            I => \N__42867\
        );

    \I__8711\ : LocalMux
    port map (
            O => \N__42867\,
            I => \N__42864\
        );

    \I__8710\ : Span4Mux_v
    port map (
            O => \N__42864\,
            I => \N__42861\
        );

    \I__8709\ : Span4Mux_v
    port map (
            O => \N__42861\,
            I => \N__42858\
        );

    \I__8708\ : Odrv4
    port map (
            O => \N__42858\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_2\
        );

    \I__8707\ : InMux
    port map (
            O => \N__42855\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1\
        );

    \I__8706\ : InMux
    port map (
            O => \N__42852\,
            I => \N__42849\
        );

    \I__8705\ : LocalMux
    port map (
            O => \N__42849\,
            I => \N__42846\
        );

    \I__8704\ : Span4Mux_v
    port map (
            O => \N__42846\,
            I => \N__42843\
        );

    \I__8703\ : Odrv4
    port map (
            O => \N__42843\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_CO\
        );

    \I__8702\ : InMux
    port map (
            O => \N__42840\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2\
        );

    \I__8701\ : InMux
    port map (
            O => \N__42837\,
            I => \N__42834\
        );

    \I__8700\ : LocalMux
    port map (
            O => \N__42834\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_4\
        );

    \I__8699\ : InMux
    port map (
            O => \N__42831\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3\
        );

    \I__8698\ : CascadeMux
    port map (
            O => \N__42828\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238DZ0Z7_cascade_\
        );

    \I__8697\ : InMux
    port map (
            O => \N__42825\,
            I => \N__42822\
        );

    \I__8696\ : LocalMux
    port map (
            O => \N__42822\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_11\
        );

    \I__8695\ : InMux
    port map (
            O => \N__42819\,
            I => \N__42816\
        );

    \I__8694\ : LocalMux
    port map (
            O => \N__42816\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_13\
        );

    \I__8693\ : InMux
    port map (
            O => \N__42813\,
            I => \N__42809\
        );

    \I__8692\ : InMux
    port map (
            O => \N__42812\,
            I => \N__42806\
        );

    \I__8691\ : LocalMux
    port map (
            O => \N__42809\,
            I => \N__42803\
        );

    \I__8690\ : LocalMux
    port map (
            O => \N__42806\,
            I => \N__42800\
        );

    \I__8689\ : Span4Mux_h
    port map (
            O => \N__42803\,
            I => \N__42797\
        );

    \I__8688\ : Span4Mux_h
    port map (
            O => \N__42800\,
            I => \N__42794\
        );

    \I__8687\ : Span4Mux_v
    port map (
            O => \N__42797\,
            I => \N__42790\
        );

    \I__8686\ : Span4Mux_h
    port map (
            O => \N__42794\,
            I => \N__42787\
        );

    \I__8685\ : InMux
    port map (
            O => \N__42793\,
            I => \N__42784\
        );

    \I__8684\ : Odrv4
    port map (
            O => \N__42790\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_13
        );

    \I__8683\ : Odrv4
    port map (
            O => \N__42787\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_13
        );

    \I__8682\ : LocalMux
    port map (
            O => \N__42784\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_13
        );

    \I__8681\ : InMux
    port map (
            O => \N__42777\,
            I => \N__42774\
        );

    \I__8680\ : LocalMux
    port map (
            O => \N__42774\,
            I => \N__42771\
        );

    \I__8679\ : Span4Mux_h
    port map (
            O => \N__42771\,
            I => \N__42768\
        );

    \I__8678\ : Odrv4
    port map (
            O => \N__42768\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_23\
        );

    \I__8677\ : InMux
    port map (
            O => \N__42765\,
            I => \N__42762\
        );

    \I__8676\ : LocalMux
    port map (
            O => \N__42762\,
            I => \N__42759\
        );

    \I__8675\ : Span4Mux_h
    port map (
            O => \N__42759\,
            I => \N__42755\
        );

    \I__8674\ : CascadeMux
    port map (
            O => \N__42758\,
            I => \N__42752\
        );

    \I__8673\ : Span4Mux_v
    port map (
            O => \N__42755\,
            I => \N__42748\
        );

    \I__8672\ : InMux
    port map (
            O => \N__42752\,
            I => \N__42743\
        );

    \I__8671\ : InMux
    port map (
            O => \N__42751\,
            I => \N__42743\
        );

    \I__8670\ : Odrv4
    port map (
            O => \N__42748\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_10
        );

    \I__8669\ : LocalMux
    port map (
            O => \N__42743\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_10
        );

    \I__8668\ : InMux
    port map (
            O => \N__42738\,
            I => \N__42735\
        );

    \I__8667\ : LocalMux
    port map (
            O => \N__42735\,
            I => \N__42732\
        );

    \I__8666\ : Span4Mux_v
    port map (
            O => \N__42732\,
            I => \N__42729\
        );

    \I__8665\ : Span4Mux_h
    port map (
            O => \N__42729\,
            I => \N__42725\
        );

    \I__8664\ : CascadeMux
    port map (
            O => \N__42728\,
            I => \N__42721\
        );

    \I__8663\ : Span4Mux_v
    port map (
            O => \N__42725\,
            I => \N__42718\
        );

    \I__8662\ : InMux
    port map (
            O => \N__42724\,
            I => \N__42715\
        );

    \I__8661\ : InMux
    port map (
            O => \N__42721\,
            I => \N__42712\
        );

    \I__8660\ : Odrv4
    port map (
            O => \N__42718\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_10
        );

    \I__8659\ : LocalMux
    port map (
            O => \N__42715\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_10
        );

    \I__8658\ : LocalMux
    port map (
            O => \N__42712\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_10
        );

    \I__8657\ : InMux
    port map (
            O => \N__42705\,
            I => \N__42702\
        );

    \I__8656\ : LocalMux
    port map (
            O => \N__42702\,
            I => \N__42698\
        );

    \I__8655\ : CascadeMux
    port map (
            O => \N__42701\,
            I => \N__42694\
        );

    \I__8654\ : Span4Mux_h
    port map (
            O => \N__42698\,
            I => \N__42691\
        );

    \I__8653\ : InMux
    port map (
            O => \N__42697\,
            I => \N__42686\
        );

    \I__8652\ : InMux
    port map (
            O => \N__42694\,
            I => \N__42686\
        );

    \I__8651\ : Odrv4
    port map (
            O => \N__42691\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_12
        );

    \I__8650\ : LocalMux
    port map (
            O => \N__42686\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_12
        );

    \I__8649\ : InMux
    port map (
            O => \N__42681\,
            I => \N__42678\
        );

    \I__8648\ : LocalMux
    port map (
            O => \N__42678\,
            I => \N__42675\
        );

    \I__8647\ : Span4Mux_v
    port map (
            O => \N__42675\,
            I => \N__42671\
        );

    \I__8646\ : CascadeMux
    port map (
            O => \N__42674\,
            I => \N__42667\
        );

    \I__8645\ : Span4Mux_v
    port map (
            O => \N__42671\,
            I => \N__42664\
        );

    \I__8644\ : InMux
    port map (
            O => \N__42670\,
            I => \N__42661\
        );

    \I__8643\ : InMux
    port map (
            O => \N__42667\,
            I => \N__42658\
        );

    \I__8642\ : Span4Mux_h
    port map (
            O => \N__42664\,
            I => \N__42655\
        );

    \I__8641\ : LocalMux
    port map (
            O => \N__42661\,
            I => \N__42650\
        );

    \I__8640\ : LocalMux
    port map (
            O => \N__42658\,
            I => \N__42650\
        );

    \I__8639\ : Odrv4
    port map (
            O => \N__42655\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_22
        );

    \I__8638\ : Odrv4
    port map (
            O => \N__42650\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_22
        );

    \I__8637\ : CascadeMux
    port map (
            O => \N__42645\,
            I => \N__42640\
        );

    \I__8636\ : CascadeMux
    port map (
            O => \N__42644\,
            I => \N__42637\
        );

    \I__8635\ : InMux
    port map (
            O => \N__42643\,
            I => \N__42634\
        );

    \I__8634\ : InMux
    port map (
            O => \N__42640\,
            I => \N__42629\
        );

    \I__8633\ : InMux
    port map (
            O => \N__42637\,
            I => \N__42629\
        );

    \I__8632\ : LocalMux
    port map (
            O => \N__42634\,
            I => \N__42626\
        );

    \I__8631\ : LocalMux
    port map (
            O => \N__42629\,
            I => \N__42623\
        );

    \I__8630\ : Span4Mux_h
    port map (
            O => \N__42626\,
            I => \N__42620\
        );

    \I__8629\ : Span4Mux_h
    port map (
            O => \N__42623\,
            I => \N__42617\
        );

    \I__8628\ : Odrv4
    port map (
            O => \N__42620\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_14
        );

    \I__8627\ : Odrv4
    port map (
            O => \N__42617\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_14
        );

    \I__8626\ : InMux
    port map (
            O => \N__42612\,
            I => \N__42609\
        );

    \I__8625\ : LocalMux
    port map (
            O => \N__42609\,
            I => \N__42605\
        );

    \I__8624\ : CascadeMux
    port map (
            O => \N__42608\,
            I => \N__42601\
        );

    \I__8623\ : Span4Mux_h
    port map (
            O => \N__42605\,
            I => \N__42598\
        );

    \I__8622\ : InMux
    port map (
            O => \N__42604\,
            I => \N__42593\
        );

    \I__8621\ : InMux
    port map (
            O => \N__42601\,
            I => \N__42593\
        );

    \I__8620\ : Span4Mux_v
    port map (
            O => \N__42598\,
            I => \N__42590\
        );

    \I__8619\ : LocalMux
    port map (
            O => \N__42593\,
            I => \N__42587\
        );

    \I__8618\ : Odrv4
    port map (
            O => \N__42590\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_15
        );

    \I__8617\ : Odrv4
    port map (
            O => \N__42587\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_15
        );

    \I__8616\ : InMux
    port map (
            O => \N__42582\,
            I => \N__42579\
        );

    \I__8615\ : LocalMux
    port map (
            O => \N__42579\,
            I => \N__42574\
        );

    \I__8614\ : InMux
    port map (
            O => \N__42578\,
            I => \N__42569\
        );

    \I__8613\ : InMux
    port map (
            O => \N__42577\,
            I => \N__42569\
        );

    \I__8612\ : Span12Mux_v
    port map (
            O => \N__42574\,
            I => \N__42566\
        );

    \I__8611\ : LocalMux
    port map (
            O => \N__42569\,
            I => \N__42563\
        );

    \I__8610\ : Odrv12
    port map (
            O => \N__42566\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_16
        );

    \I__8609\ : Odrv4
    port map (
            O => \N__42563\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_16
        );

    \I__8608\ : InMux
    port map (
            O => \N__42558\,
            I => \N__42555\
        );

    \I__8607\ : LocalMux
    port map (
            O => \N__42555\,
            I => \N__42551\
        );

    \I__8606\ : InMux
    port map (
            O => \N__42554\,
            I => \N__42547\
        );

    \I__8605\ : Span4Mux_v
    port map (
            O => \N__42551\,
            I => \N__42544\
        );

    \I__8604\ : InMux
    port map (
            O => \N__42550\,
            I => \N__42541\
        );

    \I__8603\ : LocalMux
    port map (
            O => \N__42547\,
            I => \N__42538\
        );

    \I__8602\ : Span4Mux_h
    port map (
            O => \N__42544\,
            I => \N__42531\
        );

    \I__8601\ : LocalMux
    port map (
            O => \N__42541\,
            I => \N__42531\
        );

    \I__8600\ : Span4Mux_v
    port map (
            O => \N__42538\,
            I => \N__42531\
        );

    \I__8599\ : Odrv4
    port map (
            O => \N__42531\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_11
        );

    \I__8598\ : CascadeMux
    port map (
            O => \N__42528\,
            I => \N__42524\
        );

    \I__8597\ : InMux
    port map (
            O => \N__42527\,
            I => \N__42521\
        );

    \I__8596\ : InMux
    port map (
            O => \N__42524\,
            I => \N__42518\
        );

    \I__8595\ : LocalMux
    port map (
            O => \N__42521\,
            I => \N__42515\
        );

    \I__8594\ : LocalMux
    port map (
            O => \N__42518\,
            I => \N__42511\
        );

    \I__8593\ : Span4Mux_h
    port map (
            O => \N__42515\,
            I => \N__42508\
        );

    \I__8592\ : InMux
    port map (
            O => \N__42514\,
            I => \N__42505\
        );

    \I__8591\ : Span4Mux_v
    port map (
            O => \N__42511\,
            I => \N__42502\
        );

    \I__8590\ : Span4Mux_v
    port map (
            O => \N__42508\,
            I => \N__42497\
        );

    \I__8589\ : LocalMux
    port map (
            O => \N__42505\,
            I => \N__42497\
        );

    \I__8588\ : Span4Mux_h
    port map (
            O => \N__42502\,
            I => \N__42494\
        );

    \I__8587\ : Odrv4
    port map (
            O => \N__42497\,
            I => cemf_module_64ch_ctrl_inst1_data_config_11
        );

    \I__8586\ : Odrv4
    port map (
            O => \N__42494\,
            I => cemf_module_64ch_ctrl_inst1_data_config_11
        );

    \I__8585\ : CascadeMux
    port map (
            O => \N__42489\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_11_cascade_\
        );

    \I__8584\ : InMux
    port map (
            O => \N__42486\,
            I => \N__42483\
        );

    \I__8583\ : LocalMux
    port map (
            O => \N__42483\,
            I => \N__42478\
        );

    \I__8582\ : InMux
    port map (
            O => \N__42482\,
            I => \N__42475\
        );

    \I__8581\ : CascadeMux
    port map (
            O => \N__42481\,
            I => \N__42472\
        );

    \I__8580\ : Span4Mux_v
    port map (
            O => \N__42478\,
            I => \N__42467\
        );

    \I__8579\ : LocalMux
    port map (
            O => \N__42475\,
            I => \N__42467\
        );

    \I__8578\ : InMux
    port map (
            O => \N__42472\,
            I => \N__42464\
        );

    \I__8577\ : Span4Mux_h
    port map (
            O => \N__42467\,
            I => \N__42461\
        );

    \I__8576\ : LocalMux
    port map (
            O => \N__42464\,
            I => \N__42458\
        );

    \I__8575\ : Span4Mux_h
    port map (
            O => \N__42461\,
            I => \N__42455\
        );

    \I__8574\ : Span12Mux_v
    port map (
            O => \N__42458\,
            I => \N__42452\
        );

    \I__8573\ : Odrv4
    port map (
            O => \N__42455\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_4
        );

    \I__8572\ : Odrv12
    port map (
            O => \N__42452\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_4
        );

    \I__8571\ : InMux
    port map (
            O => \N__42447\,
            I => \N__42440\
        );

    \I__8570\ : InMux
    port map (
            O => \N__42446\,
            I => \N__42440\
        );

    \I__8569\ : CascadeMux
    port map (
            O => \N__42445\,
            I => \N__42437\
        );

    \I__8568\ : LocalMux
    port map (
            O => \N__42440\,
            I => \N__42434\
        );

    \I__8567\ : InMux
    port map (
            O => \N__42437\,
            I => \N__42431\
        );

    \I__8566\ : Span4Mux_h
    port map (
            O => \N__42434\,
            I => \N__42428\
        );

    \I__8565\ : LocalMux
    port map (
            O => \N__42431\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_20
        );

    \I__8564\ : Odrv4
    port map (
            O => \N__42428\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_20
        );

    \I__8563\ : InMux
    port map (
            O => \N__42423\,
            I => \N__42420\
        );

    \I__8562\ : LocalMux
    port map (
            O => \N__42420\,
            I => \N__42416\
        );

    \I__8561\ : CascadeMux
    port map (
            O => \N__42419\,
            I => \N__42413\
        );

    \I__8560\ : Span4Mux_v
    port map (
            O => \N__42416\,
            I => \N__42409\
        );

    \I__8559\ : InMux
    port map (
            O => \N__42413\,
            I => \N__42404\
        );

    \I__8558\ : InMux
    port map (
            O => \N__42412\,
            I => \N__42404\
        );

    \I__8557\ : Sp12to4
    port map (
            O => \N__42409\,
            I => \N__42399\
        );

    \I__8556\ : LocalMux
    port map (
            O => \N__42404\,
            I => \N__42399\
        );

    \I__8555\ : Odrv12
    port map (
            O => \N__42399\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_20
        );

    \I__8554\ : InMux
    port map (
            O => \N__42396\,
            I => \N__42393\
        );

    \I__8553\ : LocalMux
    port map (
            O => \N__42393\,
            I => \N__42390\
        );

    \I__8552\ : Odrv12
    port map (
            O => \N__42390\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_15\
        );

    \I__8551\ : CascadeMux
    port map (
            O => \N__42387\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_15_cascade_\
        );

    \I__8550\ : CascadeMux
    port map (
            O => \N__42384\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8DZ0Z7_cascade_\
        );

    \I__8549\ : InMux
    port map (
            O => \N__42381\,
            I => \N__42378\
        );

    \I__8548\ : LocalMux
    port map (
            O => \N__42378\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15\
        );

    \I__8547\ : InMux
    port map (
            O => \N__42375\,
            I => \N__42372\
        );

    \I__8546\ : LocalMux
    port map (
            O => \N__42372\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_14\
        );

    \I__8545\ : CascadeMux
    port map (
            O => \N__42369\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15_cascade_\
        );

    \I__8544\ : CascadeMux
    port map (
            O => \N__42366\,
            I => \N__42363\
        );

    \I__8543\ : InMux
    port map (
            O => \N__42363\,
            I => \N__42360\
        );

    \I__8542\ : LocalMux
    port map (
            O => \N__42360\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_16\
        );

    \I__8541\ : CascadeMux
    port map (
            O => \N__42357\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8DZ0Z7_cascade_\
        );

    \I__8540\ : InMux
    port map (
            O => \N__42354\,
            I => \N__42351\
        );

    \I__8539\ : LocalMux
    port map (
            O => \N__42351\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16\
        );

    \I__8538\ : CascadeMux
    port map (
            O => \N__42348\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16_cascade_\
        );

    \I__8537\ : InMux
    port map (
            O => \N__42345\,
            I => \N__42342\
        );

    \I__8536\ : LocalMux
    port map (
            O => \N__42342\,
            I => \N__42339\
        );

    \I__8535\ : Odrv4
    port map (
            O => \N__42339\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_15\
        );

    \I__8534\ : InMux
    port map (
            O => \N__42336\,
            I => \N__42333\
        );

    \I__8533\ : LocalMux
    port map (
            O => \N__42333\,
            I => \N__42330\
        );

    \I__8532\ : Odrv12
    port map (
            O => \N__42330\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_16\
        );

    \I__8531\ : InMux
    port map (
            O => \N__42327\,
            I => \N__42324\
        );

    \I__8530\ : LocalMux
    port map (
            O => \N__42324\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_16\
        );

    \I__8529\ : CascadeMux
    port map (
            O => \N__42321\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_16_cascade_\
        );

    \I__8528\ : InMux
    port map (
            O => \N__42318\,
            I => \N__42315\
        );

    \I__8527\ : LocalMux
    port map (
            O => \N__42315\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_16\
        );

    \I__8526\ : InMux
    port map (
            O => \N__42312\,
            I => \N__42309\
        );

    \I__8525\ : LocalMux
    port map (
            O => \N__42309\,
            I => \N__42306\
        );

    \I__8524\ : Span4Mux_h
    port map (
            O => \N__42306\,
            I => \N__42303\
        );

    \I__8523\ : Span4Mux_h
    port map (
            O => \N__42303\,
            I => \N__42300\
        );

    \I__8522\ : Span4Mux_v
    port map (
            O => \N__42300\,
            I => \N__42297\
        );

    \I__8521\ : Span4Mux_h
    port map (
            O => \N__42297\,
            I => \N__42294\
        );

    \I__8520\ : Odrv4
    port map (
            O => \N__42294\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_24
        );

    \I__8519\ : InMux
    port map (
            O => \N__42291\,
            I => \N__42288\
        );

    \I__8518\ : LocalMux
    port map (
            O => \N__42288\,
            I => \N__42285\
        );

    \I__8517\ : Span4Mux_h
    port map (
            O => \N__42285\,
            I => \N__42282\
        );

    \I__8516\ : Odrv4
    port map (
            O => \N__42282\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_24\
        );

    \I__8515\ : InMux
    port map (
            O => \N__42279\,
            I => \N__42274\
        );

    \I__8514\ : InMux
    port map (
            O => \N__42278\,
            I => \N__42269\
        );

    \I__8513\ : InMux
    port map (
            O => \N__42277\,
            I => \N__42269\
        );

    \I__8512\ : LocalMux
    port map (
            O => \N__42274\,
            I => \N__42266\
        );

    \I__8511\ : LocalMux
    port map (
            O => \N__42269\,
            I => \N__42263\
        );

    \I__8510\ : Span12Mux_h
    port map (
            O => \N__42266\,
            I => \N__42260\
        );

    \I__8509\ : Span4Mux_v
    port map (
            O => \N__42263\,
            I => \N__42257\
        );

    \I__8508\ : Odrv12
    port map (
            O => \N__42260\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_22
        );

    \I__8507\ : Odrv4
    port map (
            O => \N__42257\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_22
        );

    \I__8506\ : InMux
    port map (
            O => \N__42252\,
            I => \N__42249\
        );

    \I__8505\ : LocalMux
    port map (
            O => \N__42249\,
            I => \N__42244\
        );

    \I__8504\ : InMux
    port map (
            O => \N__42248\,
            I => \N__42239\
        );

    \I__8503\ : InMux
    port map (
            O => \N__42247\,
            I => \N__42239\
        );

    \I__8502\ : Span4Mux_h
    port map (
            O => \N__42244\,
            I => \N__42236\
        );

    \I__8501\ : LocalMux
    port map (
            O => \N__42239\,
            I => \N__42233\
        );

    \I__8500\ : Span4Mux_h
    port map (
            O => \N__42236\,
            I => \N__42230\
        );

    \I__8499\ : Span4Mux_h
    port map (
            O => \N__42233\,
            I => \N__42227\
        );

    \I__8498\ : Span4Mux_h
    port map (
            O => \N__42230\,
            I => \N__42224\
        );

    \I__8497\ : Span4Mux_h
    port map (
            O => \N__42227\,
            I => \N__42221\
        );

    \I__8496\ : Odrv4
    port map (
            O => \N__42224\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_4
        );

    \I__8495\ : Odrv4
    port map (
            O => \N__42221\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_4
        );

    \I__8494\ : InMux
    port map (
            O => \N__42216\,
            I => \N__42213\
        );

    \I__8493\ : LocalMux
    port map (
            O => \N__42213\,
            I => \N__42209\
        );

    \I__8492\ : InMux
    port map (
            O => \N__42212\,
            I => \N__42205\
        );

    \I__8491\ : Span4Mux_h
    port map (
            O => \N__42209\,
            I => \N__42202\
        );

    \I__8490\ : InMux
    port map (
            O => \N__42208\,
            I => \N__42199\
        );

    \I__8489\ : LocalMux
    port map (
            O => \N__42205\,
            I => \N__42196\
        );

    \I__8488\ : Sp12to4
    port map (
            O => \N__42202\,
            I => \N__42191\
        );

    \I__8487\ : LocalMux
    port map (
            O => \N__42199\,
            I => \N__42191\
        );

    \I__8486\ : Span4Mux_h
    port map (
            O => \N__42196\,
            I => \N__42188\
        );

    \I__8485\ : Span12Mux_v
    port map (
            O => \N__42191\,
            I => \N__42185\
        );

    \I__8484\ : Span4Mux_h
    port map (
            O => \N__42188\,
            I => \N__42182\
        );

    \I__8483\ : Odrv12
    port map (
            O => \N__42185\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_5
        );

    \I__8482\ : Odrv4
    port map (
            O => \N__42182\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_5
        );

    \I__8481\ : InMux
    port map (
            O => \N__42177\,
            I => \N__42172\
        );

    \I__8480\ : CascadeMux
    port map (
            O => \N__42176\,
            I => \N__42169\
        );

    \I__8479\ : InMux
    port map (
            O => \N__42175\,
            I => \N__42166\
        );

    \I__8478\ : LocalMux
    port map (
            O => \N__42172\,
            I => \N__42163\
        );

    \I__8477\ : InMux
    port map (
            O => \N__42169\,
            I => \N__42160\
        );

    \I__8476\ : LocalMux
    port map (
            O => \N__42166\,
            I => \N__42153\
        );

    \I__8475\ : Span4Mux_v
    port map (
            O => \N__42163\,
            I => \N__42153\
        );

    \I__8474\ : LocalMux
    port map (
            O => \N__42160\,
            I => \N__42153\
        );

    \I__8473\ : Span4Mux_h
    port map (
            O => \N__42153\,
            I => \N__42150\
        );

    \I__8472\ : Span4Mux_h
    port map (
            O => \N__42150\,
            I => \N__42147\
        );

    \I__8471\ : Odrv4
    port map (
            O => \N__42147\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_6
        );

    \I__8470\ : InMux
    port map (
            O => \N__42144\,
            I => \N__42141\
        );

    \I__8469\ : LocalMux
    port map (
            O => \N__42141\,
            I => \N__42138\
        );

    \I__8468\ : Span4Mux_v
    port map (
            O => \N__42138\,
            I => \N__42135\
        );

    \I__8467\ : Span4Mux_v
    port map (
            O => \N__42135\,
            I => \N__42132\
        );

    \I__8466\ : Sp12to4
    port map (
            O => \N__42132\,
            I => \N__42129\
        );

    \I__8465\ : Odrv12
    port map (
            O => \N__42129\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_27
        );

    \I__8464\ : CascadeMux
    port map (
            O => \N__42126\,
            I => \N__42123\
        );

    \I__8463\ : InMux
    port map (
            O => \N__42123\,
            I => \N__42120\
        );

    \I__8462\ : LocalMux
    port map (
            O => \N__42120\,
            I => \N__42117\
        );

    \I__8461\ : Span4Mux_v
    port map (
            O => \N__42117\,
            I => \N__42114\
        );

    \I__8460\ : Sp12to4
    port map (
            O => \N__42114\,
            I => \N__42111\
        );

    \I__8459\ : Span12Mux_h
    port map (
            O => \N__42111\,
            I => \N__42108\
        );

    \I__8458\ : Odrv12
    port map (
            O => \N__42108\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_27
        );

    \I__8457\ : CascadeMux
    port map (
            O => \N__42105\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_27_cascade_\
        );

    \I__8456\ : InMux
    port map (
            O => \N__42102\,
            I => \N__42099\
        );

    \I__8455\ : LocalMux
    port map (
            O => \N__42099\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_27\
        );

    \I__8454\ : InMux
    port map (
            O => \N__42096\,
            I => \N__42093\
        );

    \I__8453\ : LocalMux
    port map (
            O => \N__42093\,
            I => \N__42090\
        );

    \I__8452\ : Span4Mux_h
    port map (
            O => \N__42090\,
            I => \N__42087\
        );

    \I__8451\ : Odrv4
    port map (
            O => \N__42087\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_27\
        );

    \I__8450\ : CascadeMux
    port map (
            O => \N__42084\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_27_cascade_\
        );

    \I__8449\ : InMux
    port map (
            O => \N__42081\,
            I => \N__42078\
        );

    \I__8448\ : LocalMux
    port map (
            O => \N__42078\,
            I => \N__42075\
        );

    \I__8447\ : Odrv12
    port map (
            O => \N__42075\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_654\
        );

    \I__8446\ : InMux
    port map (
            O => \N__42072\,
            I => \N__42069\
        );

    \I__8445\ : LocalMux
    port map (
            O => \N__42069\,
            I => \N__42066\
        );

    \I__8444\ : Span12Mux_h
    port map (
            O => \N__42066\,
            I => \N__42063\
        );

    \I__8443\ : Odrv12
    port map (
            O => \N__42063\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_27\
        );

    \I__8442\ : InMux
    port map (
            O => \N__42060\,
            I => \N__42057\
        );

    \I__8441\ : LocalMux
    port map (
            O => \N__42057\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_27\
        );

    \I__8440\ : InMux
    port map (
            O => \N__42054\,
            I => \N__42051\
        );

    \I__8439\ : LocalMux
    port map (
            O => \N__42051\,
            I => \N__42048\
        );

    \I__8438\ : Span4Mux_v
    port map (
            O => \N__42048\,
            I => \N__42045\
        );

    \I__8437\ : Sp12to4
    port map (
            O => \N__42045\,
            I => \N__42042\
        );

    \I__8436\ : Span12Mux_h
    port map (
            O => \N__42042\,
            I => \N__42039\
        );

    \I__8435\ : Odrv12
    port map (
            O => \N__42039\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_16
        );

    \I__8434\ : CascadeMux
    port map (
            O => \N__42036\,
            I => \N__42033\
        );

    \I__8433\ : InMux
    port map (
            O => \N__42033\,
            I => \N__42030\
        );

    \I__8432\ : LocalMux
    port map (
            O => \N__42030\,
            I => \N__42027\
        );

    \I__8431\ : Span4Mux_v
    port map (
            O => \N__42027\,
            I => \N__42024\
        );

    \I__8430\ : Span4Mux_h
    port map (
            O => \N__42024\,
            I => \N__42021\
        );

    \I__8429\ : Sp12to4
    port map (
            O => \N__42021\,
            I => \N__42018\
        );

    \I__8428\ : Odrv12
    port map (
            O => \N__42018\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_16
        );

    \I__8427\ : CascadeMux
    port map (
            O => \N__42015\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_16_cascade_\
        );

    \I__8426\ : InMux
    port map (
            O => \N__42012\,
            I => \N__42007\
        );

    \I__8425\ : CascadeMux
    port map (
            O => \N__42011\,
            I => \N__42004\
        );

    \I__8424\ : CascadeMux
    port map (
            O => \N__42010\,
            I => \N__42001\
        );

    \I__8423\ : LocalMux
    port map (
            O => \N__42007\,
            I => \N__41998\
        );

    \I__8422\ : InMux
    port map (
            O => \N__42004\,
            I => \N__41993\
        );

    \I__8421\ : InMux
    port map (
            O => \N__42001\,
            I => \N__41993\
        );

    \I__8420\ : Odrv4
    port map (
            O => \N__41998\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_16
        );

    \I__8419\ : LocalMux
    port map (
            O => \N__41993\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_16
        );

    \I__8418\ : InMux
    port map (
            O => \N__41988\,
            I => \N__41985\
        );

    \I__8417\ : LocalMux
    port map (
            O => \N__41985\,
            I => \N__41982\
        );

    \I__8416\ : Span12Mux_s10_v
    port map (
            O => \N__41982\,
            I => \N__41979\
        );

    \I__8415\ : Span12Mux_v
    port map (
            O => \N__41979\,
            I => \N__41976\
        );

    \I__8414\ : Span12Mux_h
    port map (
            O => \N__41976\,
            I => \N__41973\
        );

    \I__8413\ : Odrv12
    port map (
            O => \N__41973\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_16
        );

    \I__8412\ : InMux
    port map (
            O => \N__41970\,
            I => \N__41967\
        );

    \I__8411\ : LocalMux
    port map (
            O => \N__41967\,
            I => \N__41964\
        );

    \I__8410\ : Span4Mux_h
    port map (
            O => \N__41964\,
            I => \N__41961\
        );

    \I__8409\ : Span4Mux_v
    port map (
            O => \N__41961\,
            I => \N__41958\
        );

    \I__8408\ : Span4Mux_h
    port map (
            O => \N__41958\,
            I => \N__41955\
        );

    \I__8407\ : Odrv4
    port map (
            O => \N__41955\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_764\
        );

    \I__8406\ : CascadeMux
    port map (
            O => \N__41952\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_16_cascade_\
        );

    \I__8405\ : InMux
    port map (
            O => \N__41949\,
            I => \N__41946\
        );

    \I__8404\ : LocalMux
    port map (
            O => \N__41946\,
            I => \serializer_mod_inst.shift_regZ0Z_27\
        );

    \I__8403\ : InMux
    port map (
            O => \N__41943\,
            I => \N__41940\
        );

    \I__8402\ : LocalMux
    port map (
            O => \N__41940\,
            I => \serializer_mod_inst.shift_regZ0Z_22\
        );

    \I__8401\ : InMux
    port map (
            O => \N__41937\,
            I => \N__41934\
        );

    \I__8400\ : LocalMux
    port map (
            O => \N__41934\,
            I => \serializer_mod_inst.shift_regZ0Z_23\
        );

    \I__8399\ : InMux
    port map (
            O => \N__41931\,
            I => \N__41928\
        );

    \I__8398\ : LocalMux
    port map (
            O => \N__41928\,
            I => \N__41925\
        );

    \I__8397\ : Odrv4
    port map (
            O => \N__41925\,
            I => \serializer_mod_inst.shift_regZ0Z_108\
        );

    \I__8396\ : InMux
    port map (
            O => \N__41922\,
            I => \N__41919\
        );

    \I__8395\ : LocalMux
    port map (
            O => \N__41919\,
            I => \N__41916\
        );

    \I__8394\ : Odrv12
    port map (
            O => \N__41916\,
            I => \serializer_mod_inst.shift_regZ0Z_109\
        );

    \I__8393\ : InMux
    port map (
            O => \N__41913\,
            I => \N__41910\
        );

    \I__8392\ : LocalMux
    port map (
            O => \N__41910\,
            I => \N__41907\
        );

    \I__8391\ : Odrv4
    port map (
            O => \N__41907\,
            I => \serializer_mod_inst.shift_regZ0Z_19\
        );

    \I__8390\ : InMux
    port map (
            O => \N__41904\,
            I => \N__41901\
        );

    \I__8389\ : LocalMux
    port map (
            O => \N__41901\,
            I => \serializer_mod_inst.shift_regZ0Z_20\
        );

    \I__8388\ : InMux
    port map (
            O => \N__41898\,
            I => \N__41895\
        );

    \I__8387\ : LocalMux
    port map (
            O => \N__41895\,
            I => \serializer_mod_inst.shift_regZ0Z_24\
        );

    \I__8386\ : InMux
    port map (
            O => \N__41892\,
            I => \N__41889\
        );

    \I__8385\ : LocalMux
    port map (
            O => \N__41889\,
            I => \serializer_mod_inst.shift_regZ0Z_124\
        );

    \I__8384\ : InMux
    port map (
            O => \N__41886\,
            I => \N__41883\
        );

    \I__8383\ : LocalMux
    port map (
            O => \N__41883\,
            I => \N__41880\
        );

    \I__8382\ : Odrv4
    port map (
            O => \N__41880\,
            I => \serializer_mod_inst.shift_regZ0Z_125\
        );

    \I__8381\ : InMux
    port map (
            O => \N__41877\,
            I => \N__41874\
        );

    \I__8380\ : LocalMux
    port map (
            O => \N__41874\,
            I => \N__41871\
        );

    \I__8379\ : Span4Mux_v
    port map (
            O => \N__41871\,
            I => \N__41868\
        );

    \I__8378\ : Odrv4
    port map (
            O => \N__41868\,
            I => \serializer_mod_inst.shift_regZ0Z_122\
        );

    \I__8377\ : InMux
    port map (
            O => \N__41865\,
            I => \N__41862\
        );

    \I__8376\ : LocalMux
    port map (
            O => \N__41862\,
            I => \serializer_mod_inst.shift_regZ0Z_123\
        );

    \I__8375\ : InMux
    port map (
            O => \N__41859\,
            I => \N__41856\
        );

    \I__8374\ : LocalMux
    port map (
            O => \N__41856\,
            I => \serializer_mod_inst.shift_regZ0Z_25\
        );

    \I__8373\ : InMux
    port map (
            O => \N__41853\,
            I => \N__41850\
        );

    \I__8372\ : LocalMux
    port map (
            O => \N__41850\,
            I => \serializer_mod_inst.shift_regZ0Z_26\
        );

    \I__8371\ : InMux
    port map (
            O => \N__41847\,
            I => \N__41844\
        );

    \I__8370\ : LocalMux
    port map (
            O => \N__41844\,
            I => \N__41841\
        );

    \I__8369\ : Odrv12
    port map (
            O => \N__41841\,
            I => \serializer_mod_inst.shift_regZ0Z_6\
        );

    \I__8368\ : InMux
    port map (
            O => \N__41838\,
            I => \N__41835\
        );

    \I__8367\ : LocalMux
    port map (
            O => \N__41835\,
            I => \serializer_mod_inst.shift_regZ0Z_5\
        );

    \I__8366\ : InMux
    port map (
            O => \N__41832\,
            I => \N__41829\
        );

    \I__8365\ : LocalMux
    port map (
            O => \N__41829\,
            I => \serializer_mod_inst.shift_regZ0Z_2\
        );

    \I__8364\ : InMux
    port map (
            O => \N__41826\,
            I => \N__41823\
        );

    \I__8363\ : LocalMux
    port map (
            O => \N__41823\,
            I => \serializer_mod_inst.shift_regZ0Z_3\
        );

    \I__8362\ : InMux
    port map (
            O => \N__41820\,
            I => \N__41817\
        );

    \I__8361\ : LocalMux
    port map (
            O => \N__41817\,
            I => \serializer_mod_inst.shift_regZ0Z_4\
        );

    \I__8360\ : InMux
    port map (
            O => \N__41814\,
            I => \N__41811\
        );

    \I__8359\ : LocalMux
    port map (
            O => \N__41811\,
            I => \serializer_mod_inst.shift_regZ0Z_21\
        );

    \I__8358\ : InMux
    port map (
            O => \N__41808\,
            I => \N__41803\
        );

    \I__8357\ : InMux
    port map (
            O => \N__41807\,
            I => \N__41800\
        );

    \I__8356\ : InMux
    port map (
            O => \N__41806\,
            I => \N__41797\
        );

    \I__8355\ : LocalMux
    port map (
            O => \N__41803\,
            I => \N__41791\
        );

    \I__8354\ : LocalMux
    port map (
            O => \N__41800\,
            I => \N__41791\
        );

    \I__8353\ : LocalMux
    port map (
            O => \N__41797\,
            I => \N__41788\
        );

    \I__8352\ : InMux
    port map (
            O => \N__41796\,
            I => \N__41783\
        );

    \I__8351\ : Span12Mux_v
    port map (
            O => \N__41791\,
            I => \N__41778\
        );

    \I__8350\ : Span12Mux_v
    port map (
            O => \N__41788\,
            I => \N__41778\
        );

    \I__8349\ : InMux
    port map (
            O => \N__41787\,
            I => \N__41773\
        );

    \I__8348\ : InMux
    port map (
            O => \N__41786\,
            I => \N__41773\
        );

    \I__8347\ : LocalMux
    port map (
            O => \N__41783\,
            I => \I2C_top_level_inst1.s_data_ireg_5\
        );

    \I__8346\ : Odrv12
    port map (
            O => \N__41778\,
            I => \I2C_top_level_inst1.s_data_ireg_5\
        );

    \I__8345\ : LocalMux
    port map (
            O => \N__41773\,
            I => \I2C_top_level_inst1.s_data_ireg_5\
        );

    \I__8344\ : CascadeMux
    port map (
            O => \N__41766\,
            I => \N__41763\
        );

    \I__8343\ : InMux
    port map (
            O => \N__41763\,
            I => \N__41760\
        );

    \I__8342\ : LocalMux
    port map (
            O => \N__41760\,
            I => \I2C_top_level_inst1.s_addr0_o_5\
        );

    \I__8341\ : InMux
    port map (
            O => \N__41757\,
            I => \N__41754\
        );

    \I__8340\ : LocalMux
    port map (
            O => \N__41754\,
            I => \N__41749\
        );

    \I__8339\ : InMux
    port map (
            O => \N__41753\,
            I => \N__41746\
        );

    \I__8338\ : InMux
    port map (
            O => \N__41752\,
            I => \N__41743\
        );

    \I__8337\ : Span4Mux_v
    port map (
            O => \N__41749\,
            I => \N__41740\
        );

    \I__8336\ : LocalMux
    port map (
            O => \N__41746\,
            I => \N__41735\
        );

    \I__8335\ : LocalMux
    port map (
            O => \N__41743\,
            I => \N__41735\
        );

    \I__8334\ : Span4Mux_h
    port map (
            O => \N__41740\,
            I => \N__41730\
        );

    \I__8333\ : Span4Mux_v
    port map (
            O => \N__41735\,
            I => \N__41726\
        );

    \I__8332\ : InMux
    port map (
            O => \N__41734\,
            I => \N__41723\
        );

    \I__8331\ : InMux
    port map (
            O => \N__41733\,
            I => \N__41720\
        );

    \I__8330\ : Span4Mux_h
    port map (
            O => \N__41730\,
            I => \N__41717\
        );

    \I__8329\ : InMux
    port map (
            O => \N__41729\,
            I => \N__41714\
        );

    \I__8328\ : Odrv4
    port map (
            O => \N__41726\,
            I => \I2C_top_level_inst1.s_data_ireg_6\
        );

    \I__8327\ : LocalMux
    port map (
            O => \N__41723\,
            I => \I2C_top_level_inst1.s_data_ireg_6\
        );

    \I__8326\ : LocalMux
    port map (
            O => \N__41720\,
            I => \I2C_top_level_inst1.s_data_ireg_6\
        );

    \I__8325\ : Odrv4
    port map (
            O => \N__41717\,
            I => \I2C_top_level_inst1.s_data_ireg_6\
        );

    \I__8324\ : LocalMux
    port map (
            O => \N__41714\,
            I => \I2C_top_level_inst1.s_data_ireg_6\
        );

    \I__8323\ : CascadeMux
    port map (
            O => \N__41703\,
            I => \N__41700\
        );

    \I__8322\ : InMux
    port map (
            O => \N__41700\,
            I => \N__41697\
        );

    \I__8321\ : LocalMux
    port map (
            O => \N__41697\,
            I => \N__41694\
        );

    \I__8320\ : Odrv4
    port map (
            O => \N__41694\,
            I => \I2C_top_level_inst1.s_addr0_o_6\
        );

    \I__8319\ : InMux
    port map (
            O => \N__41691\,
            I => \N__41685\
        );

    \I__8318\ : InMux
    port map (
            O => \N__41690\,
            I => \N__41682\
        );

    \I__8317\ : InMux
    port map (
            O => \N__41689\,
            I => \N__41679\
        );

    \I__8316\ : InMux
    port map (
            O => \N__41688\,
            I => \N__41676\
        );

    \I__8315\ : LocalMux
    port map (
            O => \N__41685\,
            I => \N__41671\
        );

    \I__8314\ : LocalMux
    port map (
            O => \N__41682\,
            I => \N__41671\
        );

    \I__8313\ : LocalMux
    port map (
            O => \N__41679\,
            I => \N__41668\
        );

    \I__8312\ : LocalMux
    port map (
            O => \N__41676\,
            I => \N__41665\
        );

    \I__8311\ : Span4Mux_v
    port map (
            O => \N__41671\,
            I => \N__41662\
        );

    \I__8310\ : Span4Mux_v
    port map (
            O => \N__41668\,
            I => \N__41659\
        );

    \I__8309\ : Span4Mux_h
    port map (
            O => \N__41665\,
            I => \N__41655\
        );

    \I__8308\ : Span4Mux_h
    port map (
            O => \N__41662\,
            I => \N__41652\
        );

    \I__8307\ : Sp12to4
    port map (
            O => \N__41659\,
            I => \N__41649\
        );

    \I__8306\ : CascadeMux
    port map (
            O => \N__41658\,
            I => \N__41646\
        );

    \I__8305\ : Span4Mux_h
    port map (
            O => \N__41655\,
            I => \N__41643\
        );

    \I__8304\ : Sp12to4
    port map (
            O => \N__41652\,
            I => \N__41638\
        );

    \I__8303\ : Span12Mux_h
    port map (
            O => \N__41649\,
            I => \N__41638\
        );

    \I__8302\ : InMux
    port map (
            O => \N__41646\,
            I => \N__41635\
        );

    \I__8301\ : Odrv4
    port map (
            O => \N__41643\,
            I => \I2C_top_level_inst1.s_data_ireg_7\
        );

    \I__8300\ : Odrv12
    port map (
            O => \N__41638\,
            I => \I2C_top_level_inst1.s_data_ireg_7\
        );

    \I__8299\ : LocalMux
    port map (
            O => \N__41635\,
            I => \I2C_top_level_inst1.s_data_ireg_7\
        );

    \I__8298\ : CascadeMux
    port map (
            O => \N__41628\,
            I => \N__41625\
        );

    \I__8297\ : InMux
    port map (
            O => \N__41625\,
            I => \N__41622\
        );

    \I__8296\ : LocalMux
    port map (
            O => \N__41622\,
            I => \I2C_top_level_inst1.s_addr0_o_7\
        );

    \I__8295\ : InMux
    port map (
            O => \N__41619\,
            I => \N__41616\
        );

    \I__8294\ : LocalMux
    port map (
            O => \N__41616\,
            I => \N__41613\
        );

    \I__8293\ : Span4Mux_h
    port map (
            O => \N__41613\,
            I => \N__41610\
        );

    \I__8292\ : Span4Mux_v
    port map (
            O => \N__41610\,
            I => \N__41606\
        );

    \I__8291\ : InMux
    port map (
            O => \N__41609\,
            I => \N__41603\
        );

    \I__8290\ : Odrv4
    port map (
            O => \N__41606\,
            I => \N_396\
        );

    \I__8289\ : LocalMux
    port map (
            O => \N__41603\,
            I => \N_396\
        );

    \I__8288\ : CascadeMux
    port map (
            O => \N__41598\,
            I => \N__41595\
        );

    \I__8287\ : InMux
    port map (
            O => \N__41595\,
            I => \N__41592\
        );

    \I__8286\ : LocalMux
    port map (
            O => \N__41592\,
            I => \N__41589\
        );

    \I__8285\ : Span12Mux_h
    port map (
            O => \N__41589\,
            I => \N__41586\
        );

    \I__8284\ : Odrv12
    port map (
            O => \N__41586\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_3\
        );

    \I__8283\ : CascadeMux
    port map (
            O => \N__41583\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_4_cascade_\
        );

    \I__8282\ : CascadeMux
    port map (
            O => \N__41580\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNOZ0Z_0_cascade_\
        );

    \I__8281\ : InMux
    port map (
            O => \N__41577\,
            I => \N__41571\
        );

    \I__8280\ : InMux
    port map (
            O => \N__41576\,
            I => \N__41564\
        );

    \I__8279\ : InMux
    port map (
            O => \N__41575\,
            I => \N__41564\
        );

    \I__8278\ : InMux
    port map (
            O => \N__41574\,
            I => \N__41564\
        );

    \I__8277\ : LocalMux
    port map (
            O => \N__41571\,
            I => \N__41560\
        );

    \I__8276\ : LocalMux
    port map (
            O => \N__41564\,
            I => \N__41557\
        );

    \I__8275\ : InMux
    port map (
            O => \N__41563\,
            I => \N__41554\
        );

    \I__8274\ : Span4Mux_h
    port map (
            O => \N__41560\,
            I => \N__41551\
        );

    \I__8273\ : Span4Mux_h
    port map (
            O => \N__41557\,
            I => \N__41548\
        );

    \I__8272\ : LocalMux
    port map (
            O => \N__41554\,
            I => \I2C_top_level_inst1.s_no_restart\
        );

    \I__8271\ : Odrv4
    port map (
            O => \N__41551\,
            I => \I2C_top_level_inst1.s_no_restart\
        );

    \I__8270\ : Odrv4
    port map (
            O => \N__41548\,
            I => \I2C_top_level_inst1.s_no_restart\
        );

    \I__8269\ : InMux
    port map (
            O => \N__41541\,
            I => \N__41538\
        );

    \I__8268\ : LocalMux
    port map (
            O => \N__41538\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_1\
        );

    \I__8267\ : InMux
    port map (
            O => \N__41535\,
            I => \N__41532\
        );

    \I__8266\ : LocalMux
    port map (
            O => \N__41532\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_304_0\
        );

    \I__8265\ : CascadeMux
    port map (
            O => \N__41529\,
            I => \N__41526\
        );

    \I__8264\ : InMux
    port map (
            O => \N__41526\,
            I => \N__41523\
        );

    \I__8263\ : LocalMux
    port map (
            O => \N__41523\,
            I => \N__41518\
        );

    \I__8262\ : InMux
    port map (
            O => \N__41522\,
            I => \N__41512\
        );

    \I__8261\ : InMux
    port map (
            O => \N__41521\,
            I => \N__41512\
        );

    \I__8260\ : Span4Mux_v
    port map (
            O => \N__41518\,
            I => \N__41509\
        );

    \I__8259\ : CascadeMux
    port map (
            O => \N__41517\,
            I => \N__41506\
        );

    \I__8258\ : LocalMux
    port map (
            O => \N__41512\,
            I => \N__41503\
        );

    \I__8257\ : Span4Mux_h
    port map (
            O => \N__41509\,
            I => \N__41500\
        );

    \I__8256\ : InMux
    port map (
            O => \N__41506\,
            I => \N__41497\
        );

    \I__8255\ : Span4Mux_h
    port map (
            O => \N__41503\,
            I => \N__41494\
        );

    \I__8254\ : Odrv4
    port map (
            O => \N__41500\,
            I => \I2C_top_level_inst1.s_ack\
        );

    \I__8253\ : LocalMux
    port map (
            O => \N__41497\,
            I => \I2C_top_level_inst1.s_ack\
        );

    \I__8252\ : Odrv4
    port map (
            O => \N__41494\,
            I => \I2C_top_level_inst1.s_ack\
        );

    \I__8251\ : CascadeMux
    port map (
            O => \N__41487\,
            I => \N__41484\
        );

    \I__8250\ : InMux
    port map (
            O => \N__41484\,
            I => \N__41481\
        );

    \I__8249\ : LocalMux
    port map (
            O => \N__41481\,
            I => \N__41478\
        );

    \I__8248\ : Span4Mux_v
    port map (
            O => \N__41478\,
            I => \N__41475\
        );

    \I__8247\ : Span4Mux_h
    port map (
            O => \N__41475\,
            I => \N__41472\
        );

    \I__8246\ : Odrv4
    port map (
            O => \N__41472\,
            I => \I2C_top_level_inst1.s_addr1_o_4\
        );

    \I__8245\ : CascadeMux
    port map (
            O => \N__41469\,
            I => \N__41466\
        );

    \I__8244\ : InMux
    port map (
            O => \N__41466\,
            I => \N__41463\
        );

    \I__8243\ : LocalMux
    port map (
            O => \N__41463\,
            I => \N__41460\
        );

    \I__8242\ : Span4Mux_h
    port map (
            O => \N__41460\,
            I => \N__41457\
        );

    \I__8241\ : Odrv4
    port map (
            O => \N__41457\,
            I => \I2C_top_level_inst1.s_addr1_o_5\
        );

    \I__8240\ : CascadeMux
    port map (
            O => \N__41454\,
            I => \N__41451\
        );

    \I__8239\ : InMux
    port map (
            O => \N__41451\,
            I => \N__41448\
        );

    \I__8238\ : LocalMux
    port map (
            O => \N__41448\,
            I => \N__41445\
        );

    \I__8237\ : Span4Mux_h
    port map (
            O => \N__41445\,
            I => \N__41442\
        );

    \I__8236\ : Odrv4
    port map (
            O => \N__41442\,
            I => \I2C_top_level_inst1.s_addr1_o_6\
        );

    \I__8235\ : CascadeMux
    port map (
            O => \N__41439\,
            I => \N__41436\
        );

    \I__8234\ : InMux
    port map (
            O => \N__41436\,
            I => \N__41433\
        );

    \I__8233\ : LocalMux
    port map (
            O => \N__41433\,
            I => \N__41430\
        );

    \I__8232\ : Span4Mux_v
    port map (
            O => \N__41430\,
            I => \N__41427\
        );

    \I__8231\ : Odrv4
    port map (
            O => \N__41427\,
            I => \I2C_top_level_inst1.s_addr1_o_7\
        );

    \I__8230\ : InMux
    port map (
            O => \N__41424\,
            I => \N__41421\
        );

    \I__8229\ : LocalMux
    port map (
            O => \N__41421\,
            I => \N__41417\
        );

    \I__8228\ : CEMux
    port map (
            O => \N__41420\,
            I => \N__41414\
        );

    \I__8227\ : Span4Mux_h
    port map (
            O => \N__41417\,
            I => \N__41410\
        );

    \I__8226\ : LocalMux
    port map (
            O => \N__41414\,
            I => \N__41407\
        );

    \I__8225\ : InMux
    port map (
            O => \N__41413\,
            I => \N__41403\
        );

    \I__8224\ : Sp12to4
    port map (
            O => \N__41410\,
            I => \N__41400\
        );

    \I__8223\ : Span4Mux_h
    port map (
            O => \N__41407\,
            I => \N__41397\
        );

    \I__8222\ : InMux
    port map (
            O => \N__41406\,
            I => \N__41394\
        );

    \I__8221\ : LocalMux
    port map (
            O => \N__41403\,
            I => \I2C_top_level_inst1.s_load_addr1\
        );

    \I__8220\ : Odrv12
    port map (
            O => \N__41400\,
            I => \I2C_top_level_inst1.s_load_addr1\
        );

    \I__8219\ : Odrv4
    port map (
            O => \N__41397\,
            I => \I2C_top_level_inst1.s_load_addr1\
        );

    \I__8218\ : LocalMux
    port map (
            O => \N__41394\,
            I => \I2C_top_level_inst1.s_load_addr1\
        );

    \I__8217\ : InMux
    port map (
            O => \N__41385\,
            I => \N__41382\
        );

    \I__8216\ : LocalMux
    port map (
            O => \N__41382\,
            I => \I2C_top_level_inst1.s_addr0_o_3\
        );

    \I__8215\ : InMux
    port map (
            O => \N__41379\,
            I => \N__41372\
        );

    \I__8214\ : InMux
    port map (
            O => \N__41378\,
            I => \N__41369\
        );

    \I__8213\ : InMux
    port map (
            O => \N__41377\,
            I => \N__41366\
        );

    \I__8212\ : InMux
    port map (
            O => \N__41376\,
            I => \N__41363\
        );

    \I__8211\ : InMux
    port map (
            O => \N__41375\,
            I => \N__41360\
        );

    \I__8210\ : LocalMux
    port map (
            O => \N__41372\,
            I => \N__41355\
        );

    \I__8209\ : LocalMux
    port map (
            O => \N__41369\,
            I => \N__41355\
        );

    \I__8208\ : LocalMux
    port map (
            O => \N__41366\,
            I => \N__41352\
        );

    \I__8207\ : LocalMux
    port map (
            O => \N__41363\,
            I => \N__41349\
        );

    \I__8206\ : LocalMux
    port map (
            O => \N__41360\,
            I => \N__41343\
        );

    \I__8205\ : Span4Mux_v
    port map (
            O => \N__41355\,
            I => \N__41343\
        );

    \I__8204\ : Span4Mux_h
    port map (
            O => \N__41352\,
            I => \N__41338\
        );

    \I__8203\ : Span4Mux_v
    port map (
            O => \N__41349\,
            I => \N__41338\
        );

    \I__8202\ : InMux
    port map (
            O => \N__41348\,
            I => \N__41335\
        );

    \I__8201\ : Odrv4
    port map (
            O => \N__41343\,
            I => \I2C_top_level_inst1.s_data_ireg_4\
        );

    \I__8200\ : Odrv4
    port map (
            O => \N__41338\,
            I => \I2C_top_level_inst1.s_data_ireg_4\
        );

    \I__8199\ : LocalMux
    port map (
            O => \N__41335\,
            I => \I2C_top_level_inst1.s_data_ireg_4\
        );

    \I__8198\ : CascadeMux
    port map (
            O => \N__41328\,
            I => \N__41325\
        );

    \I__8197\ : InMux
    port map (
            O => \N__41325\,
            I => \N__41322\
        );

    \I__8196\ : LocalMux
    port map (
            O => \N__41322\,
            I => \N__41319\
        );

    \I__8195\ : Odrv4
    port map (
            O => \N__41319\,
            I => \I2C_top_level_inst1.s_addr0_o_4\
        );

    \I__8194\ : CascadeMux
    port map (
            O => \N__41316\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0_cascade_\
        );

    \I__8193\ : CascadeMux
    port map (
            O => \N__41313\,
            I => \N__41310\
        );

    \I__8192\ : InMux
    port map (
            O => \N__41310\,
            I => \N__41307\
        );

    \I__8191\ : LocalMux
    port map (
            O => \N__41307\,
            I => \I2C_top_level_inst1.s_addr1_o_1\
        );

    \I__8190\ : InMux
    port map (
            O => \N__41304\,
            I => \N__41301\
        );

    \I__8189\ : LocalMux
    port map (
            O => \N__41301\,
            I => \I2C_top_level_inst1.s_addr1_o_2\
        );

    \I__8188\ : InMux
    port map (
            O => \N__41298\,
            I => \N__41295\
        );

    \I__8187\ : LocalMux
    port map (
            O => \N__41295\,
            I => \I2C_top_level_inst1.s_addr1_o_3\
        );

    \I__8186\ : InMux
    port map (
            O => \N__41292\,
            I => \N__41289\
        );

    \I__8185\ : LocalMux
    port map (
            O => \N__41289\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11\
        );

    \I__8184\ : CascadeMux
    port map (
            O => \N__41286\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11_cascade_\
        );

    \I__8183\ : InMux
    port map (
            O => \N__41283\,
            I => \N__41280\
        );

    \I__8182\ : LocalMux
    port map (
            O => \N__41280\,
            I => \N__41277\
        );

    \I__8181\ : Odrv12
    port map (
            O => \N__41277\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_12\
        );

    \I__8180\ : CascadeMux
    port map (
            O => \N__41274\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GHZ0Z5_cascade_\
        );

    \I__8179\ : InMux
    port map (
            O => \N__41271\,
            I => \N__41268\
        );

    \I__8178\ : LocalMux
    port map (
            O => \N__41268\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12\
        );

    \I__8177\ : InMux
    port map (
            O => \N__41265\,
            I => \N__41262\
        );

    \I__8176\ : LocalMux
    port map (
            O => \N__41262\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_11\
        );

    \I__8175\ : CascadeMux
    port map (
            O => \N__41259\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12_cascade_\
        );

    \I__8174\ : InMux
    port map (
            O => \N__41256\,
            I => \N__41253\
        );

    \I__8173\ : LocalMux
    port map (
            O => \N__41253\,
            I => \N__41250\
        );

    \I__8172\ : Span4Mux_v
    port map (
            O => \N__41250\,
            I => \N__41247\
        );

    \I__8171\ : Span4Mux_h
    port map (
            O => \N__41247\,
            I => \N__41244\
        );

    \I__8170\ : Span4Mux_h
    port map (
            O => \N__41244\,
            I => \N__41241\
        );

    \I__8169\ : Odrv4
    port map (
            O => \N__41241\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_12\
        );

    \I__8168\ : CascadeMux
    port map (
            O => \N__41238\,
            I => \N__41235\
        );

    \I__8167\ : InMux
    port map (
            O => \N__41235\,
            I => \N__41231\
        );

    \I__8166\ : InMux
    port map (
            O => \N__41234\,
            I => \N__41228\
        );

    \I__8165\ : LocalMux
    port map (
            O => \N__41231\,
            I => \N__41225\
        );

    \I__8164\ : LocalMux
    port map (
            O => \N__41228\,
            I => \N__41222\
        );

    \I__8163\ : Span4Mux_v
    port map (
            O => \N__41225\,
            I => \N__41218\
        );

    \I__8162\ : Span4Mux_v
    port map (
            O => \N__41222\,
            I => \N__41215\
        );

    \I__8161\ : InMux
    port map (
            O => \N__41221\,
            I => \N__41212\
        );

    \I__8160\ : Span4Mux_h
    port map (
            O => \N__41218\,
            I => \N__41209\
        );

    \I__8159\ : Odrv4
    port map (
            O => \N__41215\,
            I => cemf_module_64ch_ctrl_inst1_data_config_12
        );

    \I__8158\ : LocalMux
    port map (
            O => \N__41212\,
            I => cemf_module_64ch_ctrl_inst1_data_config_12
        );

    \I__8157\ : Odrv4
    port map (
            O => \N__41209\,
            I => cemf_module_64ch_ctrl_inst1_data_config_12
        );

    \I__8156\ : InMux
    port map (
            O => \N__41202\,
            I => \N__41198\
        );

    \I__8155\ : InMux
    port map (
            O => \N__41201\,
            I => \N__41194\
        );

    \I__8154\ : LocalMux
    port map (
            O => \N__41198\,
            I => \N__41191\
        );

    \I__8153\ : CascadeMux
    port map (
            O => \N__41197\,
            I => \N__41188\
        );

    \I__8152\ : LocalMux
    port map (
            O => \N__41194\,
            I => \N__41185\
        );

    \I__8151\ : Span4Mux_h
    port map (
            O => \N__41191\,
            I => \N__41182\
        );

    \I__8150\ : InMux
    port map (
            O => \N__41188\,
            I => \N__41179\
        );

    \I__8149\ : Span4Mux_v
    port map (
            O => \N__41185\,
            I => \N__41176\
        );

    \I__8148\ : Odrv4
    port map (
            O => \N__41182\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_12
        );

    \I__8147\ : LocalMux
    port map (
            O => \N__41179\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_12
        );

    \I__8146\ : Odrv4
    port map (
            O => \N__41176\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_12
        );

    \I__8145\ : CascadeMux
    port map (
            O => \N__41169\,
            I => \N__41166\
        );

    \I__8144\ : InMux
    port map (
            O => \N__41166\,
            I => \N__41163\
        );

    \I__8143\ : LocalMux
    port map (
            O => \N__41163\,
            I => \N__41160\
        );

    \I__8142\ : Odrv4
    port map (
            O => \N__41160\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_12\
        );

    \I__8141\ : CascadeMux
    port map (
            O => \N__41157\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_11_cascade_\
        );

    \I__8140\ : InMux
    port map (
            O => \N__41154\,
            I => \N__41151\
        );

    \I__8139\ : LocalMux
    port map (
            O => \N__41151\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFHZ0Z5\
        );

    \I__8138\ : CascadeMux
    port map (
            O => \N__41148\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13_cascade_\
        );

    \I__8137\ : InMux
    port map (
            O => \N__41145\,
            I => \N__41142\
        );

    \I__8136\ : LocalMux
    port map (
            O => \N__41142\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_12\
        );

    \I__8135\ : InMux
    port map (
            O => \N__41139\,
            I => \N__41136\
        );

    \I__8134\ : LocalMux
    port map (
            O => \N__41136\,
            I => \N__41133\
        );

    \I__8133\ : Span4Mux_h
    port map (
            O => \N__41133\,
            I => \N__41130\
        );

    \I__8132\ : Odrv4
    port map (
            O => \N__41130\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_13\
        );

    \I__8131\ : InMux
    port map (
            O => \N__41127\,
            I => \N__41122\
        );

    \I__8130\ : CascadeMux
    port map (
            O => \N__41126\,
            I => \N__41119\
        );

    \I__8129\ : CascadeMux
    port map (
            O => \N__41125\,
            I => \N__41116\
        );

    \I__8128\ : LocalMux
    port map (
            O => \N__41122\,
            I => \N__41113\
        );

    \I__8127\ : InMux
    port map (
            O => \N__41119\,
            I => \N__41110\
        );

    \I__8126\ : InMux
    port map (
            O => \N__41116\,
            I => \N__41107\
        );

    \I__8125\ : Span4Mux_v
    port map (
            O => \N__41113\,
            I => \N__41104\
        );

    \I__8124\ : LocalMux
    port map (
            O => \N__41110\,
            I => \N__41101\
        );

    \I__8123\ : LocalMux
    port map (
            O => \N__41107\,
            I => \N__41098\
        );

    \I__8122\ : Span4Mux_h
    port map (
            O => \N__41104\,
            I => \N__41093\
        );

    \I__8121\ : Span4Mux_v
    port map (
            O => \N__41101\,
            I => \N__41093\
        );

    \I__8120\ : Odrv12
    port map (
            O => \N__41098\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_5
        );

    \I__8119\ : Odrv4
    port map (
            O => \N__41093\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_5
        );

    \I__8118\ : CascadeMux
    port map (
            O => \N__41088\,
            I => \N__41084\
        );

    \I__8117\ : InMux
    port map (
            O => \N__41087\,
            I => \N__41078\
        );

    \I__8116\ : InMux
    port map (
            O => \N__41084\,
            I => \N__41078\
        );

    \I__8115\ : InMux
    port map (
            O => \N__41083\,
            I => \N__41075\
        );

    \I__8114\ : LocalMux
    port map (
            O => \N__41078\,
            I => \N__41072\
        );

    \I__8113\ : LocalMux
    port map (
            O => \N__41075\,
            I => \N__41067\
        );

    \I__8112\ : Span4Mux_v
    port map (
            O => \N__41072\,
            I => \N__41067\
        );

    \I__8111\ : Span4Mux_v
    port map (
            O => \N__41067\,
            I => \N__41064\
        );

    \I__8110\ : Span4Mux_h
    port map (
            O => \N__41064\,
            I => \N__41061\
        );

    \I__8109\ : Odrv4
    port map (
            O => \N__41061\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_6
        );

    \I__8108\ : InMux
    port map (
            O => \N__41058\,
            I => \N__41055\
        );

    \I__8107\ : LocalMux
    port map (
            O => \N__41055\,
            I => \N__41050\
        );

    \I__8106\ : CascadeMux
    port map (
            O => \N__41054\,
            I => \N__41047\
        );

    \I__8105\ : CascadeMux
    port map (
            O => \N__41053\,
            I => \N__41044\
        );

    \I__8104\ : Span12Mux_v
    port map (
            O => \N__41050\,
            I => \N__41041\
        );

    \I__8103\ : InMux
    port map (
            O => \N__41047\,
            I => \N__41038\
        );

    \I__8102\ : InMux
    port map (
            O => \N__41044\,
            I => \N__41035\
        );

    \I__8101\ : Span12Mux_h
    port map (
            O => \N__41041\,
            I => \N__41028\
        );

    \I__8100\ : LocalMux
    port map (
            O => \N__41038\,
            I => \N__41028\
        );

    \I__8099\ : LocalMux
    port map (
            O => \N__41035\,
            I => \N__41028\
        );

    \I__8098\ : Odrv12
    port map (
            O => \N__41028\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_7
        );

    \I__8097\ : InMux
    port map (
            O => \N__41025\,
            I => \N__41022\
        );

    \I__8096\ : LocalMux
    port map (
            O => \N__41022\,
            I => \N__41017\
        );

    \I__8095\ : CascadeMux
    port map (
            O => \N__41021\,
            I => \N__41014\
        );

    \I__8094\ : CascadeMux
    port map (
            O => \N__41020\,
            I => \N__41011\
        );

    \I__8093\ : Span4Mux_h
    port map (
            O => \N__41017\,
            I => \N__41008\
        );

    \I__8092\ : InMux
    port map (
            O => \N__41014\,
            I => \N__41005\
        );

    \I__8091\ : InMux
    port map (
            O => \N__41011\,
            I => \N__41002\
        );

    \I__8090\ : Span4Mux_h
    port map (
            O => \N__41008\,
            I => \N__40997\
        );

    \I__8089\ : LocalMux
    port map (
            O => \N__41005\,
            I => \N__40997\
        );

    \I__8088\ : LocalMux
    port map (
            O => \N__41002\,
            I => \N__40994\
        );

    \I__8087\ : Span4Mux_v
    port map (
            O => \N__40997\,
            I => \N__40991\
        );

    \I__8086\ : Odrv4
    port map (
            O => \N__40994\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_8
        );

    \I__8085\ : Odrv4
    port map (
            O => \N__40991\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_8
        );

    \I__8084\ : InMux
    port map (
            O => \N__40986\,
            I => \N__40982\
        );

    \I__8083\ : InMux
    port map (
            O => \N__40985\,
            I => \N__40979\
        );

    \I__8082\ : LocalMux
    port map (
            O => \N__40982\,
            I => \N__40974\
        );

    \I__8081\ : LocalMux
    port map (
            O => \N__40979\,
            I => \N__40974\
        );

    \I__8080\ : Span4Mux_h
    port map (
            O => \N__40974\,
            I => \N__40970\
        );

    \I__8079\ : InMux
    port map (
            O => \N__40973\,
            I => \N__40967\
        );

    \I__8078\ : Odrv4
    port map (
            O => \N__40970\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_20
        );

    \I__8077\ : LocalMux
    port map (
            O => \N__40967\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_20
        );

    \I__8076\ : CascadeMux
    port map (
            O => \N__40962\,
            I => \N__40958\
        );

    \I__8075\ : InMux
    port map (
            O => \N__40961\,
            I => \N__40954\
        );

    \I__8074\ : InMux
    port map (
            O => \N__40958\,
            I => \N__40949\
        );

    \I__8073\ : InMux
    port map (
            O => \N__40957\,
            I => \N__40949\
        );

    \I__8072\ : LocalMux
    port map (
            O => \N__40954\,
            I => \N__40946\
        );

    \I__8071\ : LocalMux
    port map (
            O => \N__40949\,
            I => \N__40943\
        );

    \I__8070\ : Span4Mux_v
    port map (
            O => \N__40946\,
            I => \N__40938\
        );

    \I__8069\ : Span4Mux_h
    port map (
            O => \N__40943\,
            I => \N__40938\
        );

    \I__8068\ : Odrv4
    port map (
            O => \N__40938\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_12
        );

    \I__8067\ : CascadeMux
    port map (
            O => \N__40935\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_0_12_cascade_\
        );

    \I__8066\ : InMux
    port map (
            O => \N__40932\,
            I => \N__40929\
        );

    \I__8065\ : LocalMux
    port map (
            O => \N__40929\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_2_12\
        );

    \I__8064\ : CascadeMux
    port map (
            O => \N__40926\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_0_i_12_cascade_\
        );

    \I__8063\ : InMux
    port map (
            O => \N__40923\,
            I => \N__40920\
        );

    \I__8062\ : LocalMux
    port map (
            O => \N__40920\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12\
        );

    \I__8061\ : CascadeMux
    port map (
            O => \N__40917\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12_cascade_\
        );

    \I__8060\ : InMux
    port map (
            O => \N__40914\,
            I => \N__40911\
        );

    \I__8059\ : LocalMux
    port map (
            O => \N__40911\,
            I => \N__40908\
        );

    \I__8058\ : Span4Mux_h
    port map (
            O => \N__40908\,
            I => \N__40905\
        );

    \I__8057\ : Span4Mux_v
    port map (
            O => \N__40905\,
            I => \N__40902\
        );

    \I__8056\ : Span4Mux_h
    port map (
            O => \N__40902\,
            I => \N__40899\
        );

    \I__8055\ : Odrv4
    port map (
            O => \N__40899\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_13\
        );

    \I__8054\ : CascadeMux
    port map (
            O => \N__40896\,
            I => \N__40893\
        );

    \I__8053\ : InMux
    port map (
            O => \N__40893\,
            I => \N__40889\
        );

    \I__8052\ : CascadeMux
    port map (
            O => \N__40892\,
            I => \N__40885\
        );

    \I__8051\ : LocalMux
    port map (
            O => \N__40889\,
            I => \N__40882\
        );

    \I__8050\ : InMux
    port map (
            O => \N__40888\,
            I => \N__40879\
        );

    \I__8049\ : InMux
    port map (
            O => \N__40885\,
            I => \N__40876\
        );

    \I__8048\ : Span4Mux_v
    port map (
            O => \N__40882\,
            I => \N__40871\
        );

    \I__8047\ : LocalMux
    port map (
            O => \N__40879\,
            I => \N__40871\
        );

    \I__8046\ : LocalMux
    port map (
            O => \N__40876\,
            I => \N__40868\
        );

    \I__8045\ : Span4Mux_h
    port map (
            O => \N__40871\,
            I => \N__40865\
        );

    \I__8044\ : Odrv12
    port map (
            O => \N__40868\,
            I => cemf_module_64ch_ctrl_inst1_data_config_13
        );

    \I__8043\ : Odrv4
    port map (
            O => \N__40865\,
            I => cemf_module_64ch_ctrl_inst1_data_config_13
        );

    \I__8042\ : CascadeMux
    port map (
            O => \N__40860\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8DZ0Z7_cascade_\
        );

    \I__8041\ : InMux
    port map (
            O => \N__40857\,
            I => \N__40854\
        );

    \I__8040\ : LocalMux
    port map (
            O => \N__40854\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13\
        );

    \I__8039\ : InMux
    port map (
            O => \N__40851\,
            I => \N__40848\
        );

    \I__8038\ : LocalMux
    port map (
            O => \N__40848\,
            I => \N__40845\
        );

    \I__8037\ : Odrv4
    port map (
            O => \N__40845\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8DZ0Z7\
        );

    \I__8036\ : InMux
    port map (
            O => \N__40842\,
            I => \N__40839\
        );

    \I__8035\ : LocalMux
    port map (
            O => \N__40839\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14\
        );

    \I__8034\ : CascadeMux
    port map (
            O => \N__40836\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14_cascade_\
        );

    \I__8033\ : InMux
    port map (
            O => \N__40833\,
            I => \N__40830\
        );

    \I__8032\ : LocalMux
    port map (
            O => \N__40830\,
            I => \N__40827\
        );

    \I__8031\ : Span4Mux_h
    port map (
            O => \N__40827\,
            I => \N__40824\
        );

    \I__8030\ : Span4Mux_v
    port map (
            O => \N__40824\,
            I => \N__40819\
        );

    \I__8029\ : InMux
    port map (
            O => \N__40823\,
            I => \N__40816\
        );

    \I__8028\ : InMux
    port map (
            O => \N__40822\,
            I => \N__40813\
        );

    \I__8027\ : Odrv4
    port map (
            O => \N__40819\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_8
        );

    \I__8026\ : LocalMux
    port map (
            O => \N__40816\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_8
        );

    \I__8025\ : LocalMux
    port map (
            O => \N__40813\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_8
        );

    \I__8024\ : InMux
    port map (
            O => \N__40806\,
            I => \N__40803\
        );

    \I__8023\ : LocalMux
    port map (
            O => \N__40803\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_8\
        );

    \I__8022\ : InMux
    port map (
            O => \N__40800\,
            I => \N__40797\
        );

    \I__8021\ : LocalMux
    port map (
            O => \N__40797\,
            I => \N__40794\
        );

    \I__8020\ : Odrv4
    port map (
            O => \N__40794\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_20\
        );

    \I__8019\ : InMux
    port map (
            O => \N__40791\,
            I => \N__40788\
        );

    \I__8018\ : LocalMux
    port map (
            O => \N__40788\,
            I => \N__40785\
        );

    \I__8017\ : Odrv12
    port map (
            O => \N__40785\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_3\
        );

    \I__8016\ : InMux
    port map (
            O => \N__40782\,
            I => \N__40779\
        );

    \I__8015\ : LocalMux
    port map (
            O => \N__40779\,
            I => \N__40776\
        );

    \I__8014\ : Odrv4
    port map (
            O => \N__40776\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_8\
        );

    \I__8013\ : CascadeMux
    port map (
            O => \N__40773\,
            I => \N__40770\
        );

    \I__8012\ : InMux
    port map (
            O => \N__40770\,
            I => \N__40767\
        );

    \I__8011\ : LocalMux
    port map (
            O => \N__40767\,
            I => \N__40763\
        );

    \I__8010\ : InMux
    port map (
            O => \N__40766\,
            I => \N__40760\
        );

    \I__8009\ : Span4Mux_v
    port map (
            O => \N__40763\,
            I => \N__40754\
        );

    \I__8008\ : LocalMux
    port map (
            O => \N__40760\,
            I => \N__40754\
        );

    \I__8007\ : InMux
    port map (
            O => \N__40759\,
            I => \N__40751\
        );

    \I__8006\ : Span4Mux_h
    port map (
            O => \N__40754\,
            I => \N__40748\
        );

    \I__8005\ : LocalMux
    port map (
            O => \N__40751\,
            I => \N__40745\
        );

    \I__8004\ : Span4Mux_v
    port map (
            O => \N__40748\,
            I => \N__40742\
        );

    \I__8003\ : Span4Mux_h
    port map (
            O => \N__40745\,
            I => \N__40739\
        );

    \I__8002\ : Sp12to4
    port map (
            O => \N__40742\,
            I => \N__40736\
        );

    \I__8001\ : Odrv4
    port map (
            O => \N__40739\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_8
        );

    \I__8000\ : Odrv12
    port map (
            O => \N__40736\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_8
        );

    \I__7999\ : InMux
    port map (
            O => \N__40731\,
            I => \N__40728\
        );

    \I__7998\ : LocalMux
    port map (
            O => \N__40728\,
            I => \N__40725\
        );

    \I__7997\ : Span4Mux_h
    port map (
            O => \N__40725\,
            I => \N__40722\
        );

    \I__7996\ : Span4Mux_h
    port map (
            O => \N__40722\,
            I => \N__40718\
        );

    \I__7995\ : InMux
    port map (
            O => \N__40721\,
            I => \N__40714\
        );

    \I__7994\ : Span4Mux_v
    port map (
            O => \N__40718\,
            I => \N__40711\
        );

    \I__7993\ : InMux
    port map (
            O => \N__40717\,
            I => \N__40708\
        );

    \I__7992\ : LocalMux
    port map (
            O => \N__40714\,
            I => \N__40705\
        );

    \I__7991\ : Odrv4
    port map (
            O => \N__40711\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_8
        );

    \I__7990\ : LocalMux
    port map (
            O => \N__40708\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_8
        );

    \I__7989\ : Odrv4
    port map (
            O => \N__40705\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_8
        );

    \I__7988\ : InMux
    port map (
            O => \N__40698\,
            I => \N__40693\
        );

    \I__7987\ : InMux
    port map (
            O => \N__40697\,
            I => \N__40690\
        );

    \I__7986\ : InMux
    port map (
            O => \N__40696\,
            I => \N__40687\
        );

    \I__7985\ : LocalMux
    port map (
            O => \N__40693\,
            I => \N__40684\
        );

    \I__7984\ : LocalMux
    port map (
            O => \N__40690\,
            I => \N__40681\
        );

    \I__7983\ : LocalMux
    port map (
            O => \N__40687\,
            I => \N__40678\
        );

    \I__7982\ : Span4Mux_h
    port map (
            O => \N__40684\,
            I => \N__40675\
        );

    \I__7981\ : Span4Mux_h
    port map (
            O => \N__40681\,
            I => \N__40672\
        );

    \I__7980\ : Span4Mux_h
    port map (
            O => \N__40678\,
            I => \N__40669\
        );

    \I__7979\ : Span4Mux_v
    port map (
            O => \N__40675\,
            I => \N__40666\
        );

    \I__7978\ : Span4Mux_h
    port map (
            O => \N__40672\,
            I => \N__40663\
        );

    \I__7977\ : Span4Mux_h
    port map (
            O => \N__40669\,
            I => \N__40660\
        );

    \I__7976\ : Odrv4
    port map (
            O => \N__40666\,
            I => cemf_module_64ch_ctrl_inst1_data_config_8
        );

    \I__7975\ : Odrv4
    port map (
            O => \N__40663\,
            I => cemf_module_64ch_ctrl_inst1_data_config_8
        );

    \I__7974\ : Odrv4
    port map (
            O => \N__40660\,
            I => cemf_module_64ch_ctrl_inst1_data_config_8
        );

    \I__7973\ : CascadeMux
    port map (
            O => \N__40653\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_8_cascade_\
        );

    \I__7972\ : CascadeMux
    port map (
            O => \N__40650\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SLZ0Z7_cascade_\
        );

    \I__7971\ : InMux
    port map (
            O => \N__40647\,
            I => \N__40644\
        );

    \I__7970\ : LocalMux
    port map (
            O => \N__40644\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8\
        );

    \I__7969\ : InMux
    port map (
            O => \N__40641\,
            I => \N__40638\
        );

    \I__7968\ : LocalMux
    port map (
            O => \N__40638\,
            I => \N__40635\
        );

    \I__7967\ : Span4Mux_v
    port map (
            O => \N__40635\,
            I => \N__40632\
        );

    \I__7966\ : Span4Mux_h
    port map (
            O => \N__40632\,
            I => \N__40629\
        );

    \I__7965\ : Odrv4
    port map (
            O => \N__40629\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_7\
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__40626\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8_cascade_\
        );

    \I__7963\ : CascadeMux
    port map (
            O => \N__40623\,
            I => \N__40620\
        );

    \I__7962\ : InMux
    port map (
            O => \N__40620\,
            I => \N__40617\
        );

    \I__7961\ : LocalMux
    port map (
            O => \N__40617\,
            I => \N__40614\
        );

    \I__7960\ : Span4Mux_h
    port map (
            O => \N__40614\,
            I => \N__40611\
        );

    \I__7959\ : Span4Mux_h
    port map (
            O => \N__40611\,
            I => \N__40608\
        );

    \I__7958\ : Sp12to4
    port map (
            O => \N__40608\,
            I => \N__40605\
        );

    \I__7957\ : Odrv12
    port map (
            O => \N__40605\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_28\
        );

    \I__7956\ : InMux
    port map (
            O => \N__40602\,
            I => \N__40599\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__40599\,
            I => \N__40596\
        );

    \I__7954\ : Span4Mux_v
    port map (
            O => \N__40596\,
            I => \N__40593\
        );

    \I__7953\ : Span4Mux_v
    port map (
            O => \N__40593\,
            I => \N__40590\
        );

    \I__7952\ : Sp12to4
    port map (
            O => \N__40590\,
            I => \N__40587\
        );

    \I__7951\ : Odrv12
    port map (
            O => \N__40587\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_1Z0Z_26\
        );

    \I__7950\ : CascadeMux
    port map (
            O => \N__40584\,
            I => \N__40581\
        );

    \I__7949\ : InMux
    port map (
            O => \N__40581\,
            I => \N__40578\
        );

    \I__7948\ : LocalMux
    port map (
            O => \N__40578\,
            I => \N__40575\
        );

    \I__7947\ : Span4Mux_h
    port map (
            O => \N__40575\,
            I => \N__40572\
        );

    \I__7946\ : Odrv4
    port map (
            O => \N__40572\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_27\
        );

    \I__7945\ : InMux
    port map (
            O => \N__40569\,
            I => \N__40566\
        );

    \I__7944\ : LocalMux
    port map (
            O => \N__40566\,
            I => \N__40563\
        );

    \I__7943\ : Odrv4
    port map (
            O => \N__40563\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_7\
        );

    \I__7942\ : InMux
    port map (
            O => \N__40560\,
            I => \N__40557\
        );

    \I__7941\ : LocalMux
    port map (
            O => \N__40557\,
            I => \N__40554\
        );

    \I__7940\ : Odrv12
    port map (
            O => \N__40554\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_7\
        );

    \I__7939\ : InMux
    port map (
            O => \N__40551\,
            I => \N__40548\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__40548\,
            I => \N__40545\
        );

    \I__7937\ : Span12Mux_h
    port map (
            O => \N__40545\,
            I => \N__40540\
        );

    \I__7936\ : InMux
    port map (
            O => \N__40544\,
            I => \N__40535\
        );

    \I__7935\ : InMux
    port map (
            O => \N__40543\,
            I => \N__40535\
        );

    \I__7934\ : Odrv12
    port map (
            O => \N__40540\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_7
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__40535\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_7
        );

    \I__7932\ : CascadeMux
    port map (
            O => \N__40530\,
            I => \N__40526\
        );

    \I__7931\ : InMux
    port map (
            O => \N__40529\,
            I => \N__40523\
        );

    \I__7930\ : InMux
    port map (
            O => \N__40526\,
            I => \N__40520\
        );

    \I__7929\ : LocalMux
    port map (
            O => \N__40523\,
            I => \N__40517\
        );

    \I__7928\ : LocalMux
    port map (
            O => \N__40520\,
            I => \N__40514\
        );

    \I__7927\ : Span4Mux_h
    port map (
            O => \N__40517\,
            I => \N__40511\
        );

    \I__7926\ : Span4Mux_h
    port map (
            O => \N__40514\,
            I => \N__40507\
        );

    \I__7925\ : Span4Mux_h
    port map (
            O => \N__40511\,
            I => \N__40504\
        );

    \I__7924\ : InMux
    port map (
            O => \N__40510\,
            I => \N__40501\
        );

    \I__7923\ : Span4Mux_h
    port map (
            O => \N__40507\,
            I => \N__40498\
        );

    \I__7922\ : Odrv4
    port map (
            O => \N__40504\,
            I => cemf_module_64ch_ctrl_inst1_data_config_7
        );

    \I__7921\ : LocalMux
    port map (
            O => \N__40501\,
            I => cemf_module_64ch_ctrl_inst1_data_config_7
        );

    \I__7920\ : Odrv4
    port map (
            O => \N__40498\,
            I => cemf_module_64ch_ctrl_inst1_data_config_7
        );

    \I__7919\ : CascadeMux
    port map (
            O => \N__40491\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_8_cascade_\
        );

    \I__7918\ : CascadeMux
    port map (
            O => \N__40488\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3QZ0Z5_cascade_\
        );

    \I__7917\ : InMux
    port map (
            O => \N__40485\,
            I => \N__40482\
        );

    \I__7916\ : LocalMux
    port map (
            O => \N__40482\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__40479\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8_cascade_\
        );

    \I__7914\ : CascadeMux
    port map (
            O => \N__40476\,
            I => \N__40473\
        );

    \I__7913\ : InMux
    port map (
            O => \N__40473\,
            I => \N__40470\
        );

    \I__7912\ : LocalMux
    port map (
            O => \N__40470\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_7\
        );

    \I__7911\ : CascadeMux
    port map (
            O => \N__40467\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3QZ0Z5_cascade_\
        );

    \I__7910\ : InMux
    port map (
            O => \N__40464\,
            I => \N__40461\
        );

    \I__7909\ : LocalMux
    port map (
            O => \N__40461\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7\
        );

    \I__7908\ : InMux
    port map (
            O => \N__40458\,
            I => \N__40455\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__40455\,
            I => \N__40452\
        );

    \I__7906\ : Span12Mux_v
    port map (
            O => \N__40452\,
            I => \N__40449\
        );

    \I__7905\ : Odrv12
    port map (
            O => \N__40449\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_6\
        );

    \I__7904\ : CascadeMux
    port map (
            O => \N__40446\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7_cascade_\
        );

    \I__7903\ : InMux
    port map (
            O => \N__40443\,
            I => \N__40440\
        );

    \I__7902\ : LocalMux
    port map (
            O => \N__40440\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_7\
        );

    \I__7901\ : CascadeMux
    port map (
            O => \N__40437\,
            I => \N__40434\
        );

    \I__7900\ : InMux
    port map (
            O => \N__40434\,
            I => \N__40431\
        );

    \I__7899\ : LocalMux
    port map (
            O => \N__40431\,
            I => \N__40428\
        );

    \I__7898\ : Span4Mux_v
    port map (
            O => \N__40428\,
            I => \N__40425\
        );

    \I__7897\ : Odrv4
    port map (
            O => \N__40425\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_24\
        );

    \I__7896\ : InMux
    port map (
            O => \N__40422\,
            I => \N__40419\
        );

    \I__7895\ : LocalMux
    port map (
            O => \N__40419\,
            I => \N__40416\
        );

    \I__7894\ : Odrv4
    port map (
            O => \N__40416\,
            I => \serializer_mod_inst.shift_regZ0Z_82\
        );

    \I__7893\ : InMux
    port map (
            O => \N__40413\,
            I => \N__40410\
        );

    \I__7892\ : LocalMux
    port map (
            O => \N__40410\,
            I => \N__40407\
        );

    \I__7891\ : Span4Mux_h
    port map (
            O => \N__40407\,
            I => \N__40404\
        );

    \I__7890\ : Odrv4
    port map (
            O => \N__40404\,
            I => \serializer_mod_inst.shift_regZ0Z_80\
        );

    \I__7889\ : InMux
    port map (
            O => \N__40401\,
            I => \N__40398\
        );

    \I__7888\ : LocalMux
    port map (
            O => \N__40398\,
            I => \serializer_mod_inst.shift_regZ0Z_81\
        );

    \I__7887\ : InMux
    port map (
            O => \N__40395\,
            I => \N__40392\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__40392\,
            I => \N__40389\
        );

    \I__7885\ : Span4Mux_v
    port map (
            O => \N__40389\,
            I => \N__40386\
        );

    \I__7884\ : Span4Mux_h
    port map (
            O => \N__40386\,
            I => \N__40383\
        );

    \I__7883\ : Span4Mux_h
    port map (
            O => \N__40383\,
            I => \N__40380\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__40380\,
            I => \N__40377\
        );

    \I__7881\ : Odrv4
    port map (
            O => \N__40377\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_29
        );

    \I__7880\ : CascadeMux
    port map (
            O => \N__40374\,
            I => \N__40371\
        );

    \I__7879\ : InMux
    port map (
            O => \N__40371\,
            I => \N__40368\
        );

    \I__7878\ : LocalMux
    port map (
            O => \N__40368\,
            I => \N__40365\
        );

    \I__7877\ : Span4Mux_v
    port map (
            O => \N__40365\,
            I => \N__40362\
        );

    \I__7876\ : Span4Mux_h
    port map (
            O => \N__40362\,
            I => \N__40359\
        );

    \I__7875\ : Span4Mux_h
    port map (
            O => \N__40359\,
            I => \N__40356\
        );

    \I__7874\ : Odrv4
    port map (
            O => \N__40356\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_29
        );

    \I__7873\ : CascadeMux
    port map (
            O => \N__40353\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_29_cascade_\
        );

    \I__7872\ : InMux
    port map (
            O => \N__40350\,
            I => \N__40347\
        );

    \I__7871\ : LocalMux
    port map (
            O => \N__40347\,
            I => \N__40344\
        );

    \I__7870\ : Span4Mux_v
    port map (
            O => \N__40344\,
            I => \N__40341\
        );

    \I__7869\ : Span4Mux_h
    port map (
            O => \N__40341\,
            I => \N__40338\
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__40338\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_29\
        );

    \I__7867\ : InMux
    port map (
            O => \N__40335\,
            I => \N__40332\
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__40332\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_29\
        );

    \I__7865\ : CascadeMux
    port map (
            O => \N__40329\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_29_cascade_\
        );

    \I__7864\ : InMux
    port map (
            O => \N__40326\,
            I => \N__40323\
        );

    \I__7863\ : LocalMux
    port map (
            O => \N__40323\,
            I => \N__40320\
        );

    \I__7862\ : Span4Mux_h
    port map (
            O => \N__40320\,
            I => \N__40317\
        );

    \I__7861\ : Span4Mux_h
    port map (
            O => \N__40317\,
            I => \N__40314\
        );

    \I__7860\ : Odrv4
    port map (
            O => \N__40314\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_632\
        );

    \I__7859\ : InMux
    port map (
            O => \N__40311\,
            I => \N__40308\
        );

    \I__7858\ : LocalMux
    port map (
            O => \N__40308\,
            I => \N__40305\
        );

    \I__7857\ : Span4Mux_h
    port map (
            O => \N__40305\,
            I => \N__40302\
        );

    \I__7856\ : Span4Mux_h
    port map (
            O => \N__40302\,
            I => \N__40299\
        );

    \I__7855\ : Odrv4
    port map (
            O => \N__40299\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_29\
        );

    \I__7854\ : InMux
    port map (
            O => \N__40296\,
            I => \N__40293\
        );

    \I__7853\ : LocalMux
    port map (
            O => \N__40293\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_29\
        );

    \I__7852\ : InMux
    port map (
            O => \N__40290\,
            I => \N__40287\
        );

    \I__7851\ : LocalMux
    port map (
            O => \N__40287\,
            I => \serializer_mod_inst.shift_regZ0Z_42\
        );

    \I__7850\ : InMux
    port map (
            O => \N__40284\,
            I => \N__40281\
        );

    \I__7849\ : LocalMux
    port map (
            O => \N__40281\,
            I => \serializer_mod_inst.shift_regZ0Z_43\
        );

    \I__7848\ : InMux
    port map (
            O => \N__40278\,
            I => \N__40275\
        );

    \I__7847\ : LocalMux
    port map (
            O => \N__40275\,
            I => \serializer_mod_inst.shift_regZ0Z_44\
        );

    \I__7846\ : InMux
    port map (
            O => \N__40272\,
            I => \N__40269\
        );

    \I__7845\ : LocalMux
    port map (
            O => \N__40269\,
            I => \N__40266\
        );

    \I__7844\ : Odrv4
    port map (
            O => \N__40266\,
            I => \serializer_mod_inst.shift_regZ0Z_45\
        );

    \I__7843\ : InMux
    port map (
            O => \N__40263\,
            I => \N__40260\
        );

    \I__7842\ : LocalMux
    port map (
            O => \N__40260\,
            I => \serializer_mod_inst.shift_regZ0Z_70\
        );

    \I__7841\ : InMux
    port map (
            O => \N__40257\,
            I => \N__40254\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__40254\,
            I => \serializer_mod_inst.shift_regZ0Z_71\
        );

    \I__7839\ : InMux
    port map (
            O => \N__40251\,
            I => \N__40248\
        );

    \I__7838\ : LocalMux
    port map (
            O => \N__40248\,
            I => \serializer_mod_inst.shift_regZ0Z_74\
        );

    \I__7837\ : InMux
    port map (
            O => \N__40245\,
            I => \N__40242\
        );

    \I__7836\ : LocalMux
    port map (
            O => \N__40242\,
            I => \N__40239\
        );

    \I__7835\ : Odrv4
    port map (
            O => \N__40239\,
            I => \serializer_mod_inst.shift_regZ0Z_75\
        );

    \I__7834\ : InMux
    port map (
            O => \N__40236\,
            I => \N__40233\
        );

    \I__7833\ : LocalMux
    port map (
            O => \N__40233\,
            I => \N__40230\
        );

    \I__7832\ : Odrv4
    port map (
            O => \N__40230\,
            I => \serializer_mod_inst.shift_regZ0Z_98\
        );

    \I__7831\ : InMux
    port map (
            O => \N__40227\,
            I => \N__40224\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__40224\,
            I => \N__40221\
        );

    \I__7829\ : Odrv4
    port map (
            O => \N__40221\,
            I => \serializer_mod_inst.shift_regZ0Z_99\
        );

    \I__7828\ : InMux
    port map (
            O => \N__40218\,
            I => \N__40215\
        );

    \I__7827\ : LocalMux
    port map (
            O => \N__40215\,
            I => \serializer_mod_inst.shift_regZ0Z_72\
        );

    \I__7826\ : InMux
    port map (
            O => \N__40212\,
            I => \N__40209\
        );

    \I__7825\ : LocalMux
    port map (
            O => \N__40209\,
            I => \serializer_mod_inst.shift_regZ0Z_73\
        );

    \I__7824\ : CascadeMux
    port map (
            O => \N__40206\,
            I => \N__40203\
        );

    \I__7823\ : InMux
    port map (
            O => \N__40203\,
            I => \N__40200\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__40200\,
            I => \serializer_mod_inst.shift_regZ0Z_83\
        );

    \I__7821\ : InMux
    port map (
            O => \N__40197\,
            I => \N__40194\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__40194\,
            I => \N__40191\
        );

    \I__7819\ : Odrv4
    port map (
            O => \N__40191\,
            I => \serializer_mod_inst.shift_regZ0Z_85\
        );

    \I__7818\ : InMux
    port map (
            O => \N__40188\,
            I => \N__40185\
        );

    \I__7817\ : LocalMux
    port map (
            O => \N__40185\,
            I => \serializer_mod_inst.shift_regZ0Z_1\
        );

    \I__7816\ : InMux
    port map (
            O => \N__40182\,
            I => \N__40179\
        );

    \I__7815\ : LocalMux
    port map (
            O => \N__40179\,
            I => \serializer_mod_inst.shift_regZ0Z_101\
        );

    \I__7814\ : InMux
    port map (
            O => \N__40176\,
            I => \N__40173\
        );

    \I__7813\ : LocalMux
    port map (
            O => \N__40173\,
            I => \N__40170\
        );

    \I__7812\ : Span4Mux_h
    port map (
            O => \N__40170\,
            I => \N__40167\
        );

    \I__7811\ : Odrv4
    port map (
            O => \N__40167\,
            I => \serializer_mod_inst.shift_regZ0Z_66\
        );

    \I__7810\ : InMux
    port map (
            O => \N__40164\,
            I => \N__40161\
        );

    \I__7809\ : LocalMux
    port map (
            O => \N__40161\,
            I => \serializer_mod_inst.shift_regZ0Z_102\
        );

    \I__7808\ : CascadeMux
    port map (
            O => \N__40158\,
            I => \N__40155\
        );

    \I__7807\ : InMux
    port map (
            O => \N__40155\,
            I => \N__40152\
        );

    \I__7806\ : LocalMux
    port map (
            O => \N__40152\,
            I => \N__40149\
        );

    \I__7805\ : Odrv4
    port map (
            O => \N__40149\,
            I => \serializer_mod_inst.shift_regZ0Z_103\
        );

    \I__7804\ : InMux
    port map (
            O => \N__40146\,
            I => \N__40143\
        );

    \I__7803\ : LocalMux
    port map (
            O => \N__40143\,
            I => \serializer_mod_inst.shift_regZ0Z_84\
        );

    \I__7802\ : InMux
    port map (
            O => \N__40140\,
            I => \N__40137\
        );

    \I__7801\ : LocalMux
    port map (
            O => \N__40137\,
            I => \N__40134\
        );

    \I__7800\ : Odrv12
    port map (
            O => \N__40134\,
            I => \serializer_mod_inst.shift_regZ0Z_41\
        );

    \I__7799\ : InMux
    port map (
            O => \N__40131\,
            I => \N__40128\
        );

    \I__7798\ : LocalMux
    port map (
            O => \N__40128\,
            I => \N__40125\
        );

    \I__7797\ : Odrv4
    port map (
            O => \N__40125\,
            I => \serializer_mod_inst.shift_regZ0Z_100\
        );

    \I__7796\ : InMux
    port map (
            O => \N__40122\,
            I => \N__40119\
        );

    \I__7795\ : LocalMux
    port map (
            O => \N__40119\,
            I => \N__40116\
        );

    \I__7794\ : Odrv4
    port map (
            O => \N__40116\,
            I => \serializer_mod_inst.shift_regZ0Z_54\
        );

    \I__7793\ : InMux
    port map (
            O => \N__40113\,
            I => \N__40108\
        );

    \I__7792\ : InMux
    port map (
            O => \N__40112\,
            I => \N__40105\
        );

    \I__7791\ : InMux
    port map (
            O => \N__40111\,
            I => \N__40102\
        );

    \I__7790\ : LocalMux
    port map (
            O => \N__40108\,
            I => \N__40099\
        );

    \I__7789\ : LocalMux
    port map (
            O => \N__40105\,
            I => \N__40093\
        );

    \I__7788\ : LocalMux
    port map (
            O => \N__40102\,
            I => \N__40090\
        );

    \I__7787\ : Span4Mux_h
    port map (
            O => \N__40099\,
            I => \N__40087\
        );

    \I__7786\ : InMux
    port map (
            O => \N__40098\,
            I => \N__40080\
        );

    \I__7785\ : InMux
    port map (
            O => \N__40097\,
            I => \N__40080\
        );

    \I__7784\ : InMux
    port map (
            O => \N__40096\,
            I => \N__40080\
        );

    \I__7783\ : Span4Mux_v
    port map (
            O => \N__40093\,
            I => \N__40077\
        );

    \I__7782\ : Span4Mux_v
    port map (
            O => \N__40090\,
            I => \N__40074\
        );

    \I__7781\ : Span4Mux_v
    port map (
            O => \N__40087\,
            I => \N__40069\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__40080\,
            I => \N__40069\
        );

    \I__7779\ : Sp12to4
    port map (
            O => \N__40077\,
            I => \N__40064\
        );

    \I__7778\ : Sp12to4
    port map (
            O => \N__40074\,
            I => \N__40064\
        );

    \I__7777\ : Span4Mux_h
    port map (
            O => \N__40069\,
            I => \N__40061\
        );

    \I__7776\ : Span12Mux_h
    port map (
            O => \N__40064\,
            I => \N__40056\
        );

    \I__7775\ : Span4Mux_h
    port map (
            O => \N__40061\,
            I => \N__40053\
        );

    \I__7774\ : InMux
    port map (
            O => \N__40060\,
            I => \N__40048\
        );

    \I__7773\ : InMux
    port map (
            O => \N__40059\,
            I => \N__40048\
        );

    \I__7772\ : Odrv12
    port map (
            O => \N__40056\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_0
        );

    \I__7771\ : Odrv4
    port map (
            O => \N__40053\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_0
        );

    \I__7770\ : LocalMux
    port map (
            O => \N__40048\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_0
        );

    \I__7769\ : InMux
    port map (
            O => \N__40041\,
            I => \N__40038\
        );

    \I__7768\ : LocalMux
    port map (
            O => \N__40038\,
            I => \N__40034\
        );

    \I__7767\ : InMux
    port map (
            O => \N__40037\,
            I => \N__40030\
        );

    \I__7766\ : Span4Mux_h
    port map (
            O => \N__40034\,
            I => \N__40027\
        );

    \I__7765\ : InMux
    port map (
            O => \N__40033\,
            I => \N__40024\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__40030\,
            I => \N__40021\
        );

    \I__7763\ : Span4Mux_v
    port map (
            O => \N__40027\,
            I => \N__40018\
        );

    \I__7762\ : LocalMux
    port map (
            O => \N__40024\,
            I => \N__40015\
        );

    \I__7761\ : Span4Mux_h
    port map (
            O => \N__40021\,
            I => \N__40012\
        );

    \I__7760\ : Span4Mux_v
    port map (
            O => \N__40018\,
            I => \N__40009\
        );

    \I__7759\ : Odrv4
    port map (
            O => \N__40015\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0\
        );

    \I__7758\ : Odrv4
    port map (
            O => \N__40012\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0\
        );

    \I__7757\ : Odrv4
    port map (
            O => \N__40009\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0\
        );

    \I__7756\ : InMux
    port map (
            O => \N__40002\,
            I => \N__39997\
        );

    \I__7755\ : InMux
    port map (
            O => \N__40001\,
            I => \N__39994\
        );

    \I__7754\ : InMux
    port map (
            O => \N__40000\,
            I => \N__39991\
        );

    \I__7753\ : LocalMux
    port map (
            O => \N__39997\,
            I => \N__39988\
        );

    \I__7752\ : LocalMux
    port map (
            O => \N__39994\,
            I => \N__39985\
        );

    \I__7751\ : LocalMux
    port map (
            O => \N__39991\,
            I => \N__39982\
        );

    \I__7750\ : Span4Mux_v
    port map (
            O => \N__39988\,
            I => \N__39979\
        );

    \I__7749\ : Span4Mux_h
    port map (
            O => \N__39985\,
            I => \N__39976\
        );

    \I__7748\ : Span12Mux_h
    port map (
            O => \N__39982\,
            I => \N__39971\
        );

    \I__7747\ : Sp12to4
    port map (
            O => \N__39979\,
            I => \N__39971\
        );

    \I__7746\ : Odrv4
    port map (
            O => \N__39976\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6\
        );

    \I__7745\ : Odrv12
    port map (
            O => \N__39971\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6\
        );

    \I__7744\ : CascadeMux
    port map (
            O => \N__39966\,
            I => \N__39963\
        );

    \I__7743\ : InMux
    port map (
            O => \N__39963\,
            I => \N__39960\
        );

    \I__7742\ : LocalMux
    port map (
            O => \N__39960\,
            I => \serializer_mod_inst.shift_regZ0Z_52\
        );

    \I__7741\ : InMux
    port map (
            O => \N__39957\,
            I => \N__39954\
        );

    \I__7740\ : LocalMux
    port map (
            O => \N__39954\,
            I => \serializer_mod_inst.shift_regZ0Z_53\
        );

    \I__7739\ : CascadeMux
    port map (
            O => \N__39951\,
            I => \N__39948\
        );

    \I__7738\ : InMux
    port map (
            O => \N__39948\,
            I => \N__39945\
        );

    \I__7737\ : LocalMux
    port map (
            O => \N__39945\,
            I => \serializer_mod_inst.shift_regZ0Z_87\
        );

    \I__7736\ : InMux
    port map (
            O => \N__39942\,
            I => \N__39939\
        );

    \I__7735\ : LocalMux
    port map (
            O => \N__39939\,
            I => \serializer_mod_inst.shift_regZ0Z_88\
        );

    \I__7734\ : InMux
    port map (
            O => \N__39936\,
            I => \N__39933\
        );

    \I__7733\ : LocalMux
    port map (
            O => \N__39933\,
            I => \serializer_mod_inst.shift_regZ0Z_49\
        );

    \I__7732\ : CascadeMux
    port map (
            O => \N__39930\,
            I => \N__39927\
        );

    \I__7731\ : InMux
    port map (
            O => \N__39927\,
            I => \N__39924\
        );

    \I__7730\ : LocalMux
    port map (
            O => \N__39924\,
            I => \serializer_mod_inst.shift_regZ0Z_50\
        );

    \I__7729\ : InMux
    port map (
            O => \N__39921\,
            I => \N__39918\
        );

    \I__7728\ : LocalMux
    port map (
            O => \N__39918\,
            I => \serializer_mod_inst.shift_regZ0Z_89\
        );

    \I__7727\ : InMux
    port map (
            O => \N__39915\,
            I => \N__39912\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__39912\,
            I => \serializer_mod_inst.shift_regZ0Z_90\
        );

    \I__7725\ : InMux
    port map (
            O => \N__39909\,
            I => \N__39905\
        );

    \I__7724\ : InMux
    port map (
            O => \N__39908\,
            I => \N__39902\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__39905\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_9
        );

    \I__7722\ : LocalMux
    port map (
            O => \N__39902\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_9
        );

    \I__7721\ : InMux
    port map (
            O => \N__39897\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8\
        );

    \I__7720\ : InMux
    port map (
            O => \N__39894\,
            I => \N__39890\
        );

    \I__7719\ : InMux
    port map (
            O => \N__39893\,
            I => \N__39887\
        );

    \I__7718\ : LocalMux
    port map (
            O => \N__39890\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_10
        );

    \I__7717\ : LocalMux
    port map (
            O => \N__39887\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_10
        );

    \I__7716\ : InMux
    port map (
            O => \N__39882\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9\
        );

    \I__7715\ : InMux
    port map (
            O => \N__39879\,
            I => \N__39875\
        );

    \I__7714\ : InMux
    port map (
            O => \N__39878\,
            I => \N__39872\
        );

    \I__7713\ : LocalMux
    port map (
            O => \N__39875\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_11
        );

    \I__7712\ : LocalMux
    port map (
            O => \N__39872\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_11
        );

    \I__7711\ : InMux
    port map (
            O => \N__39867\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10\
        );

    \I__7710\ : InMux
    port map (
            O => \N__39864\,
            I => \N__39860\
        );

    \I__7709\ : InMux
    port map (
            O => \N__39863\,
            I => \N__39857\
        );

    \I__7708\ : LocalMux
    port map (
            O => \N__39860\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_12
        );

    \I__7707\ : LocalMux
    port map (
            O => \N__39857\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_12
        );

    \I__7706\ : InMux
    port map (
            O => \N__39852\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11\
        );

    \I__7705\ : InMux
    port map (
            O => \N__39849\,
            I => \N__39845\
        );

    \I__7704\ : InMux
    port map (
            O => \N__39848\,
            I => \N__39842\
        );

    \I__7703\ : LocalMux
    port map (
            O => \N__39845\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_13
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__39842\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_13
        );

    \I__7701\ : InMux
    port map (
            O => \N__39837\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12\
        );

    \I__7700\ : CascadeMux
    port map (
            O => \N__39834\,
            I => \N__39830\
        );

    \I__7699\ : InMux
    port map (
            O => \N__39833\,
            I => \N__39827\
        );

    \I__7698\ : InMux
    port map (
            O => \N__39830\,
            I => \N__39824\
        );

    \I__7697\ : LocalMux
    port map (
            O => \N__39827\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_14
        );

    \I__7696\ : LocalMux
    port map (
            O => \N__39824\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_14
        );

    \I__7695\ : InMux
    port map (
            O => \N__39819\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13\
        );

    \I__7694\ : InMux
    port map (
            O => \N__39816\,
            I => \N__39800\
        );

    \I__7693\ : InMux
    port map (
            O => \N__39815\,
            I => \N__39800\
        );

    \I__7692\ : InMux
    port map (
            O => \N__39814\,
            I => \N__39800\
        );

    \I__7691\ : InMux
    port map (
            O => \N__39813\,
            I => \N__39800\
        );

    \I__7690\ : InMux
    port map (
            O => \N__39812\,
            I => \N__39782\
        );

    \I__7689\ : InMux
    port map (
            O => \N__39811\,
            I => \N__39782\
        );

    \I__7688\ : InMux
    port map (
            O => \N__39810\,
            I => \N__39782\
        );

    \I__7687\ : InMux
    port map (
            O => \N__39809\,
            I => \N__39782\
        );

    \I__7686\ : LocalMux
    port map (
            O => \N__39800\,
            I => \N__39779\
        );

    \I__7685\ : InMux
    port map (
            O => \N__39799\,
            I => \N__39770\
        );

    \I__7684\ : InMux
    port map (
            O => \N__39798\,
            I => \N__39770\
        );

    \I__7683\ : InMux
    port map (
            O => \N__39797\,
            I => \N__39770\
        );

    \I__7682\ : InMux
    port map (
            O => \N__39796\,
            I => \N__39770\
        );

    \I__7681\ : InMux
    port map (
            O => \N__39795\,
            I => \N__39761\
        );

    \I__7680\ : InMux
    port map (
            O => \N__39794\,
            I => \N__39761\
        );

    \I__7679\ : InMux
    port map (
            O => \N__39793\,
            I => \N__39761\
        );

    \I__7678\ : InMux
    port map (
            O => \N__39792\,
            I => \N__39761\
        );

    \I__7677\ : InMux
    port map (
            O => \N__39791\,
            I => \N__39758\
        );

    \I__7676\ : LocalMux
    port map (
            O => \N__39782\,
            I => \N__39754\
        );

    \I__7675\ : Span4Mux_v
    port map (
            O => \N__39779\,
            I => \N__39747\
        );

    \I__7674\ : LocalMux
    port map (
            O => \N__39770\,
            I => \N__39747\
        );

    \I__7673\ : LocalMux
    port map (
            O => \N__39761\,
            I => \N__39747\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__39758\,
            I => \N__39744\
        );

    \I__7671\ : InMux
    port map (
            O => \N__39757\,
            I => \N__39739\
        );

    \I__7670\ : Span4Mux_h
    port map (
            O => \N__39754\,
            I => \N__39736\
        );

    \I__7669\ : Span4Mux_h
    port map (
            O => \N__39747\,
            I => \N__39733\
        );

    \I__7668\ : Span12Mux_v
    port map (
            O => \N__39744\,
            I => \N__39730\
        );

    \I__7667\ : InMux
    port map (
            O => \N__39743\,
            I => \N__39725\
        );

    \I__7666\ : InMux
    port map (
            O => \N__39742\,
            I => \N__39725\
        );

    \I__7665\ : LocalMux
    port map (
            O => \N__39739\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\
        );

    \I__7664\ : Odrv4
    port map (
            O => \N__39736\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\
        );

    \I__7663\ : Odrv4
    port map (
            O => \N__39733\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\
        );

    \I__7662\ : Odrv12
    port map (
            O => \N__39730\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__39725\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\
        );

    \I__7660\ : InMux
    port map (
            O => \N__39714\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_14\
        );

    \I__7659\ : CascadeMux
    port map (
            O => \N__39711\,
            I => \N__39707\
        );

    \I__7658\ : InMux
    port map (
            O => \N__39710\,
            I => \N__39704\
        );

    \I__7657\ : InMux
    port map (
            O => \N__39707\,
            I => \N__39701\
        );

    \I__7656\ : LocalMux
    port map (
            O => \N__39704\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_15
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__39701\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_15
        );

    \I__7654\ : CEMux
    port map (
            O => \N__39696\,
            I => \N__39692\
        );

    \I__7653\ : CEMux
    port map (
            O => \N__39695\,
            I => \N__39689\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__39692\,
            I => \N__39686\
        );

    \I__7651\ : LocalMux
    port map (
            O => \N__39689\,
            I => \N__39683\
        );

    \I__7650\ : Span4Mux_h
    port map (
            O => \N__39686\,
            I => \N__39680\
        );

    \I__7649\ : Span4Mux_h
    port map (
            O => \N__39683\,
            I => \N__39677\
        );

    \I__7648\ : Span4Mux_h
    port map (
            O => \N__39680\,
            I => \N__39674\
        );

    \I__7647\ : Span4Mux_h
    port map (
            O => \N__39677\,
            I => \N__39671\
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__39674\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0\
        );

    \I__7645\ : Odrv4
    port map (
            O => \N__39671\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0\
        );

    \I__7644\ : InMux
    port map (
            O => \N__39666\,
            I => \N__39663\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__39663\,
            I => \serializer_mod_inst.shift_regZ0Z_86\
        );

    \I__7642\ : CascadeMux
    port map (
            O => \N__39660\,
            I => \N__39657\
        );

    \I__7641\ : InMux
    port map (
            O => \N__39657\,
            I => \N__39654\
        );

    \I__7640\ : LocalMux
    port map (
            O => \N__39654\,
            I => \N__39650\
        );

    \I__7639\ : InMux
    port map (
            O => \N__39653\,
            I => \N__39647\
        );

    \I__7638\ : Span4Mux_h
    port map (
            O => \N__39650\,
            I => \N__39643\
        );

    \I__7637\ : LocalMux
    port map (
            O => \N__39647\,
            I => \N__39640\
        );

    \I__7636\ : InMux
    port map (
            O => \N__39646\,
            I => \N__39637\
        );

    \I__7635\ : Span4Mux_v
    port map (
            O => \N__39643\,
            I => \N__39634\
        );

    \I__7634\ : Span12Mux_v
    port map (
            O => \N__39640\,
            I => \N__39631\
        );

    \I__7633\ : LocalMux
    port map (
            O => \N__39637\,
            I => \cemf_module_64ch_ctrl_inst1.paddr_fsm_1\
        );

    \I__7632\ : Odrv4
    port map (
            O => \N__39634\,
            I => \cemf_module_64ch_ctrl_inst1.paddr_fsm_1\
        );

    \I__7631\ : Odrv12
    port map (
            O => \N__39631\,
            I => \cemf_module_64ch_ctrl_inst1.paddr_fsm_1\
        );

    \I__7630\ : InMux
    port map (
            O => \N__39624\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0\
        );

    \I__7629\ : InMux
    port map (
            O => \N__39621\,
            I => \N__39618\
        );

    \I__7628\ : LocalMux
    port map (
            O => \N__39618\,
            I => \N__39614\
        );

    \I__7627\ : CascadeMux
    port map (
            O => \N__39617\,
            I => \N__39608\
        );

    \I__7626\ : Span4Mux_h
    port map (
            O => \N__39614\,
            I => \N__39605\
        );

    \I__7625\ : InMux
    port map (
            O => \N__39613\,
            I => \N__39596\
        );

    \I__7624\ : InMux
    port map (
            O => \N__39612\,
            I => \N__39596\
        );

    \I__7623\ : InMux
    port map (
            O => \N__39611\,
            I => \N__39596\
        );

    \I__7622\ : InMux
    port map (
            O => \N__39608\,
            I => \N__39596\
        );

    \I__7621\ : Span4Mux_h
    port map (
            O => \N__39605\,
            I => \N__39590\
        );

    \I__7620\ : LocalMux
    port map (
            O => \N__39596\,
            I => \N__39590\
        );

    \I__7619\ : InMux
    port map (
            O => \N__39595\,
            I => \N__39587\
        );

    \I__7618\ : Span4Mux_h
    port map (
            O => \N__39590\,
            I => \N__39584\
        );

    \I__7617\ : LocalMux
    port map (
            O => \N__39587\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_2
        );

    \I__7616\ : Odrv4
    port map (
            O => \N__39584\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_2
        );

    \I__7615\ : InMux
    port map (
            O => \N__39579\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1\
        );

    \I__7614\ : InMux
    port map (
            O => \N__39576\,
            I => \N__39573\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__39573\,
            I => \N__39570\
        );

    \I__7612\ : Span4Mux_h
    port map (
            O => \N__39570\,
            I => \N__39567\
        );

    \I__7611\ : Span4Mux_h
    port map (
            O => \N__39567\,
            I => \N__39561\
        );

    \I__7610\ : InMux
    port map (
            O => \N__39566\,
            I => \N__39558\
        );

    \I__7609\ : InMux
    port map (
            O => \N__39565\,
            I => \N__39555\
        );

    \I__7608\ : InMux
    port map (
            O => \N__39564\,
            I => \N__39552\
        );

    \I__7607\ : Span4Mux_h
    port map (
            O => \N__39561\,
            I => \N__39547\
        );

    \I__7606\ : LocalMux
    port map (
            O => \N__39558\,
            I => \N__39547\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__39555\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_3
        );

    \I__7604\ : LocalMux
    port map (
            O => \N__39552\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_3
        );

    \I__7603\ : Odrv4
    port map (
            O => \N__39547\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_3
        );

    \I__7602\ : InMux
    port map (
            O => \N__39540\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2\
        );

    \I__7601\ : InMux
    port map (
            O => \N__39537\,
            I => \N__39532\
        );

    \I__7600\ : InMux
    port map (
            O => \N__39536\,
            I => \N__39529\
        );

    \I__7599\ : InMux
    port map (
            O => \N__39535\,
            I => \N__39526\
        );

    \I__7598\ : LocalMux
    port map (
            O => \N__39532\,
            I => \N__39521\
        );

    \I__7597\ : LocalMux
    port map (
            O => \N__39529\,
            I => \N__39521\
        );

    \I__7596\ : LocalMux
    port map (
            O => \N__39526\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_4
        );

    \I__7595\ : Odrv4
    port map (
            O => \N__39521\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_4
        );

    \I__7594\ : InMux
    port map (
            O => \N__39516\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3\
        );

    \I__7593\ : InMux
    port map (
            O => \N__39513\,
            I => \N__39509\
        );

    \I__7592\ : InMux
    port map (
            O => \N__39512\,
            I => \N__39506\
        );

    \I__7591\ : LocalMux
    port map (
            O => \N__39509\,
            I => \N__39500\
        );

    \I__7590\ : LocalMux
    port map (
            O => \N__39506\,
            I => \N__39500\
        );

    \I__7589\ : InMux
    port map (
            O => \N__39505\,
            I => \N__39497\
        );

    \I__7588\ : Span4Mux_v
    port map (
            O => \N__39500\,
            I => \N__39494\
        );

    \I__7587\ : LocalMux
    port map (
            O => \N__39497\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_5
        );

    \I__7586\ : Odrv4
    port map (
            O => \N__39494\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_5
        );

    \I__7585\ : InMux
    port map (
            O => \N__39489\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4\
        );

    \I__7584\ : CascadeMux
    port map (
            O => \N__39486\,
            I => \N__39482\
        );

    \I__7583\ : InMux
    port map (
            O => \N__39485\,
            I => \N__39479\
        );

    \I__7582\ : InMux
    port map (
            O => \N__39482\,
            I => \N__39476\
        );

    \I__7581\ : LocalMux
    port map (
            O => \N__39479\,
            I => \N__39470\
        );

    \I__7580\ : LocalMux
    port map (
            O => \N__39476\,
            I => \N__39470\
        );

    \I__7579\ : InMux
    port map (
            O => \N__39475\,
            I => \N__39467\
        );

    \I__7578\ : Span4Mux_h
    port map (
            O => \N__39470\,
            I => \N__39464\
        );

    \I__7577\ : LocalMux
    port map (
            O => \N__39467\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_6
        );

    \I__7576\ : Odrv4
    port map (
            O => \N__39464\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_6
        );

    \I__7575\ : InMux
    port map (
            O => \N__39459\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5\
        );

    \I__7574\ : InMux
    port map (
            O => \N__39456\,
            I => \N__39452\
        );

    \I__7573\ : InMux
    port map (
            O => \N__39455\,
            I => \N__39449\
        );

    \I__7572\ : LocalMux
    port map (
            O => \N__39452\,
            I => \N__39445\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__39449\,
            I => \N__39442\
        );

    \I__7570\ : InMux
    port map (
            O => \N__39448\,
            I => \N__39439\
        );

    \I__7569\ : Span4Mux_h
    port map (
            O => \N__39445\,
            I => \N__39434\
        );

    \I__7568\ : Span4Mux_h
    port map (
            O => \N__39442\,
            I => \N__39434\
        );

    \I__7567\ : LocalMux
    port map (
            O => \N__39439\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7\
        );

    \I__7566\ : Odrv4
    port map (
            O => \N__39434\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7\
        );

    \I__7565\ : InMux
    port map (
            O => \N__39429\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6\
        );

    \I__7564\ : InMux
    port map (
            O => \N__39426\,
            I => \N__39422\
        );

    \I__7563\ : InMux
    port map (
            O => \N__39425\,
            I => \N__39418\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__39422\,
            I => \N__39415\
        );

    \I__7561\ : InMux
    port map (
            O => \N__39421\,
            I => \N__39412\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__39418\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_8
        );

    \I__7559\ : Odrv4
    port map (
            O => \N__39415\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_8
        );

    \I__7558\ : LocalMux
    port map (
            O => \N__39412\,
            I => cemf_module_64ch_ctrl_inst1_paddr_fsm_8
        );

    \I__7557\ : InMux
    port map (
            O => \N__39405\,
            I => \bfn_18_21_0_\
        );

    \I__7556\ : SRMux
    port map (
            O => \N__39402\,
            I => \N__39397\
        );

    \I__7555\ : SRMux
    port map (
            O => \N__39401\,
            I => \N__39393\
        );

    \I__7554\ : SRMux
    port map (
            O => \N__39400\,
            I => \N__39389\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__39397\,
            I => \N__39386\
        );

    \I__7552\ : SRMux
    port map (
            O => \N__39396\,
            I => \N__39383\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__39393\,
            I => \N__39378\
        );

    \I__7550\ : SRMux
    port map (
            O => \N__39392\,
            I => \N__39375\
        );

    \I__7549\ : LocalMux
    port map (
            O => \N__39389\,
            I => \N__39366\
        );

    \I__7548\ : Span4Mux_s0_v
    port map (
            O => \N__39386\,
            I => \N__39366\
        );

    \I__7547\ : LocalMux
    port map (
            O => \N__39383\,
            I => \N__39366\
        );

    \I__7546\ : SRMux
    port map (
            O => \N__39382\,
            I => \N__39363\
        );

    \I__7545\ : SRMux
    port map (
            O => \N__39381\,
            I => \N__39359\
        );

    \I__7544\ : Span4Mux_v
    port map (
            O => \N__39378\,
            I => \N__39354\
        );

    \I__7543\ : LocalMux
    port map (
            O => \N__39375\,
            I => \N__39354\
        );

    \I__7542\ : SRMux
    port map (
            O => \N__39374\,
            I => \N__39351\
        );

    \I__7541\ : SRMux
    port map (
            O => \N__39373\,
            I => \N__39347\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__39366\,
            I => \N__39340\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__39363\,
            I => \N__39340\
        );

    \I__7538\ : SRMux
    port map (
            O => \N__39362\,
            I => \N__39337\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__39359\,
            I => \N__39329\
        );

    \I__7536\ : Span4Mux_h
    port map (
            O => \N__39354\,
            I => \N__39329\
        );

    \I__7535\ : LocalMux
    port map (
            O => \N__39351\,
            I => \N__39329\
        );

    \I__7534\ : SRMux
    port map (
            O => \N__39350\,
            I => \N__39326\
        );

    \I__7533\ : LocalMux
    port map (
            O => \N__39347\,
            I => \N__39322\
        );

    \I__7532\ : CascadeMux
    port map (
            O => \N__39346\,
            I => \N__39319\
        );

    \I__7531\ : CascadeMux
    port map (
            O => \N__39345\,
            I => \N__39316\
        );

    \I__7530\ : Span4Mux_v
    port map (
            O => \N__39340\,
            I => \N__39309\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__39337\,
            I => \N__39309\
        );

    \I__7528\ : SRMux
    port map (
            O => \N__39336\,
            I => \N__39306\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__39329\,
            I => \N__39300\
        );

    \I__7526\ : LocalMux
    port map (
            O => \N__39326\,
            I => \N__39300\
        );

    \I__7525\ : SRMux
    port map (
            O => \N__39325\,
            I => \N__39297\
        );

    \I__7524\ : Span4Mux_h
    port map (
            O => \N__39322\,
            I => \N__39293\
        );

    \I__7523\ : InMux
    port map (
            O => \N__39319\,
            I => \N__39290\
        );

    \I__7522\ : InMux
    port map (
            O => \N__39316\,
            I => \N__39287\
        );

    \I__7521\ : CascadeMux
    port map (
            O => \N__39315\,
            I => \N__39283\
        );

    \I__7520\ : SRMux
    port map (
            O => \N__39314\,
            I => \N__39278\
        );

    \I__7519\ : Span4Mux_h
    port map (
            O => \N__39309\,
            I => \N__39273\
        );

    \I__7518\ : LocalMux
    port map (
            O => \N__39306\,
            I => \N__39273\
        );

    \I__7517\ : SRMux
    port map (
            O => \N__39305\,
            I => \N__39270\
        );

    \I__7516\ : Span4Mux_v
    port map (
            O => \N__39300\,
            I => \N__39265\
        );

    \I__7515\ : LocalMux
    port map (
            O => \N__39297\,
            I => \N__39265\
        );

    \I__7514\ : SRMux
    port map (
            O => \N__39296\,
            I => \N__39262\
        );

    \I__7513\ : Span4Mux_v
    port map (
            O => \N__39293\,
            I => \N__39259\
        );

    \I__7512\ : LocalMux
    port map (
            O => \N__39290\,
            I => \N__39254\
        );

    \I__7511\ : LocalMux
    port map (
            O => \N__39287\,
            I => \N__39254\
        );

    \I__7510\ : InMux
    port map (
            O => \N__39286\,
            I => \N__39244\
        );

    \I__7509\ : InMux
    port map (
            O => \N__39283\,
            I => \N__39244\
        );

    \I__7508\ : InMux
    port map (
            O => \N__39282\,
            I => \N__39244\
        );

    \I__7507\ : InMux
    port map (
            O => \N__39281\,
            I => \N__39244\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__39278\,
            I => \N__39241\
        );

    \I__7505\ : Span4Mux_v
    port map (
            O => \N__39273\,
            I => \N__39236\
        );

    \I__7504\ : LocalMux
    port map (
            O => \N__39270\,
            I => \N__39236\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__39265\,
            I => \N__39231\
        );

    \I__7502\ : LocalMux
    port map (
            O => \N__39262\,
            I => \N__39231\
        );

    \I__7501\ : Span4Mux_v
    port map (
            O => \N__39259\,
            I => \N__39226\
        );

    \I__7500\ : Span4Mux_h
    port map (
            O => \N__39254\,
            I => \N__39226\
        );

    \I__7499\ : InMux
    port map (
            O => \N__39253\,
            I => \N__39223\
        );

    \I__7498\ : LocalMux
    port map (
            O => \N__39244\,
            I => \N__39220\
        );

    \I__7497\ : Span4Mux_v
    port map (
            O => \N__39241\,
            I => \N__39217\
        );

    \I__7496\ : Span4Mux_v
    port map (
            O => \N__39236\,
            I => \N__39212\
        );

    \I__7495\ : Span4Mux_v
    port map (
            O => \N__39231\,
            I => \N__39212\
        );

    \I__7494\ : Span4Mux_h
    port map (
            O => \N__39226\,
            I => \N__39207\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__39223\,
            I => \N__39207\
        );

    \I__7492\ : Span4Mux_v
    port map (
            O => \N__39220\,
            I => \N__39204\
        );

    \I__7491\ : Span4Mux_h
    port map (
            O => \N__39217\,
            I => \N__39199\
        );

    \I__7490\ : Span4Mux_h
    port map (
            O => \N__39212\,
            I => \N__39199\
        );

    \I__7489\ : Span4Mux_h
    port map (
            O => \N__39207\,
            I => \N__39196\
        );

    \I__7488\ : Sp12to4
    port map (
            O => \N__39204\,
            I => \N__39193\
        );

    \I__7487\ : Odrv4
    port map (
            O => \N__39199\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7486\ : Odrv4
    port map (
            O => \N__39196\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7485\ : Odrv12
    port map (
            O => \N__39193\,
            I => \CONSTANT_ONE_NET\
        );

    \I__7484\ : InMux
    port map (
            O => \N__39186\,
            I => \N__39183\
        );

    \I__7483\ : LocalMux
    port map (
            O => \N__39183\,
            I => \N__39180\
        );

    \I__7482\ : Span4Mux_v
    port map (
            O => \N__39180\,
            I => \N__39177\
        );

    \I__7481\ : Odrv4
    port map (
            O => \N__39177\,
            I => \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rstZ0\
        );

    \I__7480\ : SRMux
    port map (
            O => \N__39174\,
            I => \N__39171\
        );

    \I__7479\ : LocalMux
    port map (
            O => \N__39171\,
            I => \N__39168\
        );

    \I__7478\ : Span4Mux_v
    port map (
            O => \N__39168\,
            I => \N__39165\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__39165\,
            I => \N__39162\
        );

    \I__7476\ : Span4Mux_h
    port map (
            O => \N__39162\,
            I => \N__39159\
        );

    \I__7475\ : Span4Mux_v
    port map (
            O => \N__39159\,
            I => \N__39156\
        );

    \I__7474\ : Odrv4
    port map (
            O => \N__39156\,
            I => \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNOZ0\
        );

    \I__7473\ : CascadeMux
    port map (
            O => \N__39153\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa_cascade_\
        );

    \I__7472\ : CascadeMux
    port map (
            O => \N__39150\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_3_cascade_\
        );

    \I__7471\ : CascadeMux
    port map (
            O => \N__39147\,
            I => \N__39137\
        );

    \I__7470\ : InMux
    port map (
            O => \N__39146\,
            I => \N__39134\
        );

    \I__7469\ : InMux
    port map (
            O => \N__39145\,
            I => \N__39125\
        );

    \I__7468\ : InMux
    port map (
            O => \N__39144\,
            I => \N__39125\
        );

    \I__7467\ : InMux
    port map (
            O => \N__39143\,
            I => \N__39125\
        );

    \I__7466\ : InMux
    port map (
            O => \N__39142\,
            I => \N__39120\
        );

    \I__7465\ : InMux
    port map (
            O => \N__39141\,
            I => \N__39120\
        );

    \I__7464\ : InMux
    port map (
            O => \N__39140\,
            I => \N__39117\
        );

    \I__7463\ : InMux
    port map (
            O => \N__39137\,
            I => \N__39110\
        );

    \I__7462\ : LocalMux
    port map (
            O => \N__39134\,
            I => \N__39102\
        );

    \I__7461\ : InMux
    port map (
            O => \N__39133\,
            I => \N__39099\
        );

    \I__7460\ : InMux
    port map (
            O => \N__39132\,
            I => \N__39096\
        );

    \I__7459\ : LocalMux
    port map (
            O => \N__39125\,
            I => \N__39093\
        );

    \I__7458\ : LocalMux
    port map (
            O => \N__39120\,
            I => \N__39088\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__39117\,
            I => \N__39088\
        );

    \I__7456\ : InMux
    port map (
            O => \N__39116\,
            I => \N__39079\
        );

    \I__7455\ : InMux
    port map (
            O => \N__39115\,
            I => \N__39079\
        );

    \I__7454\ : InMux
    port map (
            O => \N__39114\,
            I => \N__39079\
        );

    \I__7453\ : InMux
    port map (
            O => \N__39113\,
            I => \N__39079\
        );

    \I__7452\ : LocalMux
    port map (
            O => \N__39110\,
            I => \N__39076\
        );

    \I__7451\ : InMux
    port map (
            O => \N__39109\,
            I => \N__39073\
        );

    \I__7450\ : InMux
    port map (
            O => \N__39108\,
            I => \N__39064\
        );

    \I__7449\ : InMux
    port map (
            O => \N__39107\,
            I => \N__39064\
        );

    \I__7448\ : InMux
    port map (
            O => \N__39106\,
            I => \N__39064\
        );

    \I__7447\ : InMux
    port map (
            O => \N__39105\,
            I => \N__39064\
        );

    \I__7446\ : Span4Mux_v
    port map (
            O => \N__39102\,
            I => \N__39059\
        );

    \I__7445\ : LocalMux
    port map (
            O => \N__39099\,
            I => \N__39059\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__39096\,
            I => \N_1975\
        );

    \I__7443\ : Odrv4
    port map (
            O => \N__39093\,
            I => \N_1975\
        );

    \I__7442\ : Odrv12
    port map (
            O => \N__39088\,
            I => \N_1975\
        );

    \I__7441\ : LocalMux
    port map (
            O => \N__39079\,
            I => \N_1975\
        );

    \I__7440\ : Odrv12
    port map (
            O => \N__39076\,
            I => \N_1975\
        );

    \I__7439\ : LocalMux
    port map (
            O => \N__39073\,
            I => \N_1975\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__39064\,
            I => \N_1975\
        );

    \I__7437\ : Odrv4
    port map (
            O => \N__39059\,
            I => \N_1975\
        );

    \I__7436\ : InMux
    port map (
            O => \N__39042\,
            I => \N__39039\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__39039\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNOZ0\
        );

    \I__7434\ : InMux
    port map (
            O => \N__39036\,
            I => \N__39033\
        );

    \I__7433\ : LocalMux
    port map (
            O => \N__39033\,
            I => \N__39029\
        );

    \I__7432\ : InMux
    port map (
            O => \N__39032\,
            I => \N__39026\
        );

    \I__7431\ : Span4Mux_h
    port map (
            O => \N__39029\,
            I => \N__39023\
        );

    \I__7430\ : LocalMux
    port map (
            O => \N__39026\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0\
        );

    \I__7429\ : Odrv4
    port map (
            O => \N__39023\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0\
        );

    \I__7428\ : InMux
    port map (
            O => \N__39018\,
            I => \bfn_18_20_0_\
        );

    \I__7427\ : InMux
    port map (
            O => \N__39015\,
            I => \N__39012\
        );

    \I__7426\ : LocalMux
    port map (
            O => \N__39012\,
            I => \N__39008\
        );

    \I__7425\ : CascadeMux
    port map (
            O => \N__39011\,
            I => \N__39005\
        );

    \I__7424\ : Span12Mux_v
    port map (
            O => \N__39008\,
            I => \N__39002\
        );

    \I__7423\ : InMux
    port map (
            O => \N__39005\,
            I => \N__38999\
        );

    \I__7422\ : Odrv12
    port map (
            O => \N__39002\,
            I => \cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4\
        );

    \I__7421\ : LocalMux
    port map (
            O => \N__38999\,
            I => \cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4\
        );

    \I__7420\ : InMux
    port map (
            O => \N__38994\,
            I => \N__38991\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__38991\,
            I => \N__38988\
        );

    \I__7418\ : Span4Mux_h
    port map (
            O => \N__38988\,
            I => \N__38985\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__38985\,
            I => \N__38982\
        );

    \I__7416\ : Span4Mux_h
    port map (
            O => \N__38982\,
            I => \N__38979\
        );

    \I__7415\ : Odrv4
    port map (
            O => \N__38979\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_CO\
        );

    \I__7414\ : InMux
    port map (
            O => \N__38976\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0\
        );

    \I__7413\ : InMux
    port map (
            O => \N__38973\,
            I => \N__38970\
        );

    \I__7412\ : LocalMux
    port map (
            O => \N__38970\,
            I => \N__38967\
        );

    \I__7411\ : Span4Mux_h
    port map (
            O => \N__38967\,
            I => \N__38964\
        );

    \I__7410\ : Span4Mux_h
    port map (
            O => \N__38964\,
            I => \N__38961\
        );

    \I__7409\ : Span4Mux_h
    port map (
            O => \N__38961\,
            I => \N__38957\
        );

    \I__7408\ : InMux
    port map (
            O => \N__38960\,
            I => \N__38954\
        );

    \I__7407\ : Odrv4
    port map (
            O => \N__38957\,
            I => \cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5\
        );

    \I__7406\ : LocalMux
    port map (
            O => \N__38954\,
            I => \cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5\
        );

    \I__7405\ : InMux
    port map (
            O => \N__38949\,
            I => \N__38946\
        );

    \I__7404\ : LocalMux
    port map (
            O => \N__38946\,
            I => \N__38943\
        );

    \I__7403\ : Span4Mux_h
    port map (
            O => \N__38943\,
            I => \N__38940\
        );

    \I__7402\ : Span4Mux_h
    port map (
            O => \N__38940\,
            I => \N__38937\
        );

    \I__7401\ : Span4Mux_h
    port map (
            O => \N__38937\,
            I => \N__38934\
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__38934\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_CO\
        );

    \I__7399\ : InMux
    port map (
            O => \N__38931\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1\
        );

    \I__7398\ : CascadeMux
    port map (
            O => \N__38928\,
            I => \N__38925\
        );

    \I__7397\ : InMux
    port map (
            O => \N__38925\,
            I => \N__38922\
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__38922\,
            I => \cemf_module_64ch_ctrl_inst1.c_addr_RNI3UAS1_6\
        );

    \I__7395\ : InMux
    port map (
            O => \N__38919\,
            I => \N__38916\
        );

    \I__7394\ : LocalMux
    port map (
            O => \N__38916\,
            I => \N__38913\
        );

    \I__7393\ : Span4Mux_s1_v
    port map (
            O => \N__38913\,
            I => \N__38909\
        );

    \I__7392\ : InMux
    port map (
            O => \N__38912\,
            I => \N__38906\
        );

    \I__7391\ : Span4Mux_v
    port map (
            O => \N__38909\,
            I => \N__38900\
        );

    \I__7390\ : LocalMux
    port map (
            O => \N__38906\,
            I => \N__38897\
        );

    \I__7389\ : InMux
    port map (
            O => \N__38905\,
            I => \N__38894\
        );

    \I__7388\ : InMux
    port map (
            O => \N__38904\,
            I => \N__38886\
        );

    \I__7387\ : InMux
    port map (
            O => \N__38903\,
            I => \N__38886\
        );

    \I__7386\ : Span4Mux_v
    port map (
            O => \N__38900\,
            I => \N__38881\
        );

    \I__7385\ : Span4Mux_h
    port map (
            O => \N__38897\,
            I => \N__38881\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__38894\,
            I => \N__38878\
        );

    \I__7383\ : InMux
    port map (
            O => \N__38893\,
            I => \N__38873\
        );

    \I__7382\ : InMux
    port map (
            O => \N__38892\,
            I => \N__38873\
        );

    \I__7381\ : InMux
    port map (
            O => \N__38891\,
            I => \N__38870\
        );

    \I__7380\ : LocalMux
    port map (
            O => \N__38886\,
            I => \N__38867\
        );

    \I__7379\ : Span4Mux_v
    port map (
            O => \N__38881\,
            I => \N__38862\
        );

    \I__7378\ : Span4Mux_h
    port map (
            O => \N__38878\,
            I => \N__38862\
        );

    \I__7377\ : LocalMux
    port map (
            O => \N__38873\,
            I => \N__38859\
        );

    \I__7376\ : LocalMux
    port map (
            O => \N__38870\,
            I => \N__38856\
        );

    \I__7375\ : Span4Mux_v
    port map (
            O => \N__38867\,
            I => \N__38851\
        );

    \I__7374\ : Span4Mux_h
    port map (
            O => \N__38862\,
            I => \N__38851\
        );

    \I__7373\ : Span4Mux_h
    port map (
            O => \N__38859\,
            I => \N__38848\
        );

    \I__7372\ : Span12Mux_h
    port map (
            O => \N__38856\,
            I => \N__38845\
        );

    \I__7371\ : Span4Mux_h
    port map (
            O => \N__38851\,
            I => \N__38842\
        );

    \I__7370\ : Odrv4
    port map (
            O => \N__38848\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1\
        );

    \I__7369\ : Odrv12
    port map (
            O => \N__38845\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1\
        );

    \I__7368\ : Odrv4
    port map (
            O => \N__38842\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1\
        );

    \I__7367\ : InMux
    port map (
            O => \N__38835\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2\
        );

    \I__7366\ : CascadeMux
    port map (
            O => \N__38832\,
            I => \N__38829\
        );

    \I__7365\ : InMux
    port map (
            O => \N__38829\,
            I => \N__38826\
        );

    \I__7364\ : LocalMux
    port map (
            O => \N__38826\,
            I => \cemf_module_64ch_ctrl_inst1.c_addr_RNI50BS1_7\
        );

    \I__7363\ : InMux
    port map (
            O => \N__38823\,
            I => \N__38817\
        );

    \I__7362\ : InMux
    port map (
            O => \N__38822\,
            I => \N__38814\
        );

    \I__7361\ : InMux
    port map (
            O => \N__38821\,
            I => \N__38809\
        );

    \I__7360\ : InMux
    port map (
            O => \N__38820\,
            I => \N__38809\
        );

    \I__7359\ : LocalMux
    port map (
            O => \N__38817\,
            I => \N__38803\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__38814\,
            I => \N__38799\
        );

    \I__7357\ : LocalMux
    port map (
            O => \N__38809\,
            I => \N__38796\
        );

    \I__7356\ : InMux
    port map (
            O => \N__38808\,
            I => \N__38791\
        );

    \I__7355\ : InMux
    port map (
            O => \N__38807\,
            I => \N__38791\
        );

    \I__7354\ : InMux
    port map (
            O => \N__38806\,
            I => \N__38788\
        );

    \I__7353\ : Sp12to4
    port map (
            O => \N__38803\,
            I => \N__38785\
        );

    \I__7352\ : InMux
    port map (
            O => \N__38802\,
            I => \N__38782\
        );

    \I__7351\ : Span4Mux_h
    port map (
            O => \N__38799\,
            I => \N__38779\
        );

    \I__7350\ : Span4Mux_v
    port map (
            O => \N__38796\,
            I => \N__38774\
        );

    \I__7349\ : LocalMux
    port map (
            O => \N__38791\,
            I => \N__38774\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__38788\,
            I => \N__38771\
        );

    \I__7347\ : Span12Mux_s5_v
    port map (
            O => \N__38785\,
            I => \N__38766\
        );

    \I__7346\ : LocalMux
    port map (
            O => \N__38782\,
            I => \N__38766\
        );

    \I__7345\ : Span4Mux_h
    port map (
            O => \N__38779\,
            I => \N__38763\
        );

    \I__7344\ : Span4Mux_h
    port map (
            O => \N__38774\,
            I => \N__38760\
        );

    \I__7343\ : Span12Mux_h
    port map (
            O => \N__38771\,
            I => \N__38757\
        );

    \I__7342\ : Span12Mux_v
    port map (
            O => \N__38766\,
            I => \N__38754\
        );

    \I__7341\ : Span4Mux_h
    port map (
            O => \N__38763\,
            I => \N__38751\
        );

    \I__7340\ : Odrv4
    port map (
            O => \N__38760\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1\
        );

    \I__7339\ : Odrv12
    port map (
            O => \N__38757\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1\
        );

    \I__7338\ : Odrv12
    port map (
            O => \N__38754\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1\
        );

    \I__7337\ : Odrv4
    port map (
            O => \N__38751\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1\
        );

    \I__7336\ : InMux
    port map (
            O => \N__38742\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3\
        );

    \I__7335\ : InMux
    port map (
            O => \N__38739\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4\
        );

    \I__7334\ : InMux
    port map (
            O => \N__38736\,
            I => \N__38733\
        );

    \I__7333\ : LocalMux
    port map (
            O => \N__38733\,
            I => \N__38730\
        );

    \I__7332\ : Span4Mux_h
    port map (
            O => \N__38730\,
            I => \N__38727\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__38727\,
            I => \N__38723\
        );

    \I__7330\ : InMux
    port map (
            O => \N__38726\,
            I => \N__38720\
        );

    \I__7329\ : Span4Mux_v
    port map (
            O => \N__38723\,
            I => \N__38715\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__38720\,
            I => \N__38715\
        );

    \I__7327\ : Span4Mux_h
    port map (
            O => \N__38715\,
            I => \N__38712\
        );

    \I__7326\ : Odrv4
    port map (
            O => \N__38712\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93STZ0Z1\
        );

    \I__7325\ : CascadeMux
    port map (
            O => \N__38709\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_8_0_m2_ns_1_cascade_\
        );

    \I__7324\ : InMux
    port map (
            O => \N__38706\,
            I => \N__38703\
        );

    \I__7323\ : LocalMux
    port map (
            O => \N__38703\,
            I => \N__38700\
        );

    \I__7322\ : Span4Mux_v
    port map (
            O => \N__38700\,
            I => \N__38696\
        );

    \I__7321\ : InMux
    port map (
            O => \N__38699\,
            I => \N__38693\
        );

    \I__7320\ : Span4Mux_h
    port map (
            O => \N__38696\,
            I => \N__38690\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__38693\,
            I => \N__38687\
        );

    \I__7318\ : Odrv4
    port map (
            O => \N__38690\,
            I => \N_1842_0\
        );

    \I__7317\ : Odrv12
    port map (
            O => \N__38687\,
            I => \N_1842_0\
        );

    \I__7316\ : CascadeMux
    port map (
            O => \N__38682\,
            I => \N_1842_0_cascade_\
        );

    \I__7315\ : InMux
    port map (
            O => \N__38679\,
            I => \N__38676\
        );

    \I__7314\ : LocalMux
    port map (
            O => \N__38676\,
            I => \N__38670\
        );

    \I__7313\ : InMux
    port map (
            O => \N__38675\,
            I => \N__38667\
        );

    \I__7312\ : InMux
    port map (
            O => \N__38674\,
            I => \N__38661\
        );

    \I__7311\ : InMux
    port map (
            O => \N__38673\,
            I => \N__38658\
        );

    \I__7310\ : Span12Mux_h
    port map (
            O => \N__38670\,
            I => \N__38653\
        );

    \I__7309\ : LocalMux
    port map (
            O => \N__38667\,
            I => \N__38650\
        );

    \I__7308\ : InMux
    port map (
            O => \N__38666\,
            I => \N__38643\
        );

    \I__7307\ : InMux
    port map (
            O => \N__38665\,
            I => \N__38643\
        );

    \I__7306\ : InMux
    port map (
            O => \N__38664\,
            I => \N__38643\
        );

    \I__7305\ : LocalMux
    port map (
            O => \N__38661\,
            I => \N__38638\
        );

    \I__7304\ : LocalMux
    port map (
            O => \N__38658\,
            I => \N__38638\
        );

    \I__7303\ : InMux
    port map (
            O => \N__38657\,
            I => \N__38634\
        );

    \I__7302\ : InMux
    port map (
            O => \N__38656\,
            I => \N__38631\
        );

    \I__7301\ : Span12Mux_v
    port map (
            O => \N__38653\,
            I => \N__38626\
        );

    \I__7300\ : Span12Mux_v
    port map (
            O => \N__38650\,
            I => \N__38626\
        );

    \I__7299\ : LocalMux
    port map (
            O => \N__38643\,
            I => \N__38621\
        );

    \I__7298\ : Span4Mux_v
    port map (
            O => \N__38638\,
            I => \N__38621\
        );

    \I__7297\ : InMux
    port map (
            O => \N__38637\,
            I => \N__38618\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__38634\,
            I => \N_1841_0\
        );

    \I__7295\ : LocalMux
    port map (
            O => \N__38631\,
            I => \N_1841_0\
        );

    \I__7294\ : Odrv12
    port map (
            O => \N__38626\,
            I => \N_1841_0\
        );

    \I__7293\ : Odrv4
    port map (
            O => \N__38621\,
            I => \N_1841_0\
        );

    \I__7292\ : LocalMux
    port map (
            O => \N__38618\,
            I => \N_1841_0\
        );

    \I__7291\ : InMux
    port map (
            O => \N__38607\,
            I => \N__38604\
        );

    \I__7290\ : LocalMux
    port map (
            O => \N__38604\,
            I => \N__38601\
        );

    \I__7289\ : Span4Mux_v
    port map (
            O => \N__38601\,
            I => \N__38598\
        );

    \I__7288\ : Span4Mux_h
    port map (
            O => \N__38598\,
            I => \N__38593\
        );

    \I__7287\ : InMux
    port map (
            O => \N__38597\,
            I => \N__38588\
        );

    \I__7286\ : InMux
    port map (
            O => \N__38596\,
            I => \N__38588\
        );

    \I__7285\ : Odrv4
    port map (
            O => \N__38593\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_22
        );

    \I__7284\ : LocalMux
    port map (
            O => \N__38588\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_22
        );

    \I__7283\ : InMux
    port map (
            O => \N__38583\,
            I => \N__38580\
        );

    \I__7282\ : LocalMux
    port map (
            O => \N__38580\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_22\
        );

    \I__7281\ : CascadeMux
    port map (
            O => \N__38577\,
            I => \N__38573\
        );

    \I__7280\ : InMux
    port map (
            O => \N__38576\,
            I => \N__38570\
        );

    \I__7279\ : InMux
    port map (
            O => \N__38573\,
            I => \N__38567\
        );

    \I__7278\ : LocalMux
    port map (
            O => \N__38570\,
            I => \N__38561\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__38567\,
            I => \N__38561\
        );

    \I__7276\ : InMux
    port map (
            O => \N__38566\,
            I => \N__38558\
        );

    \I__7275\ : Span4Mux_h
    port map (
            O => \N__38561\,
            I => \N__38555\
        );

    \I__7274\ : LocalMux
    port map (
            O => \N__38558\,
            I => cemf_module_64ch_ctrl_inst1_data_config_20
        );

    \I__7273\ : Odrv4
    port map (
            O => \N__38555\,
            I => cemf_module_64ch_ctrl_inst1_data_config_20
        );

    \I__7272\ : InMux
    port map (
            O => \N__38550\,
            I => \N__38547\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__38547\,
            I => \N__38544\
        );

    \I__7270\ : Span4Mux_v
    port map (
            O => \N__38544\,
            I => \N__38541\
        );

    \I__7269\ : Span4Mux_v
    port map (
            O => \N__38541\,
            I => \N__38538\
        );

    \I__7268\ : Sp12to4
    port map (
            O => \N__38538\,
            I => \N__38535\
        );

    \I__7267\ : Odrv12
    port map (
            O => \N__38535\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_30\
        );

    \I__7266\ : InMux
    port map (
            O => \N__38532\,
            I => \N__38529\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__38529\,
            I => \N__38526\
        );

    \I__7264\ : Span4Mux_h
    port map (
            O => \N__38526\,
            I => \N__38523\
        );

    \I__7263\ : Span4Mux_v
    port map (
            O => \N__38523\,
            I => \N__38520\
        );

    \I__7262\ : Span4Mux_v
    port map (
            O => \N__38520\,
            I => \N__38515\
        );

    \I__7261\ : InMux
    port map (
            O => \N__38519\,
            I => \N__38510\
        );

    \I__7260\ : InMux
    port map (
            O => \N__38518\,
            I => \N__38510\
        );

    \I__7259\ : Odrv4
    port map (
            O => \N__38515\,
            I => cemf_module_64ch_ctrl_inst1_data_config_22
        );

    \I__7258\ : LocalMux
    port map (
            O => \N__38510\,
            I => cemf_module_64ch_ctrl_inst1_data_config_22
        );

    \I__7257\ : CascadeMux
    port map (
            O => \N__38505\,
            I => \N__38502\
        );

    \I__7256\ : InMux
    port map (
            O => \N__38502\,
            I => \N__38499\
        );

    \I__7255\ : LocalMux
    port map (
            O => \N__38499\,
            I => \N__38496\
        );

    \I__7254\ : Span4Mux_h
    port map (
            O => \N__38496\,
            I => \N__38493\
        );

    \I__7253\ : Span4Mux_h
    port map (
            O => \N__38493\,
            I => \N__38490\
        );

    \I__7252\ : Odrv4
    port map (
            O => \N__38490\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_31\
        );

    \I__7251\ : InMux
    port map (
            O => \N__38487\,
            I => \N__38484\
        );

    \I__7250\ : LocalMux
    port map (
            O => \N__38484\,
            I => \N__38481\
        );

    \I__7249\ : Span4Mux_h
    port map (
            O => \N__38481\,
            I => \N__38476\
        );

    \I__7248\ : CascadeMux
    port map (
            O => \N__38480\,
            I => \N__38473\
        );

    \I__7247\ : InMux
    port map (
            O => \N__38479\,
            I => \N__38470\
        );

    \I__7246\ : Span4Mux_h
    port map (
            O => \N__38476\,
            I => \N__38467\
        );

    \I__7245\ : InMux
    port map (
            O => \N__38473\,
            I => \N__38464\
        );

    \I__7244\ : LocalMux
    port map (
            O => \N__38470\,
            I => \N__38461\
        );

    \I__7243\ : Sp12to4
    port map (
            O => \N__38467\,
            I => \N__38458\
        );

    \I__7242\ : LocalMux
    port map (
            O => \N__38464\,
            I => \N__38455\
        );

    \I__7241\ : Span4Mux_h
    port map (
            O => \N__38461\,
            I => \N__38452\
        );

    \I__7240\ : Odrv12
    port map (
            O => \N__38458\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_14
        );

    \I__7239\ : Odrv12
    port map (
            O => \N__38455\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_14
        );

    \I__7238\ : Odrv4
    port map (
            O => \N__38452\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_14
        );

    \I__7237\ : CascadeMux
    port map (
            O => \N__38445\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_22_cascade_\
        );

    \I__7236\ : InMux
    port map (
            O => \N__38442\,
            I => \N__38439\
        );

    \I__7235\ : LocalMux
    port map (
            O => \N__38439\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_22\
        );

    \I__7234\ : InMux
    port map (
            O => \N__38436\,
            I => \N__38433\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__38433\,
            I => \N__38430\
        );

    \I__7232\ : Span4Mux_v
    port map (
            O => \N__38430\,
            I => \N__38426\
        );

    \I__7231\ : CascadeMux
    port map (
            O => \N__38429\,
            I => \N__38422\
        );

    \I__7230\ : Span4Mux_h
    port map (
            O => \N__38426\,
            I => \N__38419\
        );

    \I__7229\ : InMux
    port map (
            O => \N__38425\,
            I => \N__38416\
        );

    \I__7228\ : InMux
    port map (
            O => \N__38422\,
            I => \N__38413\
        );

    \I__7227\ : Odrv4
    port map (
            O => \N__38419\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_22
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__38416\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_22
        );

    \I__7225\ : LocalMux
    port map (
            O => \N__38413\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_22
        );

    \I__7224\ : CascadeMux
    port map (
            O => \N__38406\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_22_cascade_\
        );

    \I__7223\ : InMux
    port map (
            O => \N__38403\,
            I => \N__38400\
        );

    \I__7222\ : LocalMux
    port map (
            O => \N__38400\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDDZ0Z7\
        );

    \I__7221\ : CascadeMux
    port map (
            O => \N__38397\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_21_cascade_\
        );

    \I__7220\ : InMux
    port map (
            O => \N__38394\,
            I => \N__38391\
        );

    \I__7219\ : LocalMux
    port map (
            O => \N__38391\,
            I => \N__38388\
        );

    \I__7218\ : Span12Mux_h
    port map (
            O => \N__38388\,
            I => \N__38385\
        );

    \I__7217\ : Odrv12
    port map (
            O => \N__38385\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_21
        );

    \I__7216\ : InMux
    port map (
            O => \N__38382\,
            I => \N__38379\
        );

    \I__7215\ : LocalMux
    port map (
            O => \N__38379\,
            I => \N__38376\
        );

    \I__7214\ : Span4Mux_v
    port map (
            O => \N__38376\,
            I => \N__38369\
        );

    \I__7213\ : InMux
    port map (
            O => \N__38375\,
            I => \N__38366\
        );

    \I__7212\ : InMux
    port map (
            O => \N__38374\,
            I => \N__38363\
        );

    \I__7211\ : InMux
    port map (
            O => \N__38373\,
            I => \N__38360\
        );

    \I__7210\ : InMux
    port map (
            O => \N__38372\,
            I => \N__38357\
        );

    \I__7209\ : Span4Mux_h
    port map (
            O => \N__38369\,
            I => \N__38352\
        );

    \I__7208\ : LocalMux
    port map (
            O => \N__38366\,
            I => \N__38352\
        );

    \I__7207\ : LocalMux
    port map (
            O => \N__38363\,
            I => \N__38347\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__38360\,
            I => \N__38347\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__38357\,
            I => \N__38344\
        );

    \I__7204\ : Span4Mux_h
    port map (
            O => \N__38352\,
            I => \N__38339\
        );

    \I__7203\ : Span4Mux_v
    port map (
            O => \N__38347\,
            I => \N__38339\
        );

    \I__7202\ : Span12Mux_v
    port map (
            O => \N__38344\,
            I => \N__38336\
        );

    \I__7201\ : Span4Mux_v
    port map (
            O => \N__38339\,
            I => \N__38333\
        );

    \I__7200\ : Odrv12
    port map (
            O => \N__38336\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1320\
        );

    \I__7199\ : Odrv4
    port map (
            O => \N__38333\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1320\
        );

    \I__7198\ : InMux
    port map (
            O => \N__38328\,
            I => \N__38325\
        );

    \I__7197\ : LocalMux
    port map (
            O => \N__38325\,
            I => \N__38322\
        );

    \I__7196\ : Odrv12
    port map (
            O => \N__38322\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1896\
        );

    \I__7195\ : CascadeMux
    port map (
            O => \N__38319\,
            I => \N__38312\
        );

    \I__7194\ : CascadeMux
    port map (
            O => \N__38318\,
            I => \N__38308\
        );

    \I__7193\ : CascadeMux
    port map (
            O => \N__38317\,
            I => \N__38305\
        );

    \I__7192\ : InMux
    port map (
            O => \N__38316\,
            I => \N__38298\
        );

    \I__7191\ : InMux
    port map (
            O => \N__38315\,
            I => \N__38295\
        );

    \I__7190\ : InMux
    port map (
            O => \N__38312\,
            I => \N__38292\
        );

    \I__7189\ : InMux
    port map (
            O => \N__38311\,
            I => \N__38285\
        );

    \I__7188\ : InMux
    port map (
            O => \N__38308\,
            I => \N__38285\
        );

    \I__7187\ : InMux
    port map (
            O => \N__38305\,
            I => \N__38285\
        );

    \I__7186\ : CascadeMux
    port map (
            O => \N__38304\,
            I => \N__38282\
        );

    \I__7185\ : InMux
    port map (
            O => \N__38303\,
            I => \N__38279\
        );

    \I__7184\ : InMux
    port map (
            O => \N__38302\,
            I => \N__38273\
        );

    \I__7183\ : InMux
    port map (
            O => \N__38301\,
            I => \N__38270\
        );

    \I__7182\ : LocalMux
    port map (
            O => \N__38298\,
            I => \N__38263\
        );

    \I__7181\ : LocalMux
    port map (
            O => \N__38295\,
            I => \N__38263\
        );

    \I__7180\ : LocalMux
    port map (
            O => \N__38292\,
            I => \N__38260\
        );

    \I__7179\ : LocalMux
    port map (
            O => \N__38285\,
            I => \N__38257\
        );

    \I__7178\ : InMux
    port map (
            O => \N__38282\,
            I => \N__38254\
        );

    \I__7177\ : LocalMux
    port map (
            O => \N__38279\,
            I => \N__38251\
        );

    \I__7176\ : InMux
    port map (
            O => \N__38278\,
            I => \N__38248\
        );

    \I__7175\ : InMux
    port map (
            O => \N__38277\,
            I => \N__38243\
        );

    \I__7174\ : InMux
    port map (
            O => \N__38276\,
            I => \N__38243\
        );

    \I__7173\ : LocalMux
    port map (
            O => \N__38273\,
            I => \N__38240\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__38270\,
            I => \N__38234\
        );

    \I__7171\ : InMux
    port map (
            O => \N__38269\,
            I => \N__38231\
        );

    \I__7170\ : InMux
    port map (
            O => \N__38268\,
            I => \N__38228\
        );

    \I__7169\ : Span4Mux_v
    port map (
            O => \N__38263\,
            I => \N__38223\
        );

    \I__7168\ : Span4Mux_v
    port map (
            O => \N__38260\,
            I => \N__38223\
        );

    \I__7167\ : Span4Mux_v
    port map (
            O => \N__38257\,
            I => \N__38208\
        );

    \I__7166\ : LocalMux
    port map (
            O => \N__38254\,
            I => \N__38203\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__38251\,
            I => \N__38203\
        );

    \I__7164\ : LocalMux
    port map (
            O => \N__38248\,
            I => \N__38196\
        );

    \I__7163\ : LocalMux
    port map (
            O => \N__38243\,
            I => \N__38196\
        );

    \I__7162\ : Span4Mux_v
    port map (
            O => \N__38240\,
            I => \N__38196\
        );

    \I__7161\ : InMux
    port map (
            O => \N__38239\,
            I => \N__38189\
        );

    \I__7160\ : InMux
    port map (
            O => \N__38238\,
            I => \N__38189\
        );

    \I__7159\ : InMux
    port map (
            O => \N__38237\,
            I => \N__38189\
        );

    \I__7158\ : Span4Mux_h
    port map (
            O => \N__38234\,
            I => \N__38184\
        );

    \I__7157\ : LocalMux
    port map (
            O => \N__38231\,
            I => \N__38184\
        );

    \I__7156\ : LocalMux
    port map (
            O => \N__38228\,
            I => \N__38179\
        );

    \I__7155\ : Span4Mux_h
    port map (
            O => \N__38223\,
            I => \N__38179\
        );

    \I__7154\ : InMux
    port map (
            O => \N__38222\,
            I => \N__38176\
        );

    \I__7153\ : InMux
    port map (
            O => \N__38221\,
            I => \N__38161\
        );

    \I__7152\ : InMux
    port map (
            O => \N__38220\,
            I => \N__38161\
        );

    \I__7151\ : InMux
    port map (
            O => \N__38219\,
            I => \N__38161\
        );

    \I__7150\ : InMux
    port map (
            O => \N__38218\,
            I => \N__38161\
        );

    \I__7149\ : InMux
    port map (
            O => \N__38217\,
            I => \N__38161\
        );

    \I__7148\ : InMux
    port map (
            O => \N__38216\,
            I => \N__38161\
        );

    \I__7147\ : InMux
    port map (
            O => \N__38215\,
            I => \N__38161\
        );

    \I__7146\ : InMux
    port map (
            O => \N__38214\,
            I => \N__38152\
        );

    \I__7145\ : InMux
    port map (
            O => \N__38213\,
            I => \N__38152\
        );

    \I__7144\ : InMux
    port map (
            O => \N__38212\,
            I => \N__38152\
        );

    \I__7143\ : InMux
    port map (
            O => \N__38211\,
            I => \N__38152\
        );

    \I__7142\ : Span4Mux_v
    port map (
            O => \N__38208\,
            I => \N__38147\
        );

    \I__7141\ : Span4Mux_h
    port map (
            O => \N__38203\,
            I => \N__38147\
        );

    \I__7140\ : Span4Mux_h
    port map (
            O => \N__38196\,
            I => \N__38138\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__38189\,
            I => \N__38138\
        );

    \I__7138\ : Span4Mux_v
    port map (
            O => \N__38184\,
            I => \N__38138\
        );

    \I__7137\ : Span4Mux_h
    port map (
            O => \N__38179\,
            I => \N__38138\
        );

    \I__7136\ : LocalMux
    port map (
            O => \N__38176\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\
        );

    \I__7135\ : LocalMux
    port map (
            O => \N__38161\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__38152\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\
        );

    \I__7133\ : Odrv4
    port map (
            O => \N__38147\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\
        );

    \I__7132\ : Odrv4
    port map (
            O => \N__38138\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\
        );

    \I__7131\ : CascadeMux
    port map (
            O => \N__38127\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_21_cascade_\
        );

    \I__7130\ : InMux
    port map (
            O => \N__38124\,
            I => \N__38121\
        );

    \I__7129\ : LocalMux
    port map (
            O => \N__38121\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_21\
        );

    \I__7128\ : InMux
    port map (
            O => \N__38118\,
            I => \N__38115\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__38115\,
            I => \N__38112\
        );

    \I__7126\ : Span4Mux_h
    port map (
            O => \N__38112\,
            I => \N__38109\
        );

    \I__7125\ : Odrv4
    port map (
            O => \N__38109\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_21\
        );

    \I__7124\ : CascadeMux
    port map (
            O => \N__38106\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_21_cascade_\
        );

    \I__7123\ : InMux
    port map (
            O => \N__38103\,
            I => \N__38100\
        );

    \I__7122\ : LocalMux
    port map (
            O => \N__38100\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_21\
        );

    \I__7121\ : CascadeMux
    port map (
            O => \N__38097\,
            I => \N__38094\
        );

    \I__7120\ : InMux
    port map (
            O => \N__38094\,
            I => \N__38091\
        );

    \I__7119\ : LocalMux
    port map (
            O => \N__38091\,
            I => \N__38088\
        );

    \I__7118\ : Sp12to4
    port map (
            O => \N__38088\,
            I => \N__38085\
        );

    \I__7117\ : Span12Mux_v
    port map (
            O => \N__38085\,
            I => \N__38082\
        );

    \I__7116\ : Odrv12
    port map (
            O => \N__38082\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_30\
        );

    \I__7115\ : InMux
    port map (
            O => \N__38079\,
            I => \N__38074\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__38078\,
            I => \N__38071\
        );

    \I__7113\ : CascadeMux
    port map (
            O => \N__38077\,
            I => \N__38068\
        );

    \I__7112\ : LocalMux
    port map (
            O => \N__38074\,
            I => \N__38065\
        );

    \I__7111\ : InMux
    port map (
            O => \N__38071\,
            I => \N__38062\
        );

    \I__7110\ : InMux
    port map (
            O => \N__38068\,
            I => \N__38059\
        );

    \I__7109\ : Span4Mux_v
    port map (
            O => \N__38065\,
            I => \N__38056\
        );

    \I__7108\ : LocalMux
    port map (
            O => \N__38062\,
            I => \N__38053\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__38059\,
            I => \N__38050\
        );

    \I__7106\ : Span4Mux_h
    port map (
            O => \N__38056\,
            I => \N__38047\
        );

    \I__7105\ : Span4Mux_v
    port map (
            O => \N__38053\,
            I => \N__38044\
        );

    \I__7104\ : Span12Mux_h
    port map (
            O => \N__38050\,
            I => \N__38041\
        );

    \I__7103\ : Odrv4
    port map (
            O => \N__38047\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_13
        );

    \I__7102\ : Odrv4
    port map (
            O => \N__38044\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_13
        );

    \I__7101\ : Odrv12
    port map (
            O => \N__38041\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_13
        );

    \I__7100\ : InMux
    port map (
            O => \N__38034\,
            I => \N__38031\
        );

    \I__7099\ : LocalMux
    port map (
            O => \N__38031\,
            I => \N__38028\
        );

    \I__7098\ : Odrv12
    port map (
            O => \N__38028\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_20\
        );

    \I__7097\ : InMux
    port map (
            O => \N__38025\,
            I => \N__38022\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__38022\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21\
        );

    \I__7095\ : CascadeMux
    port map (
            O => \N__38019\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21_cascade_\
        );

    \I__7094\ : CascadeMux
    port map (
            O => \N__38016\,
            I => \N__38013\
        );

    \I__7093\ : InMux
    port map (
            O => \N__38013\,
            I => \N__38010\
        );

    \I__7092\ : LocalMux
    port map (
            O => \N__38010\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_20\
        );

    \I__7091\ : InMux
    port map (
            O => \N__38007\,
            I => \N__38004\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__38004\,
            I => \N__38001\
        );

    \I__7089\ : Odrv4
    port map (
            O => \N__38001\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_20\
        );

    \I__7088\ : CascadeMux
    port map (
            O => \N__37998\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LHZ0Z5_cascade_\
        );

    \I__7087\ : InMux
    port map (
            O => \N__37995\,
            I => \N__37992\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__37992\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20\
        );

    \I__7085\ : CascadeMux
    port map (
            O => \N__37989\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20_cascade_\
        );

    \I__7084\ : InMux
    port map (
            O => \N__37986\,
            I => \N__37983\
        );

    \I__7083\ : LocalMux
    port map (
            O => \N__37983\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_20\
        );

    \I__7082\ : InMux
    port map (
            O => \N__37980\,
            I => \N__37977\
        );

    \I__7081\ : LocalMux
    port map (
            O => \N__37977\,
            I => \N__37974\
        );

    \I__7080\ : Span4Mux_h
    port map (
            O => \N__37974\,
            I => \N__37971\
        );

    \I__7079\ : Span4Mux_h
    port map (
            O => \N__37971\,
            I => \N__37968\
        );

    \I__7078\ : Span4Mux_v
    port map (
            O => \N__37968\,
            I => \N__37965\
        );

    \I__7077\ : Span4Mux_v
    port map (
            O => \N__37965\,
            I => \N__37962\
        );

    \I__7076\ : Odrv4
    port map (
            O => \N__37962\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_21
        );

    \I__7075\ : CascadeMux
    port map (
            O => \N__37959\,
            I => \N__37956\
        );

    \I__7074\ : InMux
    port map (
            O => \N__37956\,
            I => \N__37953\
        );

    \I__7073\ : LocalMux
    port map (
            O => \N__37953\,
            I => \N__37950\
        );

    \I__7072\ : Span4Mux_v
    port map (
            O => \N__37950\,
            I => \N__37947\
        );

    \I__7071\ : Span4Mux_h
    port map (
            O => \N__37947\,
            I => \N__37944\
        );

    \I__7070\ : Span4Mux_h
    port map (
            O => \N__37944\,
            I => \N__37941\
        );

    \I__7069\ : Odrv4
    port map (
            O => \N__37941\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_21
        );

    \I__7068\ : CascadeMux
    port map (
            O => \N__37938\,
            I => \N__37935\
        );

    \I__7067\ : InMux
    port map (
            O => \N__37935\,
            I => \N__37931\
        );

    \I__7066\ : CascadeMux
    port map (
            O => \N__37934\,
            I => \N__37928\
        );

    \I__7065\ : LocalMux
    port map (
            O => \N__37931\,
            I => \N__37925\
        );

    \I__7064\ : InMux
    port map (
            O => \N__37928\,
            I => \N__37922\
        );

    \I__7063\ : Span12Mux_v
    port map (
            O => \N__37925\,
            I => \N__37919\
        );

    \I__7062\ : LocalMux
    port map (
            O => \N__37922\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_23
        );

    \I__7061\ : Odrv12
    port map (
            O => \N__37919\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_23
        );

    \I__7060\ : InMux
    port map (
            O => \N__37914\,
            I => \N__37911\
        );

    \I__7059\ : LocalMux
    port map (
            O => \N__37911\,
            I => \N__37908\
        );

    \I__7058\ : Span4Mux_v
    port map (
            O => \N__37908\,
            I => \N__37905\
        );

    \I__7057\ : Sp12to4
    port map (
            O => \N__37905\,
            I => \N__37901\
        );

    \I__7056\ : InMux
    port map (
            O => \N__37904\,
            I => \N__37898\
        );

    \I__7055\ : Span12Mux_h
    port map (
            O => \N__37901\,
            I => \N__37895\
        );

    \I__7054\ : LocalMux
    port map (
            O => \N__37898\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_10
        );

    \I__7053\ : Odrv12
    port map (
            O => \N__37895\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_10
        );

    \I__7052\ : InMux
    port map (
            O => \N__37890\,
            I => \N__37887\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__37887\,
            I => \N__37884\
        );

    \I__7050\ : Odrv12
    port map (
            O => \N__37884\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_10\
        );

    \I__7049\ : InMux
    port map (
            O => \N__37881\,
            I => \N__37870\
        );

    \I__7048\ : InMux
    port map (
            O => \N__37880\,
            I => \N__37848\
        );

    \I__7047\ : InMux
    port map (
            O => \N__37879\,
            I => \N__37848\
        );

    \I__7046\ : InMux
    port map (
            O => \N__37878\,
            I => \N__37848\
        );

    \I__7045\ : InMux
    port map (
            O => \N__37877\,
            I => \N__37848\
        );

    \I__7044\ : InMux
    port map (
            O => \N__37876\,
            I => \N__37848\
        );

    \I__7043\ : InMux
    port map (
            O => \N__37875\,
            I => \N__37848\
        );

    \I__7042\ : InMux
    port map (
            O => \N__37874\,
            I => \N__37848\
        );

    \I__7041\ : InMux
    port map (
            O => \N__37873\,
            I => \N__37845\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__37870\,
            I => \N__37840\
        );

    \I__7039\ : InMux
    port map (
            O => \N__37869\,
            I => \N__37825\
        );

    \I__7038\ : InMux
    port map (
            O => \N__37868\,
            I => \N__37825\
        );

    \I__7037\ : InMux
    port map (
            O => \N__37867\,
            I => \N__37825\
        );

    \I__7036\ : InMux
    port map (
            O => \N__37866\,
            I => \N__37825\
        );

    \I__7035\ : InMux
    port map (
            O => \N__37865\,
            I => \N__37825\
        );

    \I__7034\ : InMux
    port map (
            O => \N__37864\,
            I => \N__37825\
        );

    \I__7033\ : InMux
    port map (
            O => \N__37863\,
            I => \N__37825\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__37848\,
            I => \N__37820\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__37845\,
            I => \N__37817\
        );

    \I__7030\ : InMux
    port map (
            O => \N__37844\,
            I => \N__37814\
        );

    \I__7029\ : InMux
    port map (
            O => \N__37843\,
            I => \N__37811\
        );

    \I__7028\ : Span4Mux_v
    port map (
            O => \N__37840\,
            I => \N__37798\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__37825\,
            I => \N__37798\
        );

    \I__7026\ : CascadeMux
    port map (
            O => \N__37824\,
            I => \N__37795\
        );

    \I__7025\ : CascadeMux
    port map (
            O => \N__37823\,
            I => \N__37792\
        );

    \I__7024\ : Span4Mux_h
    port map (
            O => \N__37820\,
            I => \N__37789\
        );

    \I__7023\ : Span4Mux_v
    port map (
            O => \N__37817\,
            I => \N__37784\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__37814\,
            I => \N__37784\
        );

    \I__7021\ : LocalMux
    port map (
            O => \N__37811\,
            I => \N__37781\
        );

    \I__7020\ : InMux
    port map (
            O => \N__37810\,
            I => \N__37768\
        );

    \I__7019\ : InMux
    port map (
            O => \N__37809\,
            I => \N__37768\
        );

    \I__7018\ : InMux
    port map (
            O => \N__37808\,
            I => \N__37768\
        );

    \I__7017\ : InMux
    port map (
            O => \N__37807\,
            I => \N__37768\
        );

    \I__7016\ : InMux
    port map (
            O => \N__37806\,
            I => \N__37768\
        );

    \I__7015\ : InMux
    port map (
            O => \N__37805\,
            I => \N__37768\
        );

    \I__7014\ : InMux
    port map (
            O => \N__37804\,
            I => \N__37765\
        );

    \I__7013\ : InMux
    port map (
            O => \N__37803\,
            I => \N__37762\
        );

    \I__7012\ : Span4Mux_v
    port map (
            O => \N__37798\,
            I => \N__37759\
        );

    \I__7011\ : InMux
    port map (
            O => \N__37795\,
            I => \N__37754\
        );

    \I__7010\ : InMux
    port map (
            O => \N__37792\,
            I => \N__37754\
        );

    \I__7009\ : Span4Mux_v
    port map (
            O => \N__37789\,
            I => \N__37749\
        );

    \I__7008\ : Span4Mux_h
    port map (
            O => \N__37784\,
            I => \N__37749\
        );

    \I__7007\ : Span12Mux_v
    port map (
            O => \N__37781\,
            I => \N__37742\
        );

    \I__7006\ : LocalMux
    port map (
            O => \N__37768\,
            I => \N__37742\
        );

    \I__7005\ : LocalMux
    port map (
            O => \N__37765\,
            I => \N__37742\
        );

    \I__7004\ : LocalMux
    port map (
            O => \N__37762\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable
        );

    \I__7003\ : Odrv4
    port map (
            O => \N__37759\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable
        );

    \I__7002\ : LocalMux
    port map (
            O => \N__37754\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable
        );

    \I__7001\ : Odrv4
    port map (
            O => \N__37749\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable
        );

    \I__7000\ : Odrv12
    port map (
            O => \N__37742\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable
        );

    \I__6999\ : CascadeMux
    port map (
            O => \N__37731\,
            I => \N__37728\
        );

    \I__6998\ : InMux
    port map (
            O => \N__37728\,
            I => \N__37725\
        );

    \I__6997\ : LocalMux
    port map (
            O => \N__37725\,
            I => \N__37722\
        );

    \I__6996\ : Span4Mux_v
    port map (
            O => \N__37722\,
            I => \N__37719\
        );

    \I__6995\ : Sp12to4
    port map (
            O => \N__37719\,
            I => \N__37716\
        );

    \I__6994\ : Odrv12
    port map (
            O => \N__37716\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_24
        );

    \I__6993\ : InMux
    port map (
            O => \N__37713\,
            I => \N__37710\
        );

    \I__6992\ : LocalMux
    port map (
            O => \N__37710\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_676\
        );

    \I__6991\ : InMux
    port map (
            O => \N__37707\,
            I => \N__37702\
        );

    \I__6990\ : InMux
    port map (
            O => \N__37706\,
            I => \N__37695\
        );

    \I__6989\ : InMux
    port map (
            O => \N__37705\,
            I => \N__37691\
        );

    \I__6988\ : LocalMux
    port map (
            O => \N__37702\,
            I => \N__37685\
        );

    \I__6987\ : InMux
    port map (
            O => \N__37701\,
            I => \N__37682\
        );

    \I__6986\ : InMux
    port map (
            O => \N__37700\,
            I => \N__37675\
        );

    \I__6985\ : InMux
    port map (
            O => \N__37699\,
            I => \N__37675\
        );

    \I__6984\ : InMux
    port map (
            O => \N__37698\,
            I => \N__37675\
        );

    \I__6983\ : LocalMux
    port map (
            O => \N__37695\,
            I => \N__37672\
        );

    \I__6982\ : InMux
    port map (
            O => \N__37694\,
            I => \N__37669\
        );

    \I__6981\ : LocalMux
    port map (
            O => \N__37691\,
            I => \N__37666\
        );

    \I__6980\ : InMux
    port map (
            O => \N__37690\,
            I => \N__37659\
        );

    \I__6979\ : InMux
    port map (
            O => \N__37689\,
            I => \N__37659\
        );

    \I__6978\ : InMux
    port map (
            O => \N__37688\,
            I => \N__37659\
        );

    \I__6977\ : Span4Mux_h
    port map (
            O => \N__37685\,
            I => \N__37635\
        );

    \I__6976\ : LocalMux
    port map (
            O => \N__37682\,
            I => \N__37635\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__37675\,
            I => \N__37632\
        );

    \I__6974\ : Span4Mux_h
    port map (
            O => \N__37672\,
            I => \N__37627\
        );

    \I__6973\ : LocalMux
    port map (
            O => \N__37669\,
            I => \N__37627\
        );

    \I__6972\ : Span4Mux_v
    port map (
            O => \N__37666\,
            I => \N__37622\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__37659\,
            I => \N__37622\
        );

    \I__6970\ : InMux
    port map (
            O => \N__37658\,
            I => \N__37613\
        );

    \I__6969\ : InMux
    port map (
            O => \N__37657\,
            I => \N__37613\
        );

    \I__6968\ : InMux
    port map (
            O => \N__37656\,
            I => \N__37613\
        );

    \I__6967\ : InMux
    port map (
            O => \N__37655\,
            I => \N__37613\
        );

    \I__6966\ : InMux
    port map (
            O => \N__37654\,
            I => \N__37604\
        );

    \I__6965\ : InMux
    port map (
            O => \N__37653\,
            I => \N__37604\
        );

    \I__6964\ : InMux
    port map (
            O => \N__37652\,
            I => \N__37604\
        );

    \I__6963\ : InMux
    port map (
            O => \N__37651\,
            I => \N__37604\
        );

    \I__6962\ : InMux
    port map (
            O => \N__37650\,
            I => \N__37589\
        );

    \I__6961\ : InMux
    port map (
            O => \N__37649\,
            I => \N__37589\
        );

    \I__6960\ : InMux
    port map (
            O => \N__37648\,
            I => \N__37589\
        );

    \I__6959\ : InMux
    port map (
            O => \N__37647\,
            I => \N__37589\
        );

    \I__6958\ : InMux
    port map (
            O => \N__37646\,
            I => \N__37589\
        );

    \I__6957\ : InMux
    port map (
            O => \N__37645\,
            I => \N__37589\
        );

    \I__6956\ : InMux
    port map (
            O => \N__37644\,
            I => \N__37589\
        );

    \I__6955\ : InMux
    port map (
            O => \N__37643\,
            I => \N__37580\
        );

    \I__6954\ : InMux
    port map (
            O => \N__37642\,
            I => \N__37580\
        );

    \I__6953\ : InMux
    port map (
            O => \N__37641\,
            I => \N__37580\
        );

    \I__6952\ : InMux
    port map (
            O => \N__37640\,
            I => \N__37580\
        );

    \I__6951\ : Span4Mux_v
    port map (
            O => \N__37635\,
            I => \N__37575\
        );

    \I__6950\ : Span4Mux_v
    port map (
            O => \N__37632\,
            I => \N__37575\
        );

    \I__6949\ : Span4Mux_v
    port map (
            O => \N__37627\,
            I => \N__37570\
        );

    \I__6948\ : Span4Mux_h
    port map (
            O => \N__37622\,
            I => \N__37570\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__37613\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__37604\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\
        );

    \I__6945\ : LocalMux
    port map (
            O => \N__37589\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__37580\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\
        );

    \I__6943\ : Odrv4
    port map (
            O => \N__37575\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\
        );

    \I__6942\ : Odrv4
    port map (
            O => \N__37570\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\
        );

    \I__6941\ : InMux
    port map (
            O => \N__37557\,
            I => \N__37554\
        );

    \I__6940\ : LocalMux
    port map (
            O => \N__37554\,
            I => \N__37551\
        );

    \I__6939\ : Odrv12
    port map (
            O => \N__37551\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_23\
        );

    \I__6938\ : CascadeMux
    port map (
            O => \N__37548\,
            I => \N__37545\
        );

    \I__6937\ : InMux
    port map (
            O => \N__37545\,
            I => \N__37542\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__37542\,
            I => \N__37539\
        );

    \I__6935\ : Span4Mux_v
    port map (
            O => \N__37539\,
            I => \N__37536\
        );

    \I__6934\ : Odrv4
    port map (
            O => \N__37536\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_687\
        );

    \I__6933\ : InMux
    port map (
            O => \N__37533\,
            I => \N__37530\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__37530\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_23\
        );

    \I__6931\ : CascadeMux
    port map (
            O => \N__37527\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_23_cascade_\
        );

    \I__6930\ : InMux
    port map (
            O => \N__37524\,
            I => \N__37521\
        );

    \I__6929\ : LocalMux
    port map (
            O => \N__37521\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_23\
        );

    \I__6928\ : InMux
    port map (
            O => \N__37518\,
            I => \N__37515\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__37515\,
            I => \N__37512\
        );

    \I__6926\ : Span4Mux_h
    port map (
            O => \N__37512\,
            I => \N__37509\
        );

    \I__6925\ : Span4Mux_h
    port map (
            O => \N__37509\,
            I => \N__37506\
        );

    \I__6924\ : Span4Mux_h
    port map (
            O => \N__37506\,
            I => \N__37503\
        );

    \I__6923\ : Span4Mux_v
    port map (
            O => \N__37503\,
            I => \N__37500\
        );

    \I__6922\ : Odrv4
    port map (
            O => \N__37500\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_23
        );

    \I__6921\ : CascadeMux
    port map (
            O => \N__37497\,
            I => \N__37494\
        );

    \I__6920\ : InMux
    port map (
            O => \N__37494\,
            I => \N__37491\
        );

    \I__6919\ : LocalMux
    port map (
            O => \N__37491\,
            I => \N__37488\
        );

    \I__6918\ : Span4Mux_v
    port map (
            O => \N__37488\,
            I => \N__37485\
        );

    \I__6917\ : Span4Mux_h
    port map (
            O => \N__37485\,
            I => \N__37482\
        );

    \I__6916\ : Span4Mux_h
    port map (
            O => \N__37482\,
            I => \N__37479\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__37479\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_23
        );

    \I__6914\ : CascadeMux
    port map (
            O => \N__37476\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_23_cascade_\
        );

    \I__6913\ : InMux
    port map (
            O => \N__37473\,
            I => \N__37470\
        );

    \I__6912\ : LocalMux
    port map (
            O => \N__37470\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_23\
        );

    \I__6911\ : InMux
    port map (
            O => \N__37467\,
            I => \N__37464\
        );

    \I__6910\ : LocalMux
    port map (
            O => \N__37464\,
            I => \serializer_mod_inst.shift_regZ0Z_95\
        );

    \I__6909\ : InMux
    port map (
            O => \N__37461\,
            I => \N__37458\
        );

    \I__6908\ : LocalMux
    port map (
            O => \N__37458\,
            I => \serializer_mod_inst.shift_regZ0Z_96\
        );

    \I__6907\ : InMux
    port map (
            O => \N__37455\,
            I => \N__37452\
        );

    \I__6906\ : LocalMux
    port map (
            O => \N__37452\,
            I => \serializer_mod_inst.shift_regZ0Z_97\
        );

    \I__6905\ : IoInMux
    port map (
            O => \N__37449\,
            I => \N__37446\
        );

    \I__6904\ : LocalMux
    port map (
            O => \N__37446\,
            I => \N__37443\
        );

    \I__6903\ : Span12Mux_s3_v
    port map (
            O => \N__37443\,
            I => \N__37440\
        );

    \I__6902\ : Odrv12
    port map (
            O => \N__37440\,
            I => enable_config_c
        );

    \I__6901\ : IoInMux
    port map (
            O => \N__37437\,
            I => \N__37434\
        );

    \I__6900\ : LocalMux
    port map (
            O => \N__37434\,
            I => \N__37431\
        );

    \I__6899\ : Span12Mux_s9_v
    port map (
            O => \N__37431\,
            I => \N__37428\
        );

    \I__6898\ : Span12Mux_h
    port map (
            O => \N__37428\,
            I => \N__37425\
        );

    \I__6897\ : Odrv12
    port map (
            O => \N__37425\,
            I => elec_config_out_c
        );

    \I__6896\ : InMux
    port map (
            O => \N__37422\,
            I => \N__37419\
        );

    \I__6895\ : LocalMux
    port map (
            O => \N__37419\,
            I => \N__37416\
        );

    \I__6894\ : Span4Mux_v
    port map (
            O => \N__37416\,
            I => \N__37413\
        );

    \I__6893\ : Odrv4
    port map (
            O => \N__37413\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_24\
        );

    \I__6892\ : CascadeMux
    port map (
            O => \N__37410\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_24_cascade_\
        );

    \I__6891\ : InMux
    port map (
            O => \N__37407\,
            I => \N__37404\
        );

    \I__6890\ : LocalMux
    port map (
            O => \N__37404\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_24\
        );

    \I__6889\ : InMux
    port map (
            O => \N__37401\,
            I => \N__37398\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__37398\,
            I => \N__37395\
        );

    \I__6887\ : Span4Mux_h
    port map (
            O => \N__37395\,
            I => \N__37392\
        );

    \I__6886\ : Sp12to4
    port map (
            O => \N__37392\,
            I => \N__37389\
        );

    \I__6885\ : Span12Mux_v
    port map (
            O => \N__37389\,
            I => \N__37386\
        );

    \I__6884\ : Odrv12
    port map (
            O => \N__37386\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_24
        );

    \I__6883\ : CascadeMux
    port map (
            O => \N__37383\,
            I => \N__37380\
        );

    \I__6882\ : InMux
    port map (
            O => \N__37380\,
            I => \N__37377\
        );

    \I__6881\ : LocalMux
    port map (
            O => \N__37377\,
            I => \N__37374\
        );

    \I__6880\ : Span4Mux_h
    port map (
            O => \N__37374\,
            I => \N__37371\
        );

    \I__6879\ : Span4Mux_h
    port map (
            O => \N__37371\,
            I => \N__37368\
        );

    \I__6878\ : Span4Mux_h
    port map (
            O => \N__37368\,
            I => \N__37365\
        );

    \I__6877\ : Odrv4
    port map (
            O => \N__37365\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_24
        );

    \I__6876\ : CascadeMux
    port map (
            O => \N__37362\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_24_cascade_\
        );

    \I__6875\ : InMux
    port map (
            O => \N__37359\,
            I => \N__37356\
        );

    \I__6874\ : LocalMux
    port map (
            O => \N__37356\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_24\
        );

    \I__6873\ : InMux
    port map (
            O => \N__37353\,
            I => \N__37350\
        );

    \I__6872\ : LocalMux
    port map (
            O => \N__37350\,
            I => \serializer_mod_inst.shift_regZ0Z_106\
        );

    \I__6871\ : InMux
    port map (
            O => \N__37347\,
            I => \N__37344\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__37344\,
            I => \N__37341\
        );

    \I__6869\ : Span4Mux_h
    port map (
            O => \N__37341\,
            I => \N__37338\
        );

    \I__6868\ : Odrv4
    port map (
            O => \N__37338\,
            I => \serializer_mod_inst.shift_regZ0Z_47\
        );

    \I__6867\ : InMux
    port map (
            O => \N__37335\,
            I => \N__37332\
        );

    \I__6866\ : LocalMux
    port map (
            O => \N__37332\,
            I => \serializer_mod_inst.shift_regZ0Z_94\
        );

    \I__6865\ : InMux
    port map (
            O => \N__37329\,
            I => \N__37326\
        );

    \I__6864\ : LocalMux
    port map (
            O => \N__37326\,
            I => \serializer_mod_inst.shift_regZ0Z_104\
        );

    \I__6863\ : CascadeMux
    port map (
            O => \N__37323\,
            I => \N__37320\
        );

    \I__6862\ : InMux
    port map (
            O => \N__37320\,
            I => \N__37317\
        );

    \I__6861\ : LocalMux
    port map (
            O => \N__37317\,
            I => \serializer_mod_inst.shift_regZ0Z_105\
        );

    \I__6860\ : InMux
    port map (
            O => \N__37314\,
            I => \N__37311\
        );

    \I__6859\ : LocalMux
    port map (
            O => \N__37311\,
            I => \serializer_mod_inst.shift_regZ0Z_46\
        );

    \I__6858\ : InMux
    port map (
            O => \N__37308\,
            I => \N__37305\
        );

    \I__6857\ : LocalMux
    port map (
            O => \N__37305\,
            I => \N__37302\
        );

    \I__6856\ : Odrv12
    port map (
            O => \N__37302\,
            I => \serializer_mod_inst.shift_regZ0Z_91\
        );

    \I__6855\ : InMux
    port map (
            O => \N__37299\,
            I => \N__37296\
        );

    \I__6854\ : LocalMux
    port map (
            O => \N__37296\,
            I => \serializer_mod_inst.shift_regZ0Z_92\
        );

    \I__6853\ : InMux
    port map (
            O => \N__37293\,
            I => \N__37290\
        );

    \I__6852\ : LocalMux
    port map (
            O => \N__37290\,
            I => \serializer_mod_inst.shift_regZ0Z_93\
        );

    \I__6851\ : InMux
    port map (
            O => \N__37287\,
            I => \N__37284\
        );

    \I__6850\ : LocalMux
    port map (
            O => \N__37284\,
            I => \serializer_mod_inst.shift_regZ0Z_15\
        );

    \I__6849\ : InMux
    port map (
            O => \N__37281\,
            I => \N__37278\
        );

    \I__6848\ : LocalMux
    port map (
            O => \N__37278\,
            I => \serializer_mod_inst.shift_regZ0Z_79\
        );

    \I__6847\ : InMux
    port map (
            O => \N__37275\,
            I => \N__37272\
        );

    \I__6846\ : LocalMux
    port map (
            O => \N__37272\,
            I => \serializer_mod_inst.shift_regZ0Z_16\
        );

    \I__6845\ : InMux
    port map (
            O => \N__37269\,
            I => \N__37266\
        );

    \I__6844\ : LocalMux
    port map (
            O => \N__37266\,
            I => \serializer_mod_inst.shift_regZ0Z_17\
        );

    \I__6843\ : InMux
    port map (
            O => \N__37263\,
            I => \N__37260\
        );

    \I__6842\ : LocalMux
    port map (
            O => \N__37260\,
            I => \serializer_mod_inst.shift_regZ0Z_18\
        );

    \I__6841\ : InMux
    port map (
            O => \N__37257\,
            I => \N__37254\
        );

    \I__6840\ : LocalMux
    port map (
            O => \N__37254\,
            I => \serializer_mod_inst.shift_regZ0Z_107\
        );

    \I__6839\ : InMux
    port map (
            O => \N__37251\,
            I => \N__37248\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__37248\,
            I => \serializer_mod_inst.shift_regZ0Z_69\
        );

    \I__6837\ : InMux
    port map (
            O => \N__37245\,
            I => \N__37242\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__37242\,
            I => \serializer_mod_inst.shift_regZ0Z_51\
        );

    \I__6835\ : InMux
    port map (
            O => \N__37239\,
            I => \N__37236\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__37236\,
            I => \serializer_mod_inst.shift_regZ0Z_10\
        );

    \I__6833\ : InMux
    port map (
            O => \N__37233\,
            I => \N__37230\
        );

    \I__6832\ : LocalMux
    port map (
            O => \N__37230\,
            I => \N__37227\
        );

    \I__6831\ : Span4Mux_h
    port map (
            O => \N__37227\,
            I => \N__37224\
        );

    \I__6830\ : Odrv4
    port map (
            O => \N__37224\,
            I => \serializer_mod_inst.shift_regZ0Z_55\
        );

    \I__6829\ : InMux
    port map (
            O => \N__37221\,
            I => \N__37218\
        );

    \I__6828\ : LocalMux
    port map (
            O => \N__37218\,
            I => \N__37215\
        );

    \I__6827\ : Odrv4
    port map (
            O => \N__37215\,
            I => \serializer_mod_inst.shift_regZ0Z_121\
        );

    \I__6826\ : InMux
    port map (
            O => \N__37212\,
            I => \N__37209\
        );

    \I__6825\ : LocalMux
    port map (
            O => \N__37209\,
            I => \serializer_mod_inst.shift_regZ0Z_14\
        );

    \I__6824\ : InMux
    port map (
            O => \N__37206\,
            I => \N__37203\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__37203\,
            I => \serializer_mod_inst.shift_regZ0Z_12\
        );

    \I__6822\ : InMux
    port map (
            O => \N__37200\,
            I => \N__37197\
        );

    \I__6821\ : LocalMux
    port map (
            O => \N__37197\,
            I => \serializer_mod_inst.shift_regZ0Z_13\
        );

    \I__6820\ : InMux
    port map (
            O => \N__37194\,
            I => \N__37191\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__37191\,
            I => \serializer_mod_inst.shift_regZ0Z_8\
        );

    \I__6818\ : InMux
    port map (
            O => \N__37188\,
            I => \N__37185\
        );

    \I__6817\ : LocalMux
    port map (
            O => \N__37185\,
            I => \serializer_mod_inst.shift_regZ0Z_9\
        );

    \I__6816\ : InMux
    port map (
            O => \N__37182\,
            I => \N__37179\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__37179\,
            I => \N__37176\
        );

    \I__6814\ : Odrv12
    port map (
            O => \N__37176\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8Z0Z_26\
        );

    \I__6813\ : InMux
    port map (
            O => \N__37173\,
            I => \N__37170\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__37170\,
            I => \N__37165\
        );

    \I__6811\ : InMux
    port map (
            O => \N__37169\,
            I => \N__37162\
        );

    \I__6810\ : InMux
    port map (
            O => \N__37168\,
            I => \N__37156\
        );

    \I__6809\ : Span4Mux_v
    port map (
            O => \N__37165\,
            I => \N__37153\
        );

    \I__6808\ : LocalMux
    port map (
            O => \N__37162\,
            I => \N__37150\
        );

    \I__6807\ : InMux
    port map (
            O => \N__37161\,
            I => \N__37145\
        );

    \I__6806\ : InMux
    port map (
            O => \N__37160\,
            I => \N__37140\
        );

    \I__6805\ : InMux
    port map (
            O => \N__37159\,
            I => \N__37140\
        );

    \I__6804\ : LocalMux
    port map (
            O => \N__37156\,
            I => \N__37137\
        );

    \I__6803\ : Sp12to4
    port map (
            O => \N__37153\,
            I => \N__37132\
        );

    \I__6802\ : Span12Mux_v
    port map (
            O => \N__37150\,
            I => \N__37132\
        );

    \I__6801\ : InMux
    port map (
            O => \N__37149\,
            I => \N__37127\
        );

    \I__6800\ : InMux
    port map (
            O => \N__37148\,
            I => \N__37127\
        );

    \I__6799\ : LocalMux
    port map (
            O => \N__37145\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\
        );

    \I__6798\ : LocalMux
    port map (
            O => \N__37140\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\
        );

    \I__6797\ : Odrv4
    port map (
            O => \N__37137\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\
        );

    \I__6796\ : Odrv12
    port map (
            O => \N__37132\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\
        );

    \I__6795\ : LocalMux
    port map (
            O => \N__37127\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\
        );

    \I__6794\ : InMux
    port map (
            O => \N__37116\,
            I => \N__37113\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__37113\,
            I => \N__37110\
        );

    \I__6792\ : Span4Mux_h
    port map (
            O => \N__37110\,
            I => \N__37103\
        );

    \I__6791\ : InMux
    port map (
            O => \N__37109\,
            I => \N__37100\
        );

    \I__6790\ : InMux
    port map (
            O => \N__37108\,
            I => \N__37097\
        );

    \I__6789\ : InMux
    port map (
            O => \N__37107\,
            I => \N__37092\
        );

    \I__6788\ : InMux
    port map (
            O => \N__37106\,
            I => \N__37092\
        );

    \I__6787\ : Odrv4
    port map (
            O => \N__37103\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_12\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__37100\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_12\
        );

    \I__6785\ : LocalMux
    port map (
            O => \N__37097\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_12\
        );

    \I__6784\ : LocalMux
    port map (
            O => \N__37092\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_12\
        );

    \I__6783\ : InMux
    port map (
            O => \N__37083\,
            I => \N__37077\
        );

    \I__6782\ : InMux
    port map (
            O => \N__37082\,
            I => \N__37077\
        );

    \I__6781\ : LocalMux
    port map (
            O => \N__37077\,
            I => \N__37074\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__37074\,
            I => \N__37071\
        );

    \I__6779\ : Odrv4
    port map (
            O => \N__37071\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1862\
        );

    \I__6778\ : InMux
    port map (
            O => \N__37068\,
            I => \N__37065\
        );

    \I__6777\ : LocalMux
    port map (
            O => \N__37065\,
            I => \N__37061\
        );

    \I__6776\ : InMux
    port map (
            O => \N__37064\,
            I => \N__37058\
        );

    \I__6775\ : Span4Mux_h
    port map (
            O => \N__37061\,
            I => \N__37053\
        );

    \I__6774\ : LocalMux
    port map (
            O => \N__37058\,
            I => \N__37053\
        );

    \I__6773\ : Odrv4
    port map (
            O => \N__37053\,
            I => \cemf_module_64ch_ctrl_inst1.N_1816_0\
        );

    \I__6772\ : CascadeMux
    port map (
            O => \N__37050\,
            I => \N__37045\
        );

    \I__6771\ : InMux
    port map (
            O => \N__37049\,
            I => \N__37042\
        );

    \I__6770\ : InMux
    port map (
            O => \N__37048\,
            I => \N__37037\
        );

    \I__6769\ : InMux
    port map (
            O => \N__37045\,
            I => \N__37037\
        );

    \I__6768\ : LocalMux
    port map (
            O => \N__37042\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_8\
        );

    \I__6767\ : LocalMux
    port map (
            O => \N__37037\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_8\
        );

    \I__6766\ : InMux
    port map (
            O => \N__37032\,
            I => \N__37028\
        );

    \I__6765\ : InMux
    port map (
            O => \N__37031\,
            I => \N__37025\
        );

    \I__6764\ : LocalMux
    port map (
            O => \N__37028\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__37025\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9\
        );

    \I__6762\ : InMux
    port map (
            O => \N__37020\,
            I => \N__37016\
        );

    \I__6761\ : InMux
    port map (
            O => \N__37019\,
            I => \N__37013\
        );

    \I__6760\ : LocalMux
    port map (
            O => \N__37016\,
            I => \N__37008\
        );

    \I__6759\ : LocalMux
    port map (
            O => \N__37013\,
            I => \N__37008\
        );

    \I__6758\ : Odrv12
    port map (
            O => \N__37008\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_reti_0\
        );

    \I__6757\ : InMux
    port map (
            O => \N__37005\,
            I => \N__37002\
        );

    \I__6756\ : LocalMux
    port map (
            O => \N__37002\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_6\
        );

    \I__6755\ : InMux
    port map (
            O => \N__36999\,
            I => \N__36996\
        );

    \I__6754\ : LocalMux
    port map (
            O => \N__36996\,
            I => \serializer_mod_inst.shift_regZ0Z_11\
        );

    \I__6753\ : InMux
    port map (
            O => \N__36993\,
            I => \N__36990\
        );

    \I__6752\ : LocalMux
    port map (
            O => \N__36990\,
            I => \serializer_mod_inst.shift_regZ0Z_48\
        );

    \I__6751\ : InMux
    port map (
            O => \N__36987\,
            I => \N__36984\
        );

    \I__6750\ : LocalMux
    port map (
            O => \N__36984\,
            I => \I2C_top_level_inst1.s_sda_o_qZ0Z_1\
        );

    \I__6749\ : InMux
    port map (
            O => \N__36981\,
            I => \N__36978\
        );

    \I__6748\ : LocalMux
    port map (
            O => \N__36978\,
            I => \I2C_top_level_inst1.s_sda_o_txZ0\
        );

    \I__6747\ : InMux
    port map (
            O => \N__36975\,
            I => \N__36972\
        );

    \I__6746\ : LocalMux
    port map (
            O => \N__36972\,
            I => \I2C_top_level_inst1.s_sda_o_qZ0Z_0\
        );

    \I__6745\ : InMux
    port map (
            O => \N__36969\,
            I => \N__36964\
        );

    \I__6744\ : CascadeMux
    port map (
            O => \N__36968\,
            I => \N__36961\
        );

    \I__6743\ : InMux
    port map (
            O => \N__36967\,
            I => \N__36951\
        );

    \I__6742\ : LocalMux
    port map (
            O => \N__36964\,
            I => \N__36948\
        );

    \I__6741\ : InMux
    port map (
            O => \N__36961\,
            I => \N__36939\
        );

    \I__6740\ : InMux
    port map (
            O => \N__36960\,
            I => \N__36939\
        );

    \I__6739\ : InMux
    port map (
            O => \N__36959\,
            I => \N__36939\
        );

    \I__6738\ : InMux
    port map (
            O => \N__36958\,
            I => \N__36939\
        );

    \I__6737\ : InMux
    port map (
            O => \N__36957\,
            I => \N__36934\
        );

    \I__6736\ : InMux
    port map (
            O => \N__36956\,
            I => \N__36934\
        );

    \I__6735\ : InMux
    port map (
            O => \N__36955\,
            I => \N__36929\
        );

    \I__6734\ : InMux
    port map (
            O => \N__36954\,
            I => \N__36929\
        );

    \I__6733\ : LocalMux
    port map (
            O => \N__36951\,
            I => \N__36926\
        );

    \I__6732\ : Span4Mux_v
    port map (
            O => \N__36948\,
            I => \N__36923\
        );

    \I__6731\ : LocalMux
    port map (
            O => \N__36939\,
            I => \N__36918\
        );

    \I__6730\ : LocalMux
    port map (
            O => \N__36934\,
            I => \N__36918\
        );

    \I__6729\ : LocalMux
    port map (
            O => \N__36929\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_a\
        );

    \I__6728\ : Odrv12
    port map (
            O => \N__36926\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_a\
        );

    \I__6727\ : Odrv4
    port map (
            O => \N__36923\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_a\
        );

    \I__6726\ : Odrv4
    port map (
            O => \N__36918\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_a\
        );

    \I__6725\ : CascadeMux
    port map (
            O => \N__36909\,
            I => \N__36905\
        );

    \I__6724\ : InMux
    port map (
            O => \N__36908\,
            I => \N__36901\
        );

    \I__6723\ : InMux
    port map (
            O => \N__36905\,
            I => \N__36897\
        );

    \I__6722\ : InMux
    port map (
            O => \N__36904\,
            I => \N__36894\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__36901\,
            I => \N__36891\
        );

    \I__6720\ : InMux
    port map (
            O => \N__36900\,
            I => \N__36888\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__36897\,
            I => \N__36883\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__36894\,
            I => \N__36883\
        );

    \I__6717\ : Span4Mux_h
    port map (
            O => \N__36891\,
            I => \N__36880\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__36888\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0\
        );

    \I__6715\ : Odrv4
    port map (
            O => \N__36883\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0\
        );

    \I__6714\ : Odrv4
    port map (
            O => \N__36880\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0\
        );

    \I__6713\ : InMux
    port map (
            O => \N__36873\,
            I => \N__36870\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__36870\,
            I => \N__36865\
        );

    \I__6711\ : InMux
    port map (
            O => \N__36869\,
            I => \N__36862\
        );

    \I__6710\ : InMux
    port map (
            O => \N__36868\,
            I => \N__36859\
        );

    \I__6709\ : Span4Mux_h
    port map (
            O => \N__36865\,
            I => \N__36856\
        );

    \I__6708\ : LocalMux
    port map (
            O => \N__36862\,
            I => \N__36851\
        );

    \I__6707\ : LocalMux
    port map (
            O => \N__36859\,
            I => \N__36851\
        );

    \I__6706\ : Odrv4
    port map (
            O => \N__36856\,
            I => \cemf_module_64ch_ctrl_inst1.N_1855_0\
        );

    \I__6705\ : Odrv12
    port map (
            O => \N__36851\,
            I => \cemf_module_64ch_ctrl_inst1.N_1855_0\
        );

    \I__6704\ : CascadeMux
    port map (
            O => \N__36846\,
            I => \cemf_module_64ch_ctrl_inst1.N_1855_0_cascade_\
        );

    \I__6703\ : CascadeMux
    port map (
            O => \N__36843\,
            I => \N__36840\
        );

    \I__6702\ : InMux
    port map (
            O => \N__36840\,
            I => \N__36831\
        );

    \I__6701\ : InMux
    port map (
            O => \N__36839\,
            I => \N__36831\
        );

    \I__6700\ : InMux
    port map (
            O => \N__36838\,
            I => \N__36828\
        );

    \I__6699\ : InMux
    port map (
            O => \N__36837\,
            I => \N__36825\
        );

    \I__6698\ : InMux
    port map (
            O => \N__36836\,
            I => \N__36822\
        );

    \I__6697\ : LocalMux
    port map (
            O => \N__36831\,
            I => \N__36819\
        );

    \I__6696\ : LocalMux
    port map (
            O => \N__36828\,
            I => \N__36816\
        );

    \I__6695\ : LocalMux
    port map (
            O => \N__36825\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0\
        );

    \I__6694\ : LocalMux
    port map (
            O => \N__36822\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0\
        );

    \I__6693\ : Odrv4
    port map (
            O => \N__36819\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0\
        );

    \I__6692\ : Odrv4
    port map (
            O => \N__36816\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0\
        );

    \I__6691\ : InMux
    port map (
            O => \N__36807\,
            I => \N__36804\
        );

    \I__6690\ : LocalMux
    port map (
            O => \N__36804\,
            I => \N__36801\
        );

    \I__6689\ : Span4Mux_h
    port map (
            O => \N__36801\,
            I => \N__36798\
        );

    \I__6688\ : Span4Mux_v
    port map (
            O => \N__36798\,
            I => \N__36795\
        );

    \I__6687\ : Odrv4
    port map (
            O => \N__36795\,
            I => \cemf_module_64ch_ctrl_inst1.N_1857_0\
        );

    \I__6686\ : CascadeMux
    port map (
            O => \N__36792\,
            I => \cemf_module_64ch_ctrl_inst1.N_1857_0_cascade_\
        );

    \I__6685\ : CascadeMux
    port map (
            O => \N__36789\,
            I => \N__36786\
        );

    \I__6684\ : InMux
    port map (
            O => \N__36786\,
            I => \N__36780\
        );

    \I__6683\ : InMux
    port map (
            O => \N__36785\,
            I => \N__36780\
        );

    \I__6682\ : LocalMux
    port map (
            O => \N__36780\,
            I => \N__36777\
        );

    \I__6681\ : Span4Mux_v
    port map (
            O => \N__36777\,
            I => \N__36774\
        );

    \I__6680\ : Odrv4
    port map (
            O => \N__36774\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_384\
        );

    \I__6679\ : InMux
    port map (
            O => \N__36771\,
            I => \N__36767\
        );

    \I__6678\ : InMux
    port map (
            O => \N__36770\,
            I => \N__36764\
        );

    \I__6677\ : LocalMux
    port map (
            O => \N__36767\,
            I => \N__36759\
        );

    \I__6676\ : LocalMux
    port map (
            O => \N__36764\,
            I => \N__36759\
        );

    \I__6675\ : Span12Mux_v
    port map (
            O => \N__36759\,
            I => \N__36756\
        );

    \I__6674\ : Odrv12
    port map (
            O => \N__36756\,
            I => \cemf_module_64ch_ctrl_inst1.N_1854_0\
        );

    \I__6673\ : InMux
    port map (
            O => \N__36753\,
            I => \N__36750\
        );

    \I__6672\ : LocalMux
    port map (
            O => \N__36750\,
            I => \N__36747\
        );

    \I__6671\ : Span4Mux_h
    port map (
            O => \N__36747\,
            I => \N__36744\
        );

    \I__6670\ : Span4Mux_v
    port map (
            O => \N__36744\,
            I => \N__36741\
        );

    \I__6669\ : Odrv4
    port map (
            O => \N__36741\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1840_0\
        );

    \I__6668\ : InMux
    port map (
            O => \N__36738\,
            I => \N__36731\
        );

    \I__6667\ : InMux
    port map (
            O => \N__36737\,
            I => \N__36722\
        );

    \I__6666\ : InMux
    port map (
            O => \N__36736\,
            I => \N__36722\
        );

    \I__6665\ : InMux
    port map (
            O => \N__36735\,
            I => \N__36722\
        );

    \I__6664\ : InMux
    port map (
            O => \N__36734\,
            I => \N__36722\
        );

    \I__6663\ : LocalMux
    port map (
            O => \N__36731\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i\
        );

    \I__6662\ : LocalMux
    port map (
            O => \N__36722\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i\
        );

    \I__6661\ : InMux
    port map (
            O => \N__36717\,
            I => \N__36711\
        );

    \I__6660\ : InMux
    port map (
            O => \N__36716\,
            I => \N__36708\
        );

    \I__6659\ : InMux
    port map (
            O => \N__36715\,
            I => \N__36703\
        );

    \I__6658\ : InMux
    port map (
            O => \N__36714\,
            I => \N__36703\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__36711\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0\
        );

    \I__6656\ : LocalMux
    port map (
            O => \N__36708\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__36703\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0\
        );

    \I__6654\ : InMux
    port map (
            O => \N__36696\,
            I => \N__36690\
        );

    \I__6653\ : InMux
    port map (
            O => \N__36695\,
            I => \N__36690\
        );

    \I__6652\ : LocalMux
    port map (
            O => \N__36690\,
            I => \N__36686\
        );

    \I__6651\ : InMux
    port map (
            O => \N__36689\,
            I => \N__36683\
        );

    \I__6650\ : Odrv4
    port map (
            O => \N__36686\,
            I => \cemf_module_64ch_ctrl_inst1.N_383\
        );

    \I__6649\ : LocalMux
    port map (
            O => \N__36683\,
            I => \cemf_module_64ch_ctrl_inst1.N_383\
        );

    \I__6648\ : InMux
    port map (
            O => \N__36678\,
            I => \N__36672\
        );

    \I__6647\ : InMux
    port map (
            O => \N__36677\,
            I => \N__36665\
        );

    \I__6646\ : InMux
    port map (
            O => \N__36676\,
            I => \N__36665\
        );

    \I__6645\ : InMux
    port map (
            O => \N__36675\,
            I => \N__36665\
        );

    \I__6644\ : LocalMux
    port map (
            O => \N__36672\,
            I => \N__36662\
        );

    \I__6643\ : LocalMux
    port map (
            O => \N__36665\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0\
        );

    \I__6642\ : Odrv4
    port map (
            O => \N__36662\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0\
        );

    \I__6641\ : InMux
    port map (
            O => \N__36657\,
            I => \N__36654\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__36654\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_6\
        );

    \I__6639\ : InMux
    port map (
            O => \N__36651\,
            I => \N__36648\
        );

    \I__6638\ : LocalMux
    port map (
            O => \N__36648\,
            I => \N__36644\
        );

    \I__6637\ : CascadeMux
    port map (
            O => \N__36647\,
            I => \N__36635\
        );

    \I__6636\ : Span4Mux_h
    port map (
            O => \N__36644\,
            I => \N__36631\
        );

    \I__6635\ : InMux
    port map (
            O => \N__36643\,
            I => \N__36626\
        );

    \I__6634\ : InMux
    port map (
            O => \N__36642\,
            I => \N__36626\
        );

    \I__6633\ : InMux
    port map (
            O => \N__36641\,
            I => \N__36623\
        );

    \I__6632\ : InMux
    port map (
            O => \N__36640\,
            I => \N__36616\
        );

    \I__6631\ : InMux
    port map (
            O => \N__36639\,
            I => \N__36616\
        );

    \I__6630\ : InMux
    port map (
            O => \N__36638\,
            I => \N__36616\
        );

    \I__6629\ : InMux
    port map (
            O => \N__36635\,
            I => \N__36611\
        );

    \I__6628\ : InMux
    port map (
            O => \N__36634\,
            I => \N__36611\
        );

    \I__6627\ : Odrv4
    port map (
            O => \N__36631\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\
        );

    \I__6626\ : LocalMux
    port map (
            O => \N__36626\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\
        );

    \I__6625\ : LocalMux
    port map (
            O => \N__36623\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\
        );

    \I__6624\ : LocalMux
    port map (
            O => \N__36616\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\
        );

    \I__6623\ : LocalMux
    port map (
            O => \N__36611\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\
        );

    \I__6622\ : InMux
    port map (
            O => \N__36600\,
            I => \N__36596\
        );

    \I__6621\ : InMux
    port map (
            O => \N__36599\,
            I => \N__36592\
        );

    \I__6620\ : LocalMux
    port map (
            O => \N__36596\,
            I => \N__36589\
        );

    \I__6619\ : InMux
    port map (
            O => \N__36595\,
            I => \N__36586\
        );

    \I__6618\ : LocalMux
    port map (
            O => \N__36592\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4\
        );

    \I__6617\ : Odrv4
    port map (
            O => \N__36589\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__36586\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4\
        );

    \I__6615\ : InMux
    port map (
            O => \N__36579\,
            I => \N__36576\
        );

    \I__6614\ : LocalMux
    port map (
            O => \N__36576\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_3_1\
        );

    \I__6613\ : InMux
    port map (
            O => \N__36573\,
            I => \N__36570\
        );

    \I__6612\ : LocalMux
    port map (
            O => \N__36570\,
            I => \N__36567\
        );

    \I__6611\ : Span4Mux_v
    port map (
            O => \N__36567\,
            I => \N__36564\
        );

    \I__6610\ : Odrv4
    port map (
            O => \N__36564\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_5_1\
        );

    \I__6609\ : InMux
    port map (
            O => \N__36561\,
            I => \N__36558\
        );

    \I__6608\ : LocalMux
    port map (
            O => \N__36558\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_2_1\
        );

    \I__6607\ : CascadeMux
    port map (
            O => \N__36555\,
            I => \I2C_top_level_inst1.N_4_0_cascade_\
        );

    \I__6606\ : InMux
    port map (
            O => \N__36552\,
            I => \N__36549\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__36549\,
            I => \N__36546\
        );

    \I__6604\ : Span12Mux_h
    port map (
            O => \N__36546\,
            I => \N__36543\
        );

    \I__6603\ : Odrv12
    port map (
            O => \N__36543\,
            I => \I2C_top_level_inst1.N_259\
        );

    \I__6602\ : InMux
    port map (
            O => \N__36540\,
            I => \N__36537\
        );

    \I__6601\ : LocalMux
    port map (
            O => \N__36537\,
            I => \N__36534\
        );

    \I__6600\ : Span4Mux_h
    port map (
            O => \N__36534\,
            I => \N__36531\
        );

    \I__6599\ : Span4Mux_v
    port map (
            O => \N__36531\,
            I => \N__36527\
        );

    \I__6598\ : InMux
    port map (
            O => \N__36530\,
            I => \N__36524\
        );

    \I__6597\ : Odrv4
    port map (
            O => \N__36527\,
            I => \cemf_module_64ch_ctrl_inst1.N_1848_0\
        );

    \I__6596\ : LocalMux
    port map (
            O => \N__36524\,
            I => \cemf_module_64ch_ctrl_inst1.N_1848_0\
        );

    \I__6595\ : InMux
    port map (
            O => \N__36519\,
            I => \N__36516\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__36516\,
            I => \N__36513\
        );

    \I__6593\ : Odrv4
    port map (
            O => \N__36513\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7Z0Z_26\
        );

    \I__6592\ : CEMux
    port map (
            O => \N__36510\,
            I => \N__36507\
        );

    \I__6591\ : LocalMux
    port map (
            O => \N__36507\,
            I => \N__36504\
        );

    \I__6590\ : Span4Mux_v
    port map (
            O => \N__36504\,
            I => \N__36500\
        );

    \I__6589\ : CEMux
    port map (
            O => \N__36503\,
            I => \N__36497\
        );

    \I__6588\ : Span4Mux_h
    port map (
            O => \N__36500\,
            I => \N__36494\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__36497\,
            I => \N__36491\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__36494\,
            I => \I2C_top_level_inst1.N_327_i\
        );

    \I__6585\ : Odrv12
    port map (
            O => \N__36491\,
            I => \I2C_top_level_inst1.N_327_i\
        );

    \I__6584\ : InMux
    port map (
            O => \N__36486\,
            I => \N__36483\
        );

    \I__6583\ : LocalMux
    port map (
            O => \N__36483\,
            I => \N__36480\
        );

    \I__6582\ : Odrv4
    port map (
            O => \N__36480\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0\
        );

    \I__6581\ : InMux
    port map (
            O => \N__36477\,
            I => \N__36474\
        );

    \I__6580\ : LocalMux
    port map (
            O => \N__36474\,
            I => \N__36469\
        );

    \I__6579\ : InMux
    port map (
            O => \N__36473\,
            I => \N__36466\
        );

    \I__6578\ : InMux
    port map (
            O => \N__36472\,
            I => \N__36463\
        );

    \I__6577\ : Span4Mux_v
    port map (
            O => \N__36469\,
            I => \N__36460\
        );

    \I__6576\ : LocalMux
    port map (
            O => \N__36466\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0\
        );

    \I__6575\ : LocalMux
    port map (
            O => \N__36463\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0\
        );

    \I__6574\ : Odrv4
    port map (
            O => \N__36460\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0\
        );

    \I__6573\ : CascadeMux
    port map (
            O => \N__36453\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0_cascade_\
        );

    \I__6572\ : InMux
    port map (
            O => \N__36450\,
            I => \N__36444\
        );

    \I__6571\ : InMux
    port map (
            O => \N__36449\,
            I => \N__36444\
        );

    \I__6570\ : LocalMux
    port map (
            O => \N__36444\,
            I => \N__36441\
        );

    \I__6569\ : Span4Mux_h
    port map (
            O => \N__36441\,
            I => \N__36438\
        );

    \I__6568\ : Odrv4
    port map (
            O => \N__36438\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_113_0\
        );

    \I__6567\ : InMux
    port map (
            O => \N__36435\,
            I => \N__36432\
        );

    \I__6566\ : LocalMux
    port map (
            O => \N__36432\,
            I => \N__36428\
        );

    \I__6565\ : InMux
    port map (
            O => \N__36431\,
            I => \N__36425\
        );

    \I__6564\ : Span4Mux_h
    port map (
            O => \N__36428\,
            I => \N__36422\
        );

    \I__6563\ : LocalMux
    port map (
            O => \N__36425\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1\
        );

    \I__6562\ : Odrv4
    port map (
            O => \N__36422\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1\
        );

    \I__6561\ : CascadeMux
    port map (
            O => \N__36417\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0_cascade_\
        );

    \I__6560\ : InMux
    port map (
            O => \N__36414\,
            I => \N__36411\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__36411\,
            I => \I2C_top_level_inst1.s_command_4\
        );

    \I__6558\ : InMux
    port map (
            O => \N__36408\,
            I => \N__36405\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__36405\,
            I => \I2C_top_level_inst1.s_command_5\
        );

    \I__6556\ : InMux
    port map (
            O => \N__36402\,
            I => \N__36399\
        );

    \I__6555\ : LocalMux
    port map (
            O => \N__36399\,
            I => \I2C_top_level_inst1.s_command_6\
        );

    \I__6554\ : InMux
    port map (
            O => \N__36396\,
            I => \N__36393\
        );

    \I__6553\ : LocalMux
    port map (
            O => \N__36393\,
            I => \N__36390\
        );

    \I__6552\ : Odrv4
    port map (
            O => \N__36390\,
            I => \N_1803\
        );

    \I__6551\ : CascadeMux
    port map (
            O => \N__36387\,
            I => \N_1803_cascade_\
        );

    \I__6550\ : CascadeMux
    port map (
            O => \N__36384\,
            I => \N__36381\
        );

    \I__6549\ : InMux
    port map (
            O => \N__36381\,
            I => \N__36378\
        );

    \I__6548\ : LocalMux
    port map (
            O => \N__36378\,
            I => \I2C_top_level_inst1.s_command_7\
        );

    \I__6547\ : InMux
    port map (
            O => \N__36375\,
            I => \N__36372\
        );

    \I__6546\ : LocalMux
    port map (
            O => \N__36372\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6Z0Z_26\
        );

    \I__6545\ : CascadeMux
    port map (
            O => \N__36369\,
            I => \N_1613_cascade_\
        );

    \I__6544\ : InMux
    port map (
            O => \N__36366\,
            I => \N__36363\
        );

    \I__6543\ : LocalMux
    port map (
            O => \N__36363\,
            I => \N__36359\
        );

    \I__6542\ : InMux
    port map (
            O => \N__36362\,
            I => \N__36356\
        );

    \I__6541\ : Sp12to4
    port map (
            O => \N__36359\,
            I => \N__36351\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__36356\,
            I => \N__36348\
        );

    \I__6539\ : InMux
    port map (
            O => \N__36355\,
            I => \N__36345\
        );

    \I__6538\ : InMux
    port map (
            O => \N__36354\,
            I => \N__36342\
        );

    \I__6537\ : Span12Mux_s7_v
    port map (
            O => \N__36351\,
            I => \N__36339\
        );

    \I__6536\ : Span4Mux_v
    port map (
            O => \N__36348\,
            I => \N__36336\
        );

    \I__6535\ : LocalMux
    port map (
            O => \N__36345\,
            I => \N__36333\
        );

    \I__6534\ : LocalMux
    port map (
            O => \N__36342\,
            I => \N_1860_0\
        );

    \I__6533\ : Odrv12
    port map (
            O => \N__36339\,
            I => \N_1860_0\
        );

    \I__6532\ : Odrv4
    port map (
            O => \N__36336\,
            I => \N_1860_0\
        );

    \I__6531\ : Odrv12
    port map (
            O => \N__36333\,
            I => \N_1860_0\
        );

    \I__6530\ : InMux
    port map (
            O => \N__36324\,
            I => \N__36321\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__36321\,
            I => \N__36318\
        );

    \I__6528\ : Span4Mux_h
    port map (
            O => \N__36318\,
            I => \N__36314\
        );

    \I__6527\ : InMux
    port map (
            O => \N__36317\,
            I => \N__36311\
        );

    \I__6526\ : Odrv4
    port map (
            O => \N__36314\,
            I => \N_202_0\
        );

    \I__6525\ : LocalMux
    port map (
            O => \N__36311\,
            I => \N_202_0\
        );

    \I__6524\ : InMux
    port map (
            O => \N__36306\,
            I => \N__36302\
        );

    \I__6523\ : InMux
    port map (
            O => \N__36305\,
            I => \N__36299\
        );

    \I__6522\ : LocalMux
    port map (
            O => \N__36302\,
            I => \N__36296\
        );

    \I__6521\ : LocalMux
    port map (
            O => \N__36299\,
            I => \N__36291\
        );

    \I__6520\ : Span4Mux_h
    port map (
            O => \N__36296\,
            I => \N__36288\
        );

    \I__6519\ : InMux
    port map (
            O => \N__36295\,
            I => \N__36283\
        );

    \I__6518\ : InMux
    port map (
            O => \N__36294\,
            I => \N__36283\
        );

    \I__6517\ : Span4Mux_v
    port map (
            O => \N__36291\,
            I => \N__36280\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__36288\,
            I => \N_1859_0\
        );

    \I__6515\ : LocalMux
    port map (
            O => \N__36283\,
            I => \N_1859_0\
        );

    \I__6514\ : Odrv4
    port map (
            O => \N__36280\,
            I => \N_1859_0\
        );

    \I__6513\ : CascadeMux
    port map (
            O => \N__36273\,
            I => \N__36269\
        );

    \I__6512\ : InMux
    port map (
            O => \N__36272\,
            I => \N__36265\
        );

    \I__6511\ : InMux
    port map (
            O => \N__36269\,
            I => \N__36260\
        );

    \I__6510\ : InMux
    port map (
            O => \N__36268\,
            I => \N__36260\
        );

    \I__6509\ : LocalMux
    port map (
            O => \N__36265\,
            I => \N__36256\
        );

    \I__6508\ : LocalMux
    port map (
            O => \N__36260\,
            I => \N__36253\
        );

    \I__6507\ : InMux
    port map (
            O => \N__36259\,
            I => \N__36250\
        );

    \I__6506\ : Span4Mux_h
    port map (
            O => \N__36256\,
            I => \N__36247\
        );

    \I__6505\ : Span4Mux_v
    port map (
            O => \N__36253\,
            I => \N__36244\
        );

    \I__6504\ : LocalMux
    port map (
            O => \N__36250\,
            I => \N_1861_0\
        );

    \I__6503\ : Odrv4
    port map (
            O => \N__36247\,
            I => \N_1861_0\
        );

    \I__6502\ : Odrv4
    port map (
            O => \N__36244\,
            I => \N_1861_0\
        );

    \I__6501\ : InMux
    port map (
            O => \N__36237\,
            I => \N__36228\
        );

    \I__6500\ : InMux
    port map (
            O => \N__36236\,
            I => \N__36228\
        );

    \I__6499\ : InMux
    port map (
            O => \N__36235\,
            I => \N__36228\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__36228\,
            I => \N__36225\
        );

    \I__6497\ : Span4Mux_h
    port map (
            O => \N__36225\,
            I => \N__36222\
        );

    \I__6496\ : Span4Mux_h
    port map (
            O => \N__36222\,
            I => \N__36215\
        );

    \I__6495\ : InMux
    port map (
            O => \N__36221\,
            I => \N__36206\
        );

    \I__6494\ : InMux
    port map (
            O => \N__36220\,
            I => \N__36206\
        );

    \I__6493\ : InMux
    port map (
            O => \N__36219\,
            I => \N__36206\
        );

    \I__6492\ : InMux
    port map (
            O => \N__36218\,
            I => \N__36206\
        );

    \I__6491\ : Odrv4
    port map (
            O => \N__36215\,
            I => \N_1613\
        );

    \I__6490\ : LocalMux
    port map (
            O => \N__36206\,
            I => \N_1613\
        );

    \I__6489\ : InMux
    port map (
            O => \N__36201\,
            I => \N__36198\
        );

    \I__6488\ : LocalMux
    port map (
            O => \N__36198\,
            I => \N__36195\
        );

    \I__6487\ : Odrv12
    port map (
            O => \N__36195\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_604\
        );

    \I__6486\ : CascadeMux
    port map (
            O => \N__36192\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20_cascade_\
        );

    \I__6485\ : InMux
    port map (
            O => \N__36189\,
            I => \N__36186\
        );

    \I__6484\ : LocalMux
    port map (
            O => \N__36186\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_20\
        );

    \I__6483\ : InMux
    port map (
            O => \N__36183\,
            I => \N__36179\
        );

    \I__6482\ : InMux
    port map (
            O => \N__36182\,
            I => \N__36176\
        );

    \I__6481\ : LocalMux
    port map (
            O => \N__36179\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21\
        );

    \I__6480\ : LocalMux
    port map (
            O => \N__36176\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21\
        );

    \I__6479\ : InMux
    port map (
            O => \N__36171\,
            I => \N__36168\
        );

    \I__6478\ : LocalMux
    port map (
            O => \N__36168\,
            I => \N__36165\
        );

    \I__6477\ : Sp12to4
    port map (
            O => \N__36165\,
            I => \N__36162\
        );

    \I__6476\ : Odrv12
    port map (
            O => \N__36162\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_21\
        );

    \I__6475\ : InMux
    port map (
            O => \N__36159\,
            I => \N__36155\
        );

    \I__6474\ : InMux
    port map (
            O => \N__36158\,
            I => \N__36152\
        );

    \I__6473\ : LocalMux
    port map (
            O => \N__36155\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22\
        );

    \I__6472\ : LocalMux
    port map (
            O => \N__36152\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22\
        );

    \I__6471\ : InMux
    port map (
            O => \N__36147\,
            I => \N__36144\
        );

    \I__6470\ : LocalMux
    port map (
            O => \N__36144\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_22\
        );

    \I__6469\ : InMux
    port map (
            O => \N__36141\,
            I => \N__36137\
        );

    \I__6468\ : InMux
    port map (
            O => \N__36140\,
            I => \N__36134\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__36137\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__36134\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23\
        );

    \I__6465\ : InMux
    port map (
            O => \N__36129\,
            I => \N__36126\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__36126\,
            I => \N__36123\
        );

    \I__6463\ : Span4Mux_v
    port map (
            O => \N__36123\,
            I => \N__36120\
        );

    \I__6462\ : Sp12to4
    port map (
            O => \N__36120\,
            I => \N__36117\
        );

    \I__6461\ : Odrv12
    port map (
            O => \N__36117\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_conf\
        );

    \I__6460\ : CascadeMux
    port map (
            O => \N__36114\,
            I => \N__36110\
        );

    \I__6459\ : CascadeMux
    port map (
            O => \N__36113\,
            I => \N__36107\
        );

    \I__6458\ : CascadeBuf
    port map (
            O => \N__36110\,
            I => \N__36104\
        );

    \I__6457\ : CascadeBuf
    port map (
            O => \N__36107\,
            I => \N__36101\
        );

    \I__6456\ : CascadeMux
    port map (
            O => \N__36104\,
            I => \N__36098\
        );

    \I__6455\ : CascadeMux
    port map (
            O => \N__36101\,
            I => \N__36095\
        );

    \I__6454\ : CascadeBuf
    port map (
            O => \N__36098\,
            I => \N__36092\
        );

    \I__6453\ : CascadeBuf
    port map (
            O => \N__36095\,
            I => \N__36089\
        );

    \I__6452\ : CascadeMux
    port map (
            O => \N__36092\,
            I => \N__36086\
        );

    \I__6451\ : CascadeMux
    port map (
            O => \N__36089\,
            I => \N__36083\
        );

    \I__6450\ : CascadeBuf
    port map (
            O => \N__36086\,
            I => \N__36080\
        );

    \I__6449\ : CascadeBuf
    port map (
            O => \N__36083\,
            I => \N__36077\
        );

    \I__6448\ : CascadeMux
    port map (
            O => \N__36080\,
            I => \N__36074\
        );

    \I__6447\ : CascadeMux
    port map (
            O => \N__36077\,
            I => \N__36071\
        );

    \I__6446\ : CascadeBuf
    port map (
            O => \N__36074\,
            I => \N__36068\
        );

    \I__6445\ : CascadeBuf
    port map (
            O => \N__36071\,
            I => \N__36065\
        );

    \I__6444\ : CascadeMux
    port map (
            O => \N__36068\,
            I => \N__36062\
        );

    \I__6443\ : CascadeMux
    port map (
            O => \N__36065\,
            I => \N__36059\
        );

    \I__6442\ : CascadeBuf
    port map (
            O => \N__36062\,
            I => \N__36056\
        );

    \I__6441\ : CascadeBuf
    port map (
            O => \N__36059\,
            I => \N__36053\
        );

    \I__6440\ : CascadeMux
    port map (
            O => \N__36056\,
            I => \N__36050\
        );

    \I__6439\ : CascadeMux
    port map (
            O => \N__36053\,
            I => \N__36047\
        );

    \I__6438\ : CascadeBuf
    port map (
            O => \N__36050\,
            I => \N__36044\
        );

    \I__6437\ : CascadeBuf
    port map (
            O => \N__36047\,
            I => \N__36041\
        );

    \I__6436\ : CascadeMux
    port map (
            O => \N__36044\,
            I => \N__36038\
        );

    \I__6435\ : CascadeMux
    port map (
            O => \N__36041\,
            I => \N__36035\
        );

    \I__6434\ : CascadeBuf
    port map (
            O => \N__36038\,
            I => \N__36032\
        );

    \I__6433\ : CascadeBuf
    port map (
            O => \N__36035\,
            I => \N__36029\
        );

    \I__6432\ : CascadeMux
    port map (
            O => \N__36032\,
            I => \N__36026\
        );

    \I__6431\ : CascadeMux
    port map (
            O => \N__36029\,
            I => \N__36023\
        );

    \I__6430\ : InMux
    port map (
            O => \N__36026\,
            I => \N__36020\
        );

    \I__6429\ : InMux
    port map (
            O => \N__36023\,
            I => \N__36017\
        );

    \I__6428\ : LocalMux
    port map (
            O => \N__36020\,
            I => \N__36014\
        );

    \I__6427\ : LocalMux
    port map (
            O => \N__36017\,
            I => \N__36011\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__36014\,
            I => \N__36006\
        );

    \I__6425\ : Span4Mux_h
    port map (
            O => \N__36011\,
            I => \N__36006\
        );

    \I__6424\ : Span4Mux_h
    port map (
            O => \N__36006\,
            I => \N__36003\
        );

    \I__6423\ : Span4Mux_h
    port map (
            O => \N__36003\,
            I => \N__36000\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__36000\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1831_0\
        );

    \I__6421\ : CascadeMux
    port map (
            O => \N__35997\,
            I => \N__35993\
        );

    \I__6420\ : InMux
    port map (
            O => \N__35996\,
            I => \N__35983\
        );

    \I__6419\ : InMux
    port map (
            O => \N__35993\,
            I => \N__35974\
        );

    \I__6418\ : InMux
    port map (
            O => \N__35992\,
            I => \N__35974\
        );

    \I__6417\ : InMux
    port map (
            O => \N__35991\,
            I => \N__35974\
        );

    \I__6416\ : InMux
    port map (
            O => \N__35990\,
            I => \N__35974\
        );

    \I__6415\ : InMux
    port map (
            O => \N__35989\,
            I => \N__35968\
        );

    \I__6414\ : InMux
    port map (
            O => \N__35988\,
            I => \N__35968\
        );

    \I__6413\ : InMux
    port map (
            O => \N__35987\,
            I => \N__35963\
        );

    \I__6412\ : InMux
    port map (
            O => \N__35986\,
            I => \N__35963\
        );

    \I__6411\ : LocalMux
    port map (
            O => \N__35983\,
            I => \N__35960\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__35974\,
            I => \N__35957\
        );

    \I__6409\ : InMux
    port map (
            O => \N__35973\,
            I => \N__35954\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__35968\,
            I => \N__35949\
        );

    \I__6407\ : LocalMux
    port map (
            O => \N__35963\,
            I => \N__35949\
        );

    \I__6406\ : Span4Mux_v
    port map (
            O => \N__35960\,
            I => \N__35944\
        );

    \I__6405\ : Span4Mux_v
    port map (
            O => \N__35957\,
            I => \N__35944\
        );

    \I__6404\ : LocalMux
    port map (
            O => \N__35954\,
            I => \N__35941\
        );

    \I__6403\ : Span4Mux_v
    port map (
            O => \N__35949\,
            I => \N__35938\
        );

    \I__6402\ : Span4Mux_h
    port map (
            O => \N__35944\,
            I => \N__35935\
        );

    \I__6401\ : Span4Mux_h
    port map (
            O => \N__35941\,
            I => \N__35930\
        );

    \I__6400\ : Span4Mux_v
    port map (
            O => \N__35938\,
            I => \N__35930\
        );

    \I__6399\ : Odrv4
    port map (
            O => \N__35935\,
            I => \N_1614\
        );

    \I__6398\ : Odrv4
    port map (
            O => \N__35930\,
            I => \N_1614\
        );

    \I__6397\ : CascadeMux
    port map (
            O => \N__35925\,
            I => \N_1841_0_cascade_\
        );

    \I__6396\ : InMux
    port map (
            O => \N__35922\,
            I => \N__35919\
        );

    \I__6395\ : LocalMux
    port map (
            O => \N__35919\,
            I => \N__35916\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__35916\,
            I => \N__35912\
        );

    \I__6393\ : InMux
    port map (
            O => \N__35915\,
            I => \N__35909\
        );

    \I__6392\ : Span4Mux_v
    port map (
            O => \N__35912\,
            I => \N__35906\
        );

    \I__6391\ : LocalMux
    port map (
            O => \N__35909\,
            I => \N__35903\
        );

    \I__6390\ : Span4Mux_v
    port map (
            O => \N__35906\,
            I => \N__35900\
        );

    \I__6389\ : Sp12to4
    port map (
            O => \N__35903\,
            I => \N__35897\
        );

    \I__6388\ : Odrv4
    port map (
            O => \N__35900\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0\
        );

    \I__6387\ : Odrv12
    port map (
            O => \N__35897\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0\
        );

    \I__6386\ : InMux
    port map (
            O => \N__35892\,
            I => \N__35889\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__35889\,
            I => \N__35885\
        );

    \I__6384\ : InMux
    port map (
            O => \N__35888\,
            I => \N__35882\
        );

    \I__6383\ : Span4Mux_h
    port map (
            O => \N__35885\,
            I => \N__35878\
        );

    \I__6382\ : LocalMux
    port map (
            O => \N__35882\,
            I => \N__35875\
        );

    \I__6381\ : InMux
    port map (
            O => \N__35881\,
            I => \N__35872\
        );

    \I__6380\ : Span4Mux_v
    port map (
            O => \N__35878\,
            I => \N__35869\
        );

    \I__6379\ : Odrv4
    port map (
            O => \N__35875\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4\
        );

    \I__6378\ : LocalMux
    port map (
            O => \N__35872\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4\
        );

    \I__6377\ : Odrv4
    port map (
            O => \N__35869\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4\
        );

    \I__6376\ : InMux
    port map (
            O => \N__35862\,
            I => \N__35857\
        );

    \I__6375\ : InMux
    port map (
            O => \N__35861\,
            I => \N__35848\
        );

    \I__6374\ : InMux
    port map (
            O => \N__35860\,
            I => \N__35848\
        );

    \I__6373\ : LocalMux
    port map (
            O => \N__35857\,
            I => \N__35845\
        );

    \I__6372\ : InMux
    port map (
            O => \N__35856\,
            I => \N__35838\
        );

    \I__6371\ : InMux
    port map (
            O => \N__35855\,
            I => \N__35838\
        );

    \I__6370\ : InMux
    port map (
            O => \N__35854\,
            I => \N__35838\
        );

    \I__6369\ : InMux
    port map (
            O => \N__35853\,
            I => \N__35835\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__35848\,
            I => \N__35832\
        );

    \I__6367\ : Span4Mux_h
    port map (
            O => \N__35845\,
            I => \N__35829\
        );

    \I__6366\ : LocalMux
    port map (
            O => \N__35838\,
            I => \N__35826\
        );

    \I__6365\ : LocalMux
    port map (
            O => \N__35835\,
            I => \N__35823\
        );

    \I__6364\ : Span4Mux_v
    port map (
            O => \N__35832\,
            I => \N__35820\
        );

    \I__6363\ : Span4Mux_v
    port map (
            O => \N__35829\,
            I => \N__35813\
        );

    \I__6362\ : Span4Mux_h
    port map (
            O => \N__35826\,
            I => \N__35813\
        );

    \I__6361\ : Span4Mux_v
    port map (
            O => \N__35823\,
            I => \N__35808\
        );

    \I__6360\ : Span4Mux_h
    port map (
            O => \N__35820\,
            I => \N__35808\
        );

    \I__6359\ : InMux
    port map (
            O => \N__35819\,
            I => \N__35803\
        );

    \I__6358\ : InMux
    port map (
            O => \N__35818\,
            I => \N__35803\
        );

    \I__6357\ : Odrv4
    port map (
            O => \N__35813\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_b\
        );

    \I__6356\ : Odrv4
    port map (
            O => \N__35808\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_b\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__35803\,
            I => \cemf_module_64ch_ctrl_inst1.start_conf_b\
        );

    \I__6354\ : InMux
    port map (
            O => \N__35796\,
            I => \N__35792\
        );

    \I__6353\ : InMux
    port map (
            O => \N__35795\,
            I => \N__35789\
        );

    \I__6352\ : LocalMux
    port map (
            O => \N__35792\,
            I => \N__35786\
        );

    \I__6351\ : LocalMux
    port map (
            O => \N__35789\,
            I => \N__35783\
        );

    \I__6350\ : Span4Mux_v
    port map (
            O => \N__35786\,
            I => \N__35780\
        );

    \I__6349\ : Sp12to4
    port map (
            O => \N__35783\,
            I => \N__35777\
        );

    \I__6348\ : Span4Mux_v
    port map (
            O => \N__35780\,
            I => \N__35774\
        );

    \I__6347\ : Span12Mux_v
    port map (
            O => \N__35777\,
            I => \N__35771\
        );

    \I__6346\ : Sp12to4
    port map (
            O => \N__35774\,
            I => \N__35768\
        );

    \I__6345\ : Odrv12
    port map (
            O => \N__35771\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0\
        );

    \I__6344\ : Odrv12
    port map (
            O => \N__35768\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0\
        );

    \I__6343\ : CascadeMux
    port map (
            O => \N__35763\,
            I => \N__35758\
        );

    \I__6342\ : InMux
    port map (
            O => \N__35762\,
            I => \N__35752\
        );

    \I__6341\ : InMux
    port map (
            O => \N__35761\,
            I => \N__35749\
        );

    \I__6340\ : InMux
    port map (
            O => \N__35758\,
            I => \N__35743\
        );

    \I__6339\ : InMux
    port map (
            O => \N__35757\,
            I => \N__35743\
        );

    \I__6338\ : InMux
    port map (
            O => \N__35756\,
            I => \N__35738\
        );

    \I__6337\ : InMux
    port map (
            O => \N__35755\,
            I => \N__35738\
        );

    \I__6336\ : LocalMux
    port map (
            O => \N__35752\,
            I => \N__35735\
        );

    \I__6335\ : LocalMux
    port map (
            O => \N__35749\,
            I => \N__35732\
        );

    \I__6334\ : InMux
    port map (
            O => \N__35748\,
            I => \N__35729\
        );

    \I__6333\ : LocalMux
    port map (
            O => \N__35743\,
            I => \N__35726\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__35738\,
            I => \N__35719\
        );

    \I__6331\ : Span4Mux_v
    port map (
            O => \N__35735\,
            I => \N__35719\
        );

    \I__6330\ : Sp12to4
    port map (
            O => \N__35732\,
            I => \N__35716\
        );

    \I__6329\ : LocalMux
    port map (
            O => \N__35729\,
            I => \N__35711\
        );

    \I__6328\ : Span4Mux_h
    port map (
            O => \N__35726\,
            I => \N__35711\
        );

    \I__6327\ : InMux
    port map (
            O => \N__35725\,
            I => \N__35708\
        );

    \I__6326\ : InMux
    port map (
            O => \N__35724\,
            I => \N__35705\
        );

    \I__6325\ : Sp12to4
    port map (
            O => \N__35719\,
            I => \N__35700\
        );

    \I__6324\ : Span12Mux_v
    port map (
            O => \N__35716\,
            I => \N__35700\
        );

    \I__6323\ : Odrv4
    port map (
            O => \N__35711\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15\
        );

    \I__6322\ : LocalMux
    port map (
            O => \N__35708\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15\
        );

    \I__6321\ : LocalMux
    port map (
            O => \N__35705\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15\
        );

    \I__6320\ : Odrv12
    port map (
            O => \N__35700\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15\
        );

    \I__6319\ : InMux
    port map (
            O => \N__35691\,
            I => \N__35688\
        );

    \I__6318\ : LocalMux
    port map (
            O => \N__35688\,
            I => \N__35685\
        );

    \I__6317\ : Span4Mux_v
    port map (
            O => \N__35685\,
            I => \N__35682\
        );

    \I__6316\ : Sp12to4
    port map (
            O => \N__35682\,
            I => \N__35677\
        );

    \I__6315\ : InMux
    port map (
            O => \N__35681\,
            I => \N__35672\
        );

    \I__6314\ : InMux
    port map (
            O => \N__35680\,
            I => \N__35672\
        );

    \I__6313\ : Odrv12
    port map (
            O => \N__35677\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_20
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__35672\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_20
        );

    \I__6311\ : CascadeMux
    port map (
            O => \N__35667\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_20_cascade_\
        );

    \I__6310\ : CascadeMux
    port map (
            O => \N__35664\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DDZ0Z7_cascade_\
        );

    \I__6309\ : InMux
    port map (
            O => \N__35661\,
            I => \N__35658\
        );

    \I__6308\ : LocalMux
    port map (
            O => \N__35658\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20\
        );

    \I__6307\ : InMux
    port map (
            O => \N__35655\,
            I => \N__35652\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__35652\,
            I => \N__35648\
        );

    \I__6305\ : InMux
    port map (
            O => \N__35651\,
            I => \N__35645\
        );

    \I__6304\ : Span4Mux_v
    port map (
            O => \N__35648\,
            I => \N__35642\
        );

    \I__6303\ : LocalMux
    port map (
            O => \N__35645\,
            I => \N__35639\
        );

    \I__6302\ : Span4Mux_h
    port map (
            O => \N__35642\,
            I => \N__35636\
        );

    \I__6301\ : Odrv4
    port map (
            O => \N__35639\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_28
        );

    \I__6300\ : Odrv4
    port map (
            O => \N__35636\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_28
        );

    \I__6299\ : InMux
    port map (
            O => \N__35631\,
            I => \N__35628\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__35628\,
            I => \N__35625\
        );

    \I__6297\ : Span4Mux_h
    port map (
            O => \N__35625\,
            I => \N__35622\
        );

    \I__6296\ : Odrv4
    port map (
            O => \N__35622\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_28\
        );

    \I__6295\ : CascadeMux
    port map (
            O => \N__35619\,
            I => \N__35616\
        );

    \I__6294\ : InMux
    port map (
            O => \N__35616\,
            I => \N__35613\
        );

    \I__6293\ : LocalMux
    port map (
            O => \N__35613\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_28\
        );

    \I__6292\ : InMux
    port map (
            O => \N__35610\,
            I => \N__35607\
        );

    \I__6291\ : LocalMux
    port map (
            O => \N__35607\,
            I => \N__35604\
        );

    \I__6290\ : Span4Mux_v
    port map (
            O => \N__35604\,
            I => \N__35600\
        );

    \I__6289\ : InMux
    port map (
            O => \N__35603\,
            I => \N__35597\
        );

    \I__6288\ : Span4Mux_h
    port map (
            O => \N__35600\,
            I => \N__35594\
        );

    \I__6287\ : LocalMux
    port map (
            O => \N__35597\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_29
        );

    \I__6286\ : Odrv4
    port map (
            O => \N__35594\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_29
        );

    \I__6285\ : CascadeMux
    port map (
            O => \N__35589\,
            I => \N__35586\
        );

    \I__6284\ : InMux
    port map (
            O => \N__35586\,
            I => \N__35583\
        );

    \I__6283\ : LocalMux
    port map (
            O => \N__35583\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_29\
        );

    \I__6282\ : InMux
    port map (
            O => \N__35580\,
            I => \N__35577\
        );

    \I__6281\ : LocalMux
    port map (
            O => \N__35577\,
            I => \N__35574\
        );

    \I__6280\ : Span4Mux_v
    port map (
            O => \N__35574\,
            I => \N__35570\
        );

    \I__6279\ : CascadeMux
    port map (
            O => \N__35573\,
            I => \N__35567\
        );

    \I__6278\ : Span4Mux_h
    port map (
            O => \N__35570\,
            I => \N__35564\
        );

    \I__6277\ : InMux
    port map (
            O => \N__35567\,
            I => \N__35561\
        );

    \I__6276\ : Sp12to4
    port map (
            O => \N__35564\,
            I => \N__35558\
        );

    \I__6275\ : LocalMux
    port map (
            O => \N__35561\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_3
        );

    \I__6274\ : Odrv12
    port map (
            O => \N__35558\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_3
        );

    \I__6273\ : InMux
    port map (
            O => \N__35553\,
            I => \N__35550\
        );

    \I__6272\ : LocalMux
    port map (
            O => \N__35550\,
            I => \N__35547\
        );

    \I__6271\ : Span4Mux_h
    port map (
            O => \N__35547\,
            I => \N__35544\
        );

    \I__6270\ : Span4Mux_h
    port map (
            O => \N__35544\,
            I => \N__35541\
        );

    \I__6269\ : Odrv4
    port map (
            O => \N__35541\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_3\
        );

    \I__6268\ : CascadeMux
    port map (
            O => \N__35538\,
            I => \N__35534\
        );

    \I__6267\ : InMux
    port map (
            O => \N__35537\,
            I => \N__35530\
        );

    \I__6266\ : InMux
    port map (
            O => \N__35534\,
            I => \N__35527\
        );

    \I__6265\ : CascadeMux
    port map (
            O => \N__35533\,
            I => \N__35524\
        );

    \I__6264\ : LocalMux
    port map (
            O => \N__35530\,
            I => \N__35519\
        );

    \I__6263\ : LocalMux
    port map (
            O => \N__35527\,
            I => \N__35519\
        );

    \I__6262\ : InMux
    port map (
            O => \N__35524\,
            I => \N__35516\
        );

    \I__6261\ : Span4Mux_h
    port map (
            O => \N__35519\,
            I => \N__35513\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__35516\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_3
        );

    \I__6259\ : Odrv4
    port map (
            O => \N__35513\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_3
        );

    \I__6258\ : IoInMux
    port map (
            O => \N__35508\,
            I => \N__35505\
        );

    \I__6257\ : LocalMux
    port map (
            O => \N__35505\,
            I => \N__35502\
        );

    \I__6256\ : IoSpan4Mux
    port map (
            O => \N__35502\,
            I => \N__35499\
        );

    \I__6255\ : Span4Mux_s2_h
    port map (
            O => \N__35499\,
            I => \N__35496\
        );

    \I__6254\ : Sp12to4
    port map (
            O => \N__35496\,
            I => \N__35493\
        );

    \I__6253\ : Span12Mux_h
    port map (
            O => \N__35493\,
            I => \N__35490\
        );

    \I__6252\ : Odrv12
    port map (
            O => \N__35490\,
            I => serial_out_testing_c
        );

    \I__6251\ : CascadeMux
    port map (
            O => \N__35487\,
            I => \N__35484\
        );

    \I__6250\ : InMux
    port map (
            O => \N__35484\,
            I => \N__35474\
        );

    \I__6249\ : InMux
    port map (
            O => \N__35483\,
            I => \N__35474\
        );

    \I__6248\ : InMux
    port map (
            O => \N__35482\,
            I => \N__35474\
        );

    \I__6247\ : CEMux
    port map (
            O => \N__35481\,
            I => \N__35471\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__35474\,
            I => \N__35468\
        );

    \I__6245\ : LocalMux
    port map (
            O => \N__35471\,
            I => \N__35465\
        );

    \I__6244\ : Span4Mux_h
    port map (
            O => \N__35468\,
            I => \N__35461\
        );

    \I__6243\ : Span4Mux_h
    port map (
            O => \N__35465\,
            I => \N__35458\
        );

    \I__6242\ : InMux
    port map (
            O => \N__35464\,
            I => \N__35454\
        );

    \I__6241\ : Span4Mux_h
    port map (
            O => \N__35461\,
            I => \N__35451\
        );

    \I__6240\ : Span4Mux_h
    port map (
            O => \N__35458\,
            I => \N__35448\
        );

    \I__6239\ : InMux
    port map (
            O => \N__35457\,
            I => \N__35445\
        );

    \I__6238\ : LocalMux
    port map (
            O => \N__35454\,
            I => \N__35442\
        );

    \I__6237\ : Sp12to4
    port map (
            O => \N__35451\,
            I => \N__35439\
        );

    \I__6236\ : Span4Mux_h
    port map (
            O => \N__35448\,
            I => \N__35436\
        );

    \I__6235\ : LocalMux
    port map (
            O => \N__35445\,
            I => \N__35433\
        );

    \I__6234\ : Span4Mux_h
    port map (
            O => \N__35442\,
            I => \N__35430\
        );

    \I__6233\ : Span12Mux_v
    port map (
            O => \N__35439\,
            I => \N__35427\
        );

    \I__6232\ : Sp12to4
    port map (
            O => \N__35436\,
            I => \N__35424\
        );

    \I__6231\ : Span12Mux_h
    port map (
            O => \N__35433\,
            I => \N__35421\
        );

    \I__6230\ : Span4Mux_h
    port map (
            O => \N__35430\,
            I => \N__35418\
        );

    \I__6229\ : Span12Mux_h
    port map (
            O => \N__35427\,
            I => \N__35415\
        );

    \I__6228\ : Span12Mux_v
    port map (
            O => \N__35424\,
            I => \N__35410\
        );

    \I__6227\ : Span12Mux_h
    port map (
            O => \N__35421\,
            I => \N__35410\
        );

    \I__6226\ : Span4Mux_h
    port map (
            O => \N__35418\,
            I => \N__35407\
        );

    \I__6225\ : Odrv12
    port map (
            O => \N__35415\,
            I => rst_n_c
        );

    \I__6224\ : Odrv12
    port map (
            O => \N__35410\,
            I => rst_n_c
        );

    \I__6223\ : Odrv4
    port map (
            O => \N__35407\,
            I => rst_n_c
        );

    \I__6222\ : InMux
    port map (
            O => \N__35400\,
            I => \N__35397\
        );

    \I__6221\ : LocalMux
    port map (
            O => \N__35397\,
            I => \N__35391\
        );

    \I__6220\ : InMux
    port map (
            O => \N__35396\,
            I => \N__35388\
        );

    \I__6219\ : InMux
    port map (
            O => \N__35395\,
            I => \N__35383\
        );

    \I__6218\ : InMux
    port map (
            O => \N__35394\,
            I => \N__35383\
        );

    \I__6217\ : Span4Mux_h
    port map (
            O => \N__35391\,
            I => \N__35380\
        );

    \I__6216\ : LocalMux
    port map (
            O => \N__35388\,
            I => \N__35375\
        );

    \I__6215\ : LocalMux
    port map (
            O => \N__35383\,
            I => \N__35375\
        );

    \I__6214\ : Sp12to4
    port map (
            O => \N__35380\,
            I => \N__35370\
        );

    \I__6213\ : Span12Mux_h
    port map (
            O => \N__35375\,
            I => \N__35370\
        );

    \I__6212\ : Odrv12
    port map (
            O => \N__35370\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1965\
        );

    \I__6211\ : InMux
    port map (
            O => \N__35367\,
            I => \N__35364\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__35364\,
            I => \N__35361\
        );

    \I__6209\ : Span4Mux_v
    port map (
            O => \N__35361\,
            I => \N__35357\
        );

    \I__6208\ : InMux
    port map (
            O => \N__35360\,
            I => \N__35354\
        );

    \I__6207\ : Sp12to4
    port map (
            O => \N__35357\,
            I => \N__35351\
        );

    \I__6206\ : LocalMux
    port map (
            O => \N__35354\,
            I => \N__35348\
        );

    \I__6205\ : Span12Mux_h
    port map (
            O => \N__35351\,
            I => \N__35343\
        );

    \I__6204\ : Sp12to4
    port map (
            O => \N__35348\,
            I => \N__35343\
        );

    \I__6203\ : Odrv12
    port map (
            O => \N__35343\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_522_0\
        );

    \I__6202\ : CascadeMux
    port map (
            O => \N__35340\,
            I => \N__35337\
        );

    \I__6201\ : InMux
    port map (
            O => \N__35337\,
            I => \N__35334\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__35334\,
            I => \N__35331\
        );

    \I__6199\ : Span4Mux_h
    port map (
            O => \N__35331\,
            I => \N__35327\
        );

    \I__6198\ : InMux
    port map (
            O => \N__35330\,
            I => \N__35324\
        );

    \I__6197\ : Span4Mux_h
    port map (
            O => \N__35327\,
            I => \N__35321\
        );

    \I__6196\ : LocalMux
    port map (
            O => \N__35324\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_17
        );

    \I__6195\ : Odrv4
    port map (
            O => \N__35321\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_17
        );

    \I__6194\ : InMux
    port map (
            O => \N__35316\,
            I => \N__35313\
        );

    \I__6193\ : LocalMux
    port map (
            O => \N__35313\,
            I => \N__35310\
        );

    \I__6192\ : Span4Mux_h
    port map (
            O => \N__35310\,
            I => \N__35307\
        );

    \I__6191\ : Odrv4
    port map (
            O => \N__35307\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_17\
        );

    \I__6190\ : InMux
    port map (
            O => \N__35304\,
            I => \N__35300\
        );

    \I__6189\ : CascadeMux
    port map (
            O => \N__35303\,
            I => \N__35297\
        );

    \I__6188\ : LocalMux
    port map (
            O => \N__35300\,
            I => \N__35294\
        );

    \I__6187\ : InMux
    port map (
            O => \N__35297\,
            I => \N__35291\
        );

    \I__6186\ : Span4Mux_v
    port map (
            O => \N__35294\,
            I => \N__35288\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__35291\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_2
        );

    \I__6184\ : Odrv4
    port map (
            O => \N__35288\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_2
        );

    \I__6183\ : CascadeMux
    port map (
            O => \N__35283\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0_cascade_\
        );

    \I__6182\ : InMux
    port map (
            O => \N__35280\,
            I => \N__35277\
        );

    \I__6181\ : LocalMux
    port map (
            O => \N__35277\,
            I => \N__35274\
        );

    \I__6180\ : Span4Mux_h
    port map (
            O => \N__35274\,
            I => \N__35271\
        );

    \I__6179\ : Odrv4
    port map (
            O => \N__35271\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_2\
        );

    \I__6178\ : InMux
    port map (
            O => \N__35268\,
            I => \N__35265\
        );

    \I__6177\ : LocalMux
    port map (
            O => \N__35265\,
            I => \N__35261\
        );

    \I__6176\ : InMux
    port map (
            O => \N__35264\,
            I => \N__35258\
        );

    \I__6175\ : Span4Mux_h
    port map (
            O => \N__35261\,
            I => \N__35255\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__35258\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_24
        );

    \I__6173\ : Odrv4
    port map (
            O => \N__35255\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_24
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__35250\,
            I => \N__35247\
        );

    \I__6171\ : InMux
    port map (
            O => \N__35247\,
            I => \N__35244\
        );

    \I__6170\ : LocalMux
    port map (
            O => \N__35244\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_24\
        );

    \I__6169\ : CascadeMux
    port map (
            O => \N__35241\,
            I => \N__35238\
        );

    \I__6168\ : InMux
    port map (
            O => \N__35238\,
            I => \N__35235\
        );

    \I__6167\ : LocalMux
    port map (
            O => \N__35235\,
            I => \N__35231\
        );

    \I__6166\ : InMux
    port map (
            O => \N__35234\,
            I => \N__35228\
        );

    \I__6165\ : Sp12to4
    port map (
            O => \N__35231\,
            I => \N__35225\
        );

    \I__6164\ : LocalMux
    port map (
            O => \N__35228\,
            I => \N__35220\
        );

    \I__6163\ : Span12Mux_v
    port map (
            O => \N__35225\,
            I => \N__35220\
        );

    \I__6162\ : Odrv12
    port map (
            O => \N__35220\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_19
        );

    \I__6161\ : InMux
    port map (
            O => \N__35217\,
            I => \N__35214\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__35214\,
            I => \N__35211\
        );

    \I__6159\ : Span4Mux_v
    port map (
            O => \N__35211\,
            I => \N__35208\
        );

    \I__6158\ : Odrv4
    port map (
            O => \N__35208\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_19\
        );

    \I__6157\ : InMux
    port map (
            O => \N__35205\,
            I => \N__35202\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__35202\,
            I => \N__35199\
        );

    \I__6155\ : Span4Mux_v
    port map (
            O => \N__35199\,
            I => \N__35195\
        );

    \I__6154\ : InMux
    port map (
            O => \N__35198\,
            I => \N__35192\
        );

    \I__6153\ : Span4Mux_h
    port map (
            O => \N__35195\,
            I => \N__35189\
        );

    \I__6152\ : LocalMux
    port map (
            O => \N__35192\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_25
        );

    \I__6151\ : Odrv4
    port map (
            O => \N__35189\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_25
        );

    \I__6150\ : InMux
    port map (
            O => \N__35184\,
            I => \N__35181\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__35181\,
            I => \N__35178\
        );

    \I__6148\ : Span4Mux_h
    port map (
            O => \N__35178\,
            I => \N__35174\
        );

    \I__6147\ : InMux
    port map (
            O => \N__35177\,
            I => \N__35171\
        );

    \I__6146\ : Span4Mux_h
    port map (
            O => \N__35174\,
            I => \N__35168\
        );

    \I__6145\ : LocalMux
    port map (
            O => \N__35171\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_27
        );

    \I__6144\ : Odrv4
    port map (
            O => \N__35168\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_27
        );

    \I__6143\ : CascadeMux
    port map (
            O => \N__35163\,
            I => \N__35160\
        );

    \I__6142\ : InMux
    port map (
            O => \N__35160\,
            I => \N__35157\
        );

    \I__6141\ : LocalMux
    port map (
            O => \N__35157\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_27\
        );

    \I__6140\ : InMux
    port map (
            O => \N__35154\,
            I => \N__35151\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__35151\,
            I => \N__35148\
        );

    \I__6138\ : Span4Mux_h
    port map (
            O => \N__35148\,
            I => \N__35145\
        );

    \I__6137\ : Span4Mux_h
    port map (
            O => \N__35145\,
            I => \N__35142\
        );

    \I__6136\ : Span4Mux_h
    port map (
            O => \N__35142\,
            I => \N__35139\
        );

    \I__6135\ : Odrv4
    port map (
            O => \N__35139\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_12
        );

    \I__6134\ : InMux
    port map (
            O => \N__35136\,
            I => \N__35133\
        );

    \I__6133\ : LocalMux
    port map (
            O => \N__35133\,
            I => \N__35130\
        );

    \I__6132\ : Span12Mux_v
    port map (
            O => \N__35130\,
            I => \N__35127\
        );

    \I__6131\ : Odrv12
    port map (
            O => \N__35127\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_808\
        );

    \I__6130\ : CascadeMux
    port map (
            O => \N__35124\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_12_cascade_\
        );

    \I__6129\ : InMux
    port map (
            O => \N__35121\,
            I => \N__35118\
        );

    \I__6128\ : LocalMux
    port map (
            O => \N__35118\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_12\
        );

    \I__6127\ : CascadeMux
    port map (
            O => \N__35115\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_12_cascade_\
        );

    \I__6126\ : InMux
    port map (
            O => \N__35112\,
            I => \N__35109\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__35109\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_12\
        );

    \I__6124\ : CascadeMux
    port map (
            O => \N__35106\,
            I => \N__35103\
        );

    \I__6123\ : InMux
    port map (
            O => \N__35103\,
            I => \N__35100\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__35100\,
            I => \N__35096\
        );

    \I__6121\ : CascadeMux
    port map (
            O => \N__35099\,
            I => \N__35093\
        );

    \I__6120\ : Span4Mux_v
    port map (
            O => \N__35096\,
            I => \N__35090\
        );

    \I__6119\ : InMux
    port map (
            O => \N__35093\,
            I => \N__35087\
        );

    \I__6118\ : Span4Mux_v
    port map (
            O => \N__35090\,
            I => \N__35084\
        );

    \I__6117\ : LocalMux
    port map (
            O => \N__35087\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_11
        );

    \I__6116\ : Odrv4
    port map (
            O => \N__35084\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_11
        );

    \I__6115\ : InMux
    port map (
            O => \N__35079\,
            I => \N__35076\
        );

    \I__6114\ : LocalMux
    port map (
            O => \N__35076\,
            I => \N__35073\
        );

    \I__6113\ : Odrv4
    port map (
            O => \N__35073\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_11\
        );

    \I__6112\ : CascadeMux
    port map (
            O => \N__35070\,
            I => \N__35067\
        );

    \I__6111\ : InMux
    port map (
            O => \N__35067\,
            I => \N__35064\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__35064\,
            I => \N__35061\
        );

    \I__6109\ : Span4Mux_h
    port map (
            O => \N__35061\,
            I => \N__35057\
        );

    \I__6108\ : CascadeMux
    port map (
            O => \N__35060\,
            I => \N__35054\
        );

    \I__6107\ : Span4Mux_v
    port map (
            O => \N__35057\,
            I => \N__35051\
        );

    \I__6106\ : InMux
    port map (
            O => \N__35054\,
            I => \N__35048\
        );

    \I__6105\ : Sp12to4
    port map (
            O => \N__35051\,
            I => \N__35045\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__35048\,
            I => \N__35040\
        );

    \I__6103\ : Span12Mux_v
    port map (
            O => \N__35045\,
            I => \N__35040\
        );

    \I__6102\ : Odrv12
    port map (
            O => \N__35040\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_12
        );

    \I__6101\ : InMux
    port map (
            O => \N__35037\,
            I => \N__35034\
        );

    \I__6100\ : LocalMux
    port map (
            O => \N__35034\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_12\
        );

    \I__6099\ : CascadeMux
    port map (
            O => \N__35031\,
            I => \N__35028\
        );

    \I__6098\ : InMux
    port map (
            O => \N__35028\,
            I => \N__35025\
        );

    \I__6097\ : LocalMux
    port map (
            O => \N__35025\,
            I => \N__35022\
        );

    \I__6096\ : Span4Mux_v
    port map (
            O => \N__35022\,
            I => \N__35019\
        );

    \I__6095\ : Span4Mux_v
    port map (
            O => \N__35019\,
            I => \N__35015\
        );

    \I__6094\ : InMux
    port map (
            O => \N__35018\,
            I => \N__35012\
        );

    \I__6093\ : Sp12to4
    port map (
            O => \N__35015\,
            I => \N__35009\
        );

    \I__6092\ : LocalMux
    port map (
            O => \N__35012\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_13
        );

    \I__6091\ : Odrv12
    port map (
            O => \N__35009\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_13
        );

    \I__6090\ : InMux
    port map (
            O => \N__35004\,
            I => \N__35001\
        );

    \I__6089\ : LocalMux
    port map (
            O => \N__35001\,
            I => \N__34998\
        );

    \I__6088\ : Span4Mux_h
    port map (
            O => \N__34998\,
            I => \N__34995\
        );

    \I__6087\ : Odrv4
    port map (
            O => \N__34995\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_13\
        );

    \I__6086\ : CascadeMux
    port map (
            O => \N__34992\,
            I => \N__34989\
        );

    \I__6085\ : InMux
    port map (
            O => \N__34989\,
            I => \N__34985\
        );

    \I__6084\ : CascadeMux
    port map (
            O => \N__34988\,
            I => \N__34982\
        );

    \I__6083\ : LocalMux
    port map (
            O => \N__34985\,
            I => \N__34979\
        );

    \I__6082\ : InMux
    port map (
            O => \N__34982\,
            I => \N__34976\
        );

    \I__6081\ : Span12Mux_v
    port map (
            O => \N__34979\,
            I => \N__34973\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__34976\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_14
        );

    \I__6079\ : Odrv12
    port map (
            O => \N__34973\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_14
        );

    \I__6078\ : InMux
    port map (
            O => \N__34968\,
            I => \N__34965\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__34965\,
            I => \N__34962\
        );

    \I__6076\ : Span4Mux_h
    port map (
            O => \N__34962\,
            I => \N__34959\
        );

    \I__6075\ : Span4Mux_h
    port map (
            O => \N__34959\,
            I => \N__34956\
        );

    \I__6074\ : Odrv4
    port map (
            O => \N__34956\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_14\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__34953\,
            I => \N__34950\
        );

    \I__6072\ : InMux
    port map (
            O => \N__34950\,
            I => \N__34947\
        );

    \I__6071\ : LocalMux
    port map (
            O => \N__34947\,
            I => \N__34944\
        );

    \I__6070\ : Span4Mux_h
    port map (
            O => \N__34944\,
            I => \N__34940\
        );

    \I__6069\ : CascadeMux
    port map (
            O => \N__34943\,
            I => \N__34937\
        );

    \I__6068\ : Span4Mux_v
    port map (
            O => \N__34940\,
            I => \N__34934\
        );

    \I__6067\ : InMux
    port map (
            O => \N__34937\,
            I => \N__34931\
        );

    \I__6066\ : Span4Mux_v
    port map (
            O => \N__34934\,
            I => \N__34928\
        );

    \I__6065\ : LocalMux
    port map (
            O => \N__34931\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_15
        );

    \I__6064\ : Odrv4
    port map (
            O => \N__34928\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_15
        );

    \I__6063\ : InMux
    port map (
            O => \N__34923\,
            I => \N__34920\
        );

    \I__6062\ : LocalMux
    port map (
            O => \N__34920\,
            I => \N__34917\
        );

    \I__6061\ : Odrv12
    port map (
            O => \N__34917\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_15\
        );

    \I__6060\ : CascadeMux
    port map (
            O => \N__34914\,
            I => \N__34911\
        );

    \I__6059\ : InMux
    port map (
            O => \N__34911\,
            I => \N__34907\
        );

    \I__6058\ : CascadeMux
    port map (
            O => \N__34910\,
            I => \N__34904\
        );

    \I__6057\ : LocalMux
    port map (
            O => \N__34907\,
            I => \N__34901\
        );

    \I__6056\ : InMux
    port map (
            O => \N__34904\,
            I => \N__34898\
        );

    \I__6055\ : Span4Mux_v
    port map (
            O => \N__34901\,
            I => \N__34895\
        );

    \I__6054\ : LocalMux
    port map (
            O => \N__34898\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_16
        );

    \I__6053\ : Odrv4
    port map (
            O => \N__34895\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_16
        );

    \I__6052\ : InMux
    port map (
            O => \N__34890\,
            I => \N__34887\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__34887\,
            I => \serializer_mod_inst.shift_regZ0Z_67\
        );

    \I__6050\ : InMux
    port map (
            O => \N__34884\,
            I => \N__34881\
        );

    \I__6049\ : LocalMux
    port map (
            O => \N__34881\,
            I => \serializer_mod_inst.shift_regZ0Z_68\
        );

    \I__6048\ : InMux
    port map (
            O => \N__34878\,
            I => \N__34875\
        );

    \I__6047\ : LocalMux
    port map (
            O => \N__34875\,
            I => \N__34872\
        );

    \I__6046\ : Odrv4
    port map (
            O => \N__34872\,
            I => \serializer_mod_inst.shift_regZ0Z_115\
        );

    \I__6045\ : InMux
    port map (
            O => \N__34869\,
            I => \N__34866\
        );

    \I__6044\ : LocalMux
    port map (
            O => \N__34866\,
            I => \serializer_mod_inst.shift_regZ0Z_116\
        );

    \I__6043\ : InMux
    port map (
            O => \N__34863\,
            I => \N__34860\
        );

    \I__6042\ : LocalMux
    port map (
            O => \N__34860\,
            I => \serializer_mod_inst.shift_regZ0Z_117\
        );

    \I__6041\ : InMux
    port map (
            O => \N__34857\,
            I => \N__34853\
        );

    \I__6040\ : InMux
    port map (
            O => \N__34856\,
            I => \N__34848\
        );

    \I__6039\ : LocalMux
    port map (
            O => \N__34853\,
            I => \N__34845\
        );

    \I__6038\ : InMux
    port map (
            O => \N__34852\,
            I => \N__34840\
        );

    \I__6037\ : InMux
    port map (
            O => \N__34851\,
            I => \N__34837\
        );

    \I__6036\ : LocalMux
    port map (
            O => \N__34848\,
            I => \N__34832\
        );

    \I__6035\ : Span12Mux_s6_v
    port map (
            O => \N__34845\,
            I => \N__34832\
        );

    \I__6034\ : InMux
    port map (
            O => \N__34844\,
            I => \N__34827\
        );

    \I__6033\ : InMux
    port map (
            O => \N__34843\,
            I => \N__34827\
        );

    \I__6032\ : LocalMux
    port map (
            O => \N__34840\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0\
        );

    \I__6031\ : LocalMux
    port map (
            O => \N__34837\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0\
        );

    \I__6030\ : Odrv12
    port map (
            O => \N__34832\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__34827\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0\
        );

    \I__6028\ : IoInMux
    port map (
            O => \N__34818\,
            I => \N__34815\
        );

    \I__6027\ : LocalMux
    port map (
            O => \N__34815\,
            I => \N__34812\
        );

    \I__6026\ : Span4Mux_s2_v
    port map (
            O => \N__34812\,
            I => \N__34809\
        );

    \I__6025\ : Odrv4
    port map (
            O => \N__34809\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa\
        );

    \I__6024\ : IoInMux
    port map (
            O => \N__34806\,
            I => \N__34803\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__34803\,
            I => rst_n_c_i
        );

    \I__6022\ : InMux
    port map (
            O => \N__34800\,
            I => \N__34797\
        );

    \I__6021\ : LocalMux
    port map (
            O => \N__34797\,
            I => \N__34794\
        );

    \I__6020\ : Span4Mux_h
    port map (
            O => \N__34794\,
            I => \N__34791\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__34791\,
            I => \N__34788\
        );

    \I__6018\ : Span4Mux_v
    port map (
            O => \N__34788\,
            I => \N__34785\
        );

    \I__6017\ : Span4Mux_v
    port map (
            O => \N__34785\,
            I => \N__34782\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__34782\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_12
        );

    \I__6015\ : CascadeMux
    port map (
            O => \N__34779\,
            I => \N__34776\
        );

    \I__6014\ : InMux
    port map (
            O => \N__34776\,
            I => \N__34773\
        );

    \I__6013\ : LocalMux
    port map (
            O => \N__34773\,
            I => \N__34770\
        );

    \I__6012\ : Span4Mux_h
    port map (
            O => \N__34770\,
            I => \N__34767\
        );

    \I__6011\ : Span4Mux_v
    port map (
            O => \N__34767\,
            I => \N__34764\
        );

    \I__6010\ : Span4Mux_h
    port map (
            O => \N__34764\,
            I => \N__34761\
        );

    \I__6009\ : Odrv4
    port map (
            O => \N__34761\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_12
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__34758\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_12_cascade_\
        );

    \I__6007\ : InMux
    port map (
            O => \N__34755\,
            I => \N__34752\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__34752\,
            I => \N__34749\
        );

    \I__6005\ : Odrv4
    port map (
            O => \N__34749\,
            I => \serializer_mod_inst.shift_regZ0Z_113\
        );

    \I__6004\ : InMux
    port map (
            O => \N__34746\,
            I => \N__34743\
        );

    \I__6003\ : LocalMux
    port map (
            O => \N__34743\,
            I => \serializer_mod_inst.shift_regZ0Z_114\
        );

    \I__6002\ : InMux
    port map (
            O => \N__34740\,
            I => \N__34737\
        );

    \I__6001\ : LocalMux
    port map (
            O => \N__34737\,
            I => \serializer_mod_inst.shift_regZ0Z_110\
        );

    \I__6000\ : InMux
    port map (
            O => \N__34734\,
            I => \N__34731\
        );

    \I__5999\ : LocalMux
    port map (
            O => \N__34731\,
            I => \serializer_mod_inst.shift_regZ0Z_39\
        );

    \I__5998\ : InMux
    port map (
            O => \N__34728\,
            I => \N__34725\
        );

    \I__5997\ : LocalMux
    port map (
            O => \N__34725\,
            I => \serializer_mod_inst.shift_regZ0Z_77\
        );

    \I__5996\ : InMux
    port map (
            O => \N__34722\,
            I => \N__34719\
        );

    \I__5995\ : LocalMux
    port map (
            O => \N__34719\,
            I => \serializer_mod_inst.shift_regZ0Z_78\
        );

    \I__5994\ : InMux
    port map (
            O => \N__34716\,
            I => \N__34713\
        );

    \I__5993\ : LocalMux
    port map (
            O => \N__34713\,
            I => \serializer_mod_inst.shift_regZ0Z_40\
        );

    \I__5992\ : CascadeMux
    port map (
            O => \N__34710\,
            I => \N__34707\
        );

    \I__5991\ : InMux
    port map (
            O => \N__34707\,
            I => \N__34704\
        );

    \I__5990\ : LocalMux
    port map (
            O => \N__34704\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0\
        );

    \I__5989\ : InMux
    port map (
            O => \N__34701\,
            I => \N__34698\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__34698\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_2\
        );

    \I__5987\ : InMux
    port map (
            O => \N__34695\,
            I => \N__34692\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__34692\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_12\
        );

    \I__5985\ : InMux
    port map (
            O => \N__34689\,
            I => \N__34686\
        );

    \I__5984\ : LocalMux
    port map (
            O => \N__34686\,
            I => \N__34683\
        );

    \I__5983\ : Odrv4
    port map (
            O => \N__34683\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_li_0_1\
        );

    \I__5982\ : InMux
    port map (
            O => \N__34680\,
            I => \N__34677\
        );

    \I__5981\ : LocalMux
    port map (
            O => \N__34677\,
            I => \c_state_ret_12_RNIDMPS1_0\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__34674\,
            I => \c_state_ret_12_RNIDMPS1_0_cascade_\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__34671\,
            I => \N__34667\
        );

    \I__5978\ : InMux
    port map (
            O => \N__34670\,
            I => \N__34662\
        );

    \I__5977\ : InMux
    port map (
            O => \N__34667\,
            I => \N__34662\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__34662\,
            I => \N__34659\
        );

    \I__5975\ : Span4Mux_v
    port map (
            O => \N__34659\,
            I => \N__34656\
        );

    \I__5974\ : Span4Mux_v
    port map (
            O => \N__34656\,
            I => \N__34651\
        );

    \I__5973\ : InMux
    port map (
            O => \N__34655\,
            I => \N__34646\
        );

    \I__5972\ : InMux
    port map (
            O => \N__34654\,
            I => \N__34646\
        );

    \I__5971\ : Odrv4
    port map (
            O => \N__34651\,
            I => \cemf_module_64ch_ctrl_inst1.clr_sys_reg\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__34646\,
            I => \cemf_module_64ch_ctrl_inst1.clr_sys_reg\
        );

    \I__5969\ : CascadeMux
    port map (
            O => \N__34641\,
            I => \N__34636\
        );

    \I__5968\ : CascadeMux
    port map (
            O => \N__34640\,
            I => \N__34633\
        );

    \I__5967\ : CascadeMux
    port map (
            O => \N__34639\,
            I => \N__34630\
        );

    \I__5966\ : InMux
    port map (
            O => \N__34636\,
            I => \N__34626\
        );

    \I__5965\ : InMux
    port map (
            O => \N__34633\,
            I => \N__34621\
        );

    \I__5964\ : InMux
    port map (
            O => \N__34630\,
            I => \N__34621\
        );

    \I__5963\ : InMux
    port map (
            O => \N__34629\,
            I => \N__34618\
        );

    \I__5962\ : LocalMux
    port map (
            O => \N__34626\,
            I => \N__34615\
        );

    \I__5961\ : LocalMux
    port map (
            O => \N__34621\,
            I => \N__34612\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__34618\,
            I => \N__34609\
        );

    \I__5959\ : Span4Mux_v
    port map (
            O => \N__34615\,
            I => \N__34604\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__34612\,
            I => \N__34604\
        );

    \I__5957\ : Odrv12
    port map (
            O => \N__34609\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_1
        );

    \I__5956\ : Odrv4
    port map (
            O => \N__34604\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_1
        );

    \I__5955\ : InMux
    port map (
            O => \N__34599\,
            I => \N__34594\
        );

    \I__5954\ : InMux
    port map (
            O => \N__34598\,
            I => \N__34589\
        );

    \I__5953\ : InMux
    port map (
            O => \N__34597\,
            I => \N__34589\
        );

    \I__5952\ : LocalMux
    port map (
            O => \N__34594\,
            I => \N__34584\
        );

    \I__5951\ : LocalMux
    port map (
            O => \N__34589\,
            I => \N__34584\
        );

    \I__5950\ : Span4Mux_v
    port map (
            O => \N__34584\,
            I => \N__34581\
        );

    \I__5949\ : Span4Mux_v
    port map (
            O => \N__34581\,
            I => \N__34578\
        );

    \I__5948\ : Odrv4
    port map (
            O => \N__34578\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_349\
        );

    \I__5947\ : InMux
    port map (
            O => \N__34575\,
            I => \N__34572\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__34572\,
            I => \serializer_mod_inst.shift_regZ0Z_7\
        );

    \I__5945\ : InMux
    port map (
            O => \N__34569\,
            I => \N__34566\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__34566\,
            I => \serializer_mod_inst.shift_regZ0Z_31\
        );

    \I__5943\ : InMux
    port map (
            O => \N__34563\,
            I => \N__34560\
        );

    \I__5942\ : LocalMux
    port map (
            O => \N__34560\,
            I => \serializer_mod_inst.shift_regZ0Z_32\
        );

    \I__5941\ : CascadeMux
    port map (
            O => \N__34557\,
            I => \N__34552\
        );

    \I__5940\ : InMux
    port map (
            O => \N__34556\,
            I => \N__34544\
        );

    \I__5939\ : InMux
    port map (
            O => \N__34555\,
            I => \N__34544\
        );

    \I__5938\ : InMux
    port map (
            O => \N__34552\,
            I => \N__34544\
        );

    \I__5937\ : CascadeMux
    port map (
            O => \N__34551\,
            I => \N__34540\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__34544\,
            I => \N__34537\
        );

    \I__5935\ : InMux
    port map (
            O => \N__34543\,
            I => \N__34532\
        );

    \I__5934\ : InMux
    port map (
            O => \N__34540\,
            I => \N__34532\
        );

    \I__5933\ : Span4Mux_h
    port map (
            O => \N__34537\,
            I => \N__34529\
        );

    \I__5932\ : LocalMux
    port map (
            O => \N__34532\,
            I => \N__34526\
        );

    \I__5931\ : Odrv4
    port map (
            O => \N__34529\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13\
        );

    \I__5930\ : Odrv4
    port map (
            O => \N__34526\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13\
        );

    \I__5929\ : InMux
    port map (
            O => \N__34521\,
            I => \N__34518\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__34518\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1880\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__34515\,
            I => \cemf_module_64ch_ctrl_inst1.N_1848_0_cascade_\
        );

    \I__5926\ : InMux
    port map (
            O => \N__34512\,
            I => \N__34508\
        );

    \I__5925\ : InMux
    port map (
            O => \N__34511\,
            I => \N__34505\
        );

    \I__5924\ : LocalMux
    port map (
            O => \N__34508\,
            I => \N__34502\
        );

    \I__5923\ : LocalMux
    port map (
            O => \N__34505\,
            I => \N__34497\
        );

    \I__5922\ : Span4Mux_v
    port map (
            O => \N__34502\,
            I => \N__34497\
        );

    \I__5921\ : Odrv4
    port map (
            O => \N__34497\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1884_0\
        );

    \I__5920\ : InMux
    port map (
            O => \N__34494\,
            I => \N__34491\
        );

    \I__5919\ : LocalMux
    port map (
            O => \N__34491\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0\
        );

    \I__5918\ : CascadeMux
    port map (
            O => \N__34488\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0_cascade_\
        );

    \I__5917\ : InMux
    port map (
            O => \N__34485\,
            I => \N__34482\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__34482\,
            I => \N__34479\
        );

    \I__5915\ : Odrv4
    port map (
            O => \N__34479\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392_reti\
        );

    \I__5914\ : CascadeMux
    port map (
            O => \N__34476\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0_a2_6_1_cascade_\
        );

    \I__5913\ : CascadeMux
    port map (
            O => \N__34473\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1399_cascade_\
        );

    \I__5912\ : CascadeMux
    port map (
            O => \N__34470\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0_cascade_\
        );

    \I__5911\ : CascadeMux
    port map (
            O => \N__34467\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1395_cascade_\
        );

    \I__5910\ : InMux
    port map (
            O => \N__34464\,
            I => \N__34461\
        );

    \I__5909\ : LocalMux
    port map (
            O => \N__34461\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_0_10\
        );

    \I__5908\ : CascadeMux
    port map (
            O => \N__34458\,
            I => \N__34450\
        );

    \I__5907\ : InMux
    port map (
            O => \N__34457\,
            I => \N__34442\
        );

    \I__5906\ : InMux
    port map (
            O => \N__34456\,
            I => \N__34442\
        );

    \I__5905\ : InMux
    port map (
            O => \N__34455\,
            I => \N__34442\
        );

    \I__5904\ : InMux
    port map (
            O => \N__34454\,
            I => \N__34433\
        );

    \I__5903\ : InMux
    port map (
            O => \N__34453\,
            I => \N__34433\
        );

    \I__5902\ : InMux
    port map (
            O => \N__34450\,
            I => \N__34433\
        );

    \I__5901\ : InMux
    port map (
            O => \N__34449\,
            I => \N__34433\
        );

    \I__5900\ : LocalMux
    port map (
            O => \N__34442\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__34433\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10\
        );

    \I__5898\ : InMux
    port map (
            O => \N__34428\,
            I => \N__34425\
        );

    \I__5897\ : LocalMux
    port map (
            O => \N__34425\,
            I => \N__34422\
        );

    \I__5896\ : Span4Mux_v
    port map (
            O => \N__34422\,
            I => \N__34417\
        );

    \I__5895\ : InMux
    port map (
            O => \N__34421\,
            I => \N__34414\
        );

    \I__5894\ : InMux
    port map (
            O => \N__34420\,
            I => \N__34411\
        );

    \I__5893\ : Odrv4
    port map (
            O => \N__34417\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__34414\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8\
        );

    \I__5891\ : LocalMux
    port map (
            O => \N__34411\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8\
        );

    \I__5890\ : InMux
    port map (
            O => \N__34404\,
            I => \N__34400\
        );

    \I__5889\ : InMux
    port map (
            O => \N__34403\,
            I => \N__34397\
        );

    \I__5888\ : LocalMux
    port map (
            O => \N__34400\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__34397\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0\
        );

    \I__5886\ : InMux
    port map (
            O => \N__34392\,
            I => \N__34389\
        );

    \I__5885\ : LocalMux
    port map (
            O => \N__34389\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_14\
        );

    \I__5884\ : CascadeMux
    port map (
            O => \N__34386\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1409_cascade_\
        );

    \I__5883\ : InMux
    port map (
            O => \N__34383\,
            I => \N__34376\
        );

    \I__5882\ : InMux
    port map (
            O => \N__34382\,
            I => \N__34376\
        );

    \I__5881\ : InMux
    port map (
            O => \N__34381\,
            I => \N__34372\
        );

    \I__5880\ : LocalMux
    port map (
            O => \N__34376\,
            I => \N__34369\
        );

    \I__5879\ : InMux
    port map (
            O => \N__34375\,
            I => \N__34366\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__34372\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1372_0\
        );

    \I__5877\ : Odrv4
    port map (
            O => \N__34369\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1372_0\
        );

    \I__5876\ : LocalMux
    port map (
            O => \N__34366\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1372_0\
        );

    \I__5875\ : InMux
    port map (
            O => \N__34359\,
            I => \N__34355\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__34358\,
            I => \N__34351\
        );

    \I__5873\ : LocalMux
    port map (
            O => \N__34355\,
            I => \N__34348\
        );

    \I__5872\ : InMux
    port map (
            O => \N__34354\,
            I => \N__34343\
        );

    \I__5871\ : InMux
    port map (
            O => \N__34351\,
            I => \N__34343\
        );

    \I__5870\ : Span4Mux_h
    port map (
            O => \N__34348\,
            I => \N__34340\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__34343\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14\
        );

    \I__5868\ : Odrv4
    port map (
            O => \N__34340\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14\
        );

    \I__5867\ : InMux
    port map (
            O => \N__34335\,
            I => \N__34317\
        );

    \I__5866\ : InMux
    port map (
            O => \N__34334\,
            I => \N__34317\
        );

    \I__5865\ : InMux
    port map (
            O => \N__34333\,
            I => \N__34317\
        );

    \I__5864\ : InMux
    port map (
            O => \N__34332\,
            I => \N__34317\
        );

    \I__5863\ : InMux
    port map (
            O => \N__34331\,
            I => \N__34317\
        );

    \I__5862\ : InMux
    port map (
            O => \N__34330\,
            I => \N__34317\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__34317\,
            I => \N__34314\
        );

    \I__5860\ : Span4Mux_v
    port map (
            O => \N__34314\,
            I => \N__34310\
        );

    \I__5859\ : InMux
    port map (
            O => \N__34313\,
            I => \N__34307\
        );

    \I__5858\ : Odrv4
    port map (
            O => \N__34310\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1379_0\
        );

    \I__5857\ : LocalMux
    port map (
            O => \N__34307\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1379_0\
        );

    \I__5856\ : CascadeMux
    port map (
            O => \N__34302\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1400_cascade_\
        );

    \I__5855\ : InMux
    port map (
            O => \N__34299\,
            I => \N__34296\
        );

    \I__5854\ : LocalMux
    port map (
            O => \N__34296\,
            I => \N__34292\
        );

    \I__5853\ : InMux
    port map (
            O => \N__34295\,
            I => \N__34289\
        );

    \I__5852\ : Span4Mux_v
    port map (
            O => \N__34292\,
            I => \N__34286\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__34289\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1374_0\
        );

    \I__5850\ : Odrv4
    port map (
            O => \N__34286\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1374_0\
        );

    \I__5849\ : InMux
    port map (
            O => \N__34281\,
            I => \N__34277\
        );

    \I__5848\ : InMux
    port map (
            O => \N__34280\,
            I => \N__34273\
        );

    \I__5847\ : LocalMux
    port map (
            O => \N__34277\,
            I => \N__34269\
        );

    \I__5846\ : InMux
    port map (
            O => \N__34276\,
            I => \N__34266\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__34273\,
            I => \N__34263\
        );

    \I__5844\ : InMux
    port map (
            O => \N__34272\,
            I => \N__34260\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__34269\,
            I => \N__34257\
        );

    \I__5842\ : LocalMux
    port map (
            O => \N__34266\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0\
        );

    \I__5841\ : Odrv12
    port map (
            O => \N__34263\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0\
        );

    \I__5840\ : LocalMux
    port map (
            O => \N__34260\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0\
        );

    \I__5839\ : Odrv4
    port map (
            O => \N__34257\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0\
        );

    \I__5838\ : InMux
    port map (
            O => \N__34248\,
            I => \N__34245\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__34245\,
            I => \N__34241\
        );

    \I__5836\ : InMux
    port map (
            O => \N__34244\,
            I => \N__34237\
        );

    \I__5835\ : Span4Mux_h
    port map (
            O => \N__34241\,
            I => \N__34234\
        );

    \I__5834\ : InMux
    port map (
            O => \N__34240\,
            I => \N__34231\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__34237\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__34234\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2\
        );

    \I__5831\ : LocalMux
    port map (
            O => \N__34231\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2\
        );

    \I__5830\ : CascadeMux
    port map (
            O => \N__34224\,
            I => \N__34221\
        );

    \I__5829\ : InMux
    port map (
            O => \N__34221\,
            I => \N__34218\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__34218\,
            I => \N__34213\
        );

    \I__5827\ : InMux
    port map (
            O => \N__34217\,
            I => \N__34210\
        );

    \I__5826\ : InMux
    port map (
            O => \N__34216\,
            I => \N__34207\
        );

    \I__5825\ : Span4Mux_h
    port map (
            O => \N__34213\,
            I => \N__34204\
        );

    \I__5824\ : LocalMux
    port map (
            O => \N__34210\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3\
        );

    \I__5823\ : LocalMux
    port map (
            O => \N__34207\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3\
        );

    \I__5822\ : Odrv4
    port map (
            O => \N__34204\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3\
        );

    \I__5821\ : InMux
    port map (
            O => \N__34197\,
            I => \N__34194\
        );

    \I__5820\ : LocalMux
    port map (
            O => \N__34194\,
            I => \N__34191\
        );

    \I__5819\ : Span4Mux_h
    port map (
            O => \N__34191\,
            I => \N__34186\
        );

    \I__5818\ : InMux
    port map (
            O => \N__34190\,
            I => \N__34183\
        );

    \I__5817\ : InMux
    port map (
            O => \N__34189\,
            I => \N__34180\
        );

    \I__5816\ : Odrv4
    port map (
            O => \N__34186\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__34183\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1\
        );

    \I__5814\ : LocalMux
    port map (
            O => \N__34180\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1\
        );

    \I__5813\ : CascadeMux
    port map (
            O => \N__34173\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0_cascade_\
        );

    \I__5812\ : InMux
    port map (
            O => \N__34170\,
            I => \N__34163\
        );

    \I__5811\ : InMux
    port map (
            O => \N__34169\,
            I => \N__34154\
        );

    \I__5810\ : InMux
    port map (
            O => \N__34168\,
            I => \N__34154\
        );

    \I__5809\ : InMux
    port map (
            O => \N__34167\,
            I => \N__34154\
        );

    \I__5808\ : InMux
    port map (
            O => \N__34166\,
            I => \N__34154\
        );

    \I__5807\ : LocalMux
    port map (
            O => \N__34163\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6\
        );

    \I__5806\ : LocalMux
    port map (
            O => \N__34154\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6\
        );

    \I__5805\ : CascadeMux
    port map (
            O => \N__34149\,
            I => \N__34143\
        );

    \I__5804\ : InMux
    port map (
            O => \N__34148\,
            I => \N__34140\
        );

    \I__5803\ : InMux
    port map (
            O => \N__34147\,
            I => \N__34137\
        );

    \I__5802\ : InMux
    port map (
            O => \N__34146\,
            I => \N__34132\
        );

    \I__5801\ : InMux
    port map (
            O => \N__34143\,
            I => \N__34132\
        );

    \I__5800\ : LocalMux
    port map (
            O => \N__34140\,
            I => \N__34129\
        );

    \I__5799\ : LocalMux
    port map (
            O => \N__34137\,
            I => \N__34126\
        );

    \I__5798\ : LocalMux
    port map (
            O => \N__34132\,
            I => \N__34122\
        );

    \I__5797\ : Span4Mux_v
    port map (
            O => \N__34129\,
            I => \N__34117\
        );

    \I__5796\ : Span4Mux_h
    port map (
            O => \N__34126\,
            I => \N__34117\
        );

    \I__5795\ : CascadeMux
    port map (
            O => \N__34125\,
            I => \N__34113\
        );

    \I__5794\ : Span4Mux_v
    port map (
            O => \N__34122\,
            I => \N__34110\
        );

    \I__5793\ : Span4Mux_v
    port map (
            O => \N__34117\,
            I => \N__34107\
        );

    \I__5792\ : InMux
    port map (
            O => \N__34116\,
            I => \N__34102\
        );

    \I__5791\ : InMux
    port map (
            O => \N__34113\,
            I => \N__34102\
        );

    \I__5790\ : Span4Mux_v
    port map (
            O => \N__34110\,
            I => \N__34099\
        );

    \I__5789\ : Odrv4
    port map (
            O => \N__34107\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1\
        );

    \I__5788\ : LocalMux
    port map (
            O => \N__34102\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1\
        );

    \I__5787\ : Odrv4
    port map (
            O => \N__34099\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1\
        );

    \I__5786\ : InMux
    port map (
            O => \N__34092\,
            I => \N__34086\
        );

    \I__5785\ : InMux
    port map (
            O => \N__34091\,
            I => \N__34086\
        );

    \I__5784\ : LocalMux
    port map (
            O => \N__34086\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_1786_2\
        );

    \I__5783\ : InMux
    port map (
            O => \N__34083\,
            I => \N__34080\
        );

    \I__5782\ : LocalMux
    port map (
            O => \N__34080\,
            I => \N__34077\
        );

    \I__5781\ : Odrv4
    port map (
            O => \N__34077\,
            I => \N_979\
        );

    \I__5780\ : InMux
    port map (
            O => \N__34074\,
            I => \N__34071\
        );

    \I__5779\ : LocalMux
    port map (
            O => \N__34071\,
            I => \N__34068\
        );

    \I__5778\ : Span4Mux_h
    port map (
            O => \N__34068\,
            I => \N__34065\
        );

    \I__5777\ : Odrv4
    port map (
            O => \N__34065\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_id_prdata_1_4_u_i_0\
        );

    \I__5776\ : InMux
    port map (
            O => \N__34062\,
            I => \N__34059\
        );

    \I__5775\ : LocalMux
    port map (
            O => \N__34059\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2
        );

    \I__5774\ : CascadeMux
    port map (
            O => \N__34056\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2_cascade_\
        );

    \I__5773\ : CascadeMux
    port map (
            O => \N__34053\,
            I => \N_1838_0_cascade_\
        );

    \I__5772\ : InMux
    port map (
            O => \N__34050\,
            I => \N__34046\
        );

    \I__5771\ : InMux
    port map (
            O => \N__34049\,
            I => \N__34043\
        );

    \I__5770\ : LocalMux
    port map (
            O => \N__34046\,
            I => \N__34040\
        );

    \I__5769\ : LocalMux
    port map (
            O => \N__34043\,
            I => \N__34037\
        );

    \I__5768\ : Span4Mux_h
    port map (
            O => \N__34040\,
            I => \N__34034\
        );

    \I__5767\ : Span4Mux_h
    port map (
            O => \N__34037\,
            I => \N__34031\
        );

    \I__5766\ : Odrv4
    port map (
            O => \N__34034\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable
        );

    \I__5765\ : Odrv4
    port map (
            O => \N__34031\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable
        );

    \I__5764\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34023\
        );

    \I__5763\ : LocalMux
    port map (
            O => \N__34023\,
            I => \N__34020\
        );

    \I__5762\ : Span4Mux_v
    port map (
            O => \N__34020\,
            I => \N__34017\
        );

    \I__5761\ : Span4Mux_h
    port map (
            O => \N__34017\,
            I => \N__34014\
        );

    \I__5760\ : Odrv4
    port map (
            O => \N__34014\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_30\
        );

    \I__5759\ : CascadeMux
    port map (
            O => \N__34011\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1654_cascade_\
        );

    \I__5758\ : CascadeMux
    port map (
            O => \N__34008\,
            I => \N_12_0_cascade_\
        );

    \I__5757\ : InMux
    port map (
            O => \N__34005\,
            I => \N__34002\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__34002\,
            I => \N__33998\
        );

    \I__5755\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33995\
        );

    \I__5754\ : Span4Mux_h
    port map (
            O => \N__33998\,
            I => \N__33991\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__33995\,
            I => \N__33988\
        );

    \I__5752\ : InMux
    port map (
            O => \N__33994\,
            I => \N__33985\
        );

    \I__5751\ : Span4Mux_v
    port map (
            O => \N__33991\,
            I => \N__33980\
        );

    \I__5750\ : Span4Mux_h
    port map (
            O => \N__33988\,
            I => \N__33980\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__33985\,
            I => \N__33977\
        );

    \I__5748\ : Span4Mux_v
    port map (
            O => \N__33980\,
            I => \N__33971\
        );

    \I__5747\ : Span4Mux_h
    port map (
            O => \N__33977\,
            I => \N__33971\
        );

    \I__5746\ : InMux
    port map (
            O => \N__33976\,
            I => \N__33968\
        );

    \I__5745\ : Span4Mux_v
    port map (
            O => \N__33971\,
            I => \N__33965\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__33968\,
            I => \N__33962\
        );

    \I__5743\ : Span4Mux_h
    port map (
            O => \N__33965\,
            I => \N__33959\
        );

    \I__5742\ : Span12Mux_h
    port map (
            O => \N__33962\,
            I => \N__33956\
        );

    \I__5741\ : Odrv4
    port map (
            O => \N__33959\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7\
        );

    \I__5740\ : Odrv12
    port map (
            O => \N__33956\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7\
        );

    \I__5739\ : InMux
    port map (
            O => \N__33951\,
            I => \N__33926\
        );

    \I__5738\ : CascadeMux
    port map (
            O => \N__33950\,
            I => \N__33923\
        );

    \I__5737\ : InMux
    port map (
            O => \N__33949\,
            I => \N__33901\
        );

    \I__5736\ : InMux
    port map (
            O => \N__33948\,
            I => \N__33901\
        );

    \I__5735\ : InMux
    port map (
            O => \N__33947\,
            I => \N__33901\
        );

    \I__5734\ : InMux
    port map (
            O => \N__33946\,
            I => \N__33901\
        );

    \I__5733\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33901\
        );

    \I__5732\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33901\
        );

    \I__5731\ : InMux
    port map (
            O => \N__33943\,
            I => \N__33901\
        );

    \I__5730\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33886\
        );

    \I__5729\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33886\
        );

    \I__5728\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33886\
        );

    \I__5727\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33886\
        );

    \I__5726\ : InMux
    port map (
            O => \N__33938\,
            I => \N__33886\
        );

    \I__5725\ : InMux
    port map (
            O => \N__33937\,
            I => \N__33886\
        );

    \I__5724\ : InMux
    port map (
            O => \N__33936\,
            I => \N__33886\
        );

    \I__5723\ : InMux
    port map (
            O => \N__33935\,
            I => \N__33871\
        );

    \I__5722\ : InMux
    port map (
            O => \N__33934\,
            I => \N__33871\
        );

    \I__5721\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33871\
        );

    \I__5720\ : InMux
    port map (
            O => \N__33932\,
            I => \N__33871\
        );

    \I__5719\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33871\
        );

    \I__5718\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33871\
        );

    \I__5717\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33871\
        );

    \I__5716\ : LocalMux
    port map (
            O => \N__33926\,
            I => \N__33868\
        );

    \I__5715\ : InMux
    port map (
            O => \N__33923\,
            I => \N__33865\
        );

    \I__5714\ : InMux
    port map (
            O => \N__33922\,
            I => \N__33862\
        );

    \I__5713\ : InMux
    port map (
            O => \N__33921\,
            I => \N__33849\
        );

    \I__5712\ : InMux
    port map (
            O => \N__33920\,
            I => \N__33849\
        );

    \I__5711\ : InMux
    port map (
            O => \N__33919\,
            I => \N__33849\
        );

    \I__5710\ : InMux
    port map (
            O => \N__33918\,
            I => \N__33849\
        );

    \I__5709\ : InMux
    port map (
            O => \N__33917\,
            I => \N__33849\
        );

    \I__5708\ : InMux
    port map (
            O => \N__33916\,
            I => \N__33849\
        );

    \I__5707\ : LocalMux
    port map (
            O => \N__33901\,
            I => \N__33846\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__33886\,
            I => \N__33841\
        );

    \I__5705\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33841\
        );

    \I__5704\ : Span12Mux_h
    port map (
            O => \N__33868\,
            I => \N__33838\
        );

    \I__5703\ : LocalMux
    port map (
            O => \N__33865\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__33862\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__33849\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\
        );

    \I__5700\ : Odrv4
    port map (
            O => \N__33846\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\
        );

    \I__5699\ : Odrv12
    port map (
            O => \N__33841\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\
        );

    \I__5698\ : Odrv12
    port map (
            O => \N__33838\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\
        );

    \I__5697\ : InMux
    port map (
            O => \N__33825\,
            I => \N__33822\
        );

    \I__5696\ : LocalMux
    port map (
            O => \N__33822\,
            I => \N__33818\
        );

    \I__5695\ : InMux
    port map (
            O => \N__33821\,
            I => \N__33815\
        );

    \I__5694\ : Span4Mux_v
    port map (
            O => \N__33818\,
            I => \N__33812\
        );

    \I__5693\ : LocalMux
    port map (
            O => \N__33815\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_7
        );

    \I__5692\ : Odrv4
    port map (
            O => \N__33812\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_7
        );

    \I__5691\ : CascadeMux
    port map (
            O => \N__33807\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0_cascade_\
        );

    \I__5690\ : InMux
    port map (
            O => \N__33804\,
            I => \N__33801\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__33801\,
            I => \N_12_0\
        );

    \I__5688\ : InMux
    port map (
            O => \N__33798\,
            I => \N__33795\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__33795\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_0_7\
        );

    \I__5686\ : CascadeMux
    port map (
            O => \N__33792\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_23_cascade_\
        );

    \I__5685\ : CascadeMux
    port map (
            O => \N__33789\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDDZ0Z7_cascade_\
        );

    \I__5684\ : CascadeMux
    port map (
            O => \N__33786\,
            I => \N__33783\
        );

    \I__5683\ : InMux
    port map (
            O => \N__33783\,
            I => \N__33780\
        );

    \I__5682\ : LocalMux
    port map (
            O => \N__33780\,
            I => \N__33776\
        );

    \I__5681\ : InMux
    port map (
            O => \N__33779\,
            I => \N__33772\
        );

    \I__5680\ : Span4Mux_h
    port map (
            O => \N__33776\,
            I => \N__33769\
        );

    \I__5679\ : InMux
    port map (
            O => \N__33775\,
            I => \N__33766\
        );

    \I__5678\ : LocalMux
    port map (
            O => \N__33772\,
            I => \N__33761\
        );

    \I__5677\ : Span4Mux_h
    port map (
            O => \N__33769\,
            I => \N__33761\
        );

    \I__5676\ : LocalMux
    port map (
            O => \N__33766\,
            I => \N__33758\
        );

    \I__5675\ : Span4Mux_v
    port map (
            O => \N__33761\,
            I => \N__33755\
        );

    \I__5674\ : Span12Mux_h
    port map (
            O => \N__33758\,
            I => \N__33752\
        );

    \I__5673\ : Odrv4
    port map (
            O => \N__33755\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_6
        );

    \I__5672\ : Odrv12
    port map (
            O => \N__33752\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_6
        );

    \I__5671\ : InMux
    port map (
            O => \N__33747\,
            I => \N__33744\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__33744\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_6\
        );

    \I__5669\ : InMux
    port map (
            O => \N__33741\,
            I => \N__33738\
        );

    \I__5668\ : LocalMux
    port map (
            O => \N__33738\,
            I => \N__33734\
        );

    \I__5667\ : CascadeMux
    port map (
            O => \N__33737\,
            I => \N__33731\
        );

    \I__5666\ : Span4Mux_h
    port map (
            O => \N__33734\,
            I => \N__33727\
        );

    \I__5665\ : InMux
    port map (
            O => \N__33731\,
            I => \N__33722\
        );

    \I__5664\ : InMux
    port map (
            O => \N__33730\,
            I => \N__33722\
        );

    \I__5663\ : Span4Mux_v
    port map (
            O => \N__33727\,
            I => \N__33717\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__33722\,
            I => \N__33717\
        );

    \I__5661\ : Odrv4
    port map (
            O => \N__33717\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_3
        );

    \I__5660\ : CascadeMux
    port map (
            O => \N__33714\,
            I => \N__33711\
        );

    \I__5659\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33707\
        );

    \I__5658\ : InMux
    port map (
            O => \N__33710\,
            I => \N__33704\
        );

    \I__5657\ : LocalMux
    port map (
            O => \N__33707\,
            I => \N__33700\
        );

    \I__5656\ : LocalMux
    port map (
            O => \N__33704\,
            I => \N__33697\
        );

    \I__5655\ : InMux
    port map (
            O => \N__33703\,
            I => \N__33694\
        );

    \I__5654\ : Span4Mux_v
    port map (
            O => \N__33700\,
            I => \N__33691\
        );

    \I__5653\ : Span4Mux_h
    port map (
            O => \N__33697\,
            I => \N__33688\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33683\
        );

    \I__5651\ : Sp12to4
    port map (
            O => \N__33691\,
            I => \N__33683\
        );

    \I__5650\ : Odrv4
    port map (
            O => \N__33688\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_4
        );

    \I__5649\ : Odrv12
    port map (
            O => \N__33683\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_4
        );

    \I__5648\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33675\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__33675\,
            I => \N__33670\
        );

    \I__5646\ : InMux
    port map (
            O => \N__33674\,
            I => \N__33665\
        );

    \I__5645\ : InMux
    port map (
            O => \N__33673\,
            I => \N__33665\
        );

    \I__5644\ : Span4Mux_h
    port map (
            O => \N__33670\,
            I => \N__33662\
        );

    \I__5643\ : LocalMux
    port map (
            O => \N__33665\,
            I => \N__33659\
        );

    \I__5642\ : Odrv4
    port map (
            O => \N__33662\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_6
        );

    \I__5641\ : Odrv4
    port map (
            O => \N__33659\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_6
        );

    \I__5640\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33651\
        );

    \I__5639\ : LocalMux
    port map (
            O => \N__33651\,
            I => \N__33648\
        );

    \I__5638\ : Span4Mux_h
    port map (
            O => \N__33648\,
            I => \N__33645\
        );

    \I__5637\ : Span4Mux_h
    port map (
            O => \N__33645\,
            I => \N__33642\
        );

    \I__5636\ : Odrv4
    port map (
            O => \N__33642\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_0Z0Z_26\
        );

    \I__5635\ : CascadeMux
    port map (
            O => \N__33639\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGHZ0Z5_cascade_\
        );

    \I__5634\ : InMux
    port map (
            O => \N__33636\,
            I => \N__33630\
        );

    \I__5633\ : InMux
    port map (
            O => \N__33635\,
            I => \N__33630\
        );

    \I__5632\ : LocalMux
    port map (
            O => \N__33630\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_15\
        );

    \I__5631\ : InMux
    port map (
            O => \N__33627\,
            I => \N__33624\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__33624\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14\
        );

    \I__5629\ : InMux
    port map (
            O => \N__33621\,
            I => \N__33618\
        );

    \I__5628\ : LocalMux
    port map (
            O => \N__33618\,
            I => \N__33615\
        );

    \I__5627\ : Span4Mux_h
    port map (
            O => \N__33615\,
            I => \N__33612\
        );

    \I__5626\ : Sp12to4
    port map (
            O => \N__33612\,
            I => \N__33609\
        );

    \I__5625\ : Span12Mux_h
    port map (
            O => \N__33609\,
            I => \N__33606\
        );

    \I__5624\ : Odrv12
    port map (
            O => \N__33606\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_13\
        );

    \I__5623\ : CascadeMux
    port map (
            O => \N__33603\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14_cascade_\
        );

    \I__5622\ : CascadeMux
    port map (
            O => \N__33600\,
            I => \N__33597\
        );

    \I__5621\ : InMux
    port map (
            O => \N__33597\,
            I => \N__33594\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__33594\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_14\
        );

    \I__5619\ : CascadeMux
    port map (
            O => \N__33591\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_14_cascade_\
        );

    \I__5618\ : InMux
    port map (
            O => \N__33588\,
            I => \N__33585\
        );

    \I__5617\ : LocalMux
    port map (
            O => \N__33585\,
            I => \N__33582\
        );

    \I__5616\ : Odrv4
    port map (
            O => \N__33582\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_14\
        );

    \I__5615\ : InMux
    port map (
            O => \N__33579\,
            I => \N__33576\
        );

    \I__5614\ : LocalMux
    port map (
            O => \N__33576\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGHZ0Z5\
        );

    \I__5613\ : CascadeMux
    port map (
            O => \N__33573\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_14_cascade_\
        );

    \I__5612\ : InMux
    port map (
            O => \N__33570\,
            I => \N__33567\
        );

    \I__5611\ : LocalMux
    port map (
            O => \N__33567\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_14\
        );

    \I__5610\ : InMux
    port map (
            O => \N__33564\,
            I => \N__33561\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__33561\,
            I => \N__33558\
        );

    \I__5608\ : Span4Mux_v
    port map (
            O => \N__33558\,
            I => \N__33553\
        );

    \I__5607\ : InMux
    port map (
            O => \N__33557\,
            I => \N__33550\
        );

    \I__5606\ : InMux
    port map (
            O => \N__33556\,
            I => \N__33547\
        );

    \I__5605\ : Odrv4
    port map (
            O => \N__33553\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_14
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__33550\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_14
        );

    \I__5603\ : LocalMux
    port map (
            O => \N__33547\,
            I => cemf_module_64ch_ctrl_inst1_data_coarseovf_14
        );

    \I__5602\ : InMux
    port map (
            O => \N__33540\,
            I => \N__33537\
        );

    \I__5601\ : LocalMux
    port map (
            O => \N__33537\,
            I => \N__33534\
        );

    \I__5600\ : Span4Mux_v
    port map (
            O => \N__33534\,
            I => \N__33531\
        );

    \I__5599\ : Span4Mux_h
    port map (
            O => \N__33531\,
            I => \N__33528\
        );

    \I__5598\ : Odrv4
    port map (
            O => \N__33528\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_1\
        );

    \I__5597\ : InMux
    port map (
            O => \N__33525\,
            I => \N__33522\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__33522\,
            I => \N__33518\
        );

    \I__5595\ : CascadeMux
    port map (
            O => \N__33521\,
            I => \N__33515\
        );

    \I__5594\ : Span4Mux_v
    port map (
            O => \N__33518\,
            I => \N__33512\
        );

    \I__5593\ : InMux
    port map (
            O => \N__33515\,
            I => \N__33509\
        );

    \I__5592\ : Span4Mux_h
    port map (
            O => \N__33512\,
            I => \N__33506\
        );

    \I__5591\ : LocalMux
    port map (
            O => \N__33509\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_18
        );

    \I__5590\ : Odrv4
    port map (
            O => \N__33506\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_18
        );

    \I__5589\ : CascadeMux
    port map (
            O => \N__33501\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0_cascade_\
        );

    \I__5588\ : InMux
    port map (
            O => \N__33498\,
            I => \N__33495\
        );

    \I__5587\ : LocalMux
    port map (
            O => \N__33495\,
            I => \N__33492\
        );

    \I__5586\ : Span4Mux_h
    port map (
            O => \N__33492\,
            I => \N__33489\
        );

    \I__5585\ : Odrv4
    port map (
            O => \N__33489\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_18\
        );

    \I__5584\ : CascadeMux
    port map (
            O => \N__33486\,
            I => \N__33483\
        );

    \I__5583\ : InMux
    port map (
            O => \N__33483\,
            I => \N__33480\
        );

    \I__5582\ : LocalMux
    port map (
            O => \N__33480\,
            I => \N__33476\
        );

    \I__5581\ : InMux
    port map (
            O => \N__33479\,
            I => \N__33473\
        );

    \I__5580\ : Span4Mux_v
    port map (
            O => \N__33476\,
            I => \N__33470\
        );

    \I__5579\ : LocalMux
    port map (
            O => \N__33473\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_20
        );

    \I__5578\ : Odrv4
    port map (
            O => \N__33470\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_20
        );

    \I__5577\ : InMux
    port map (
            O => \N__33465\,
            I => \N__33462\
        );

    \I__5576\ : LocalMux
    port map (
            O => \N__33462\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_20\
        );

    \I__5575\ : CascadeMux
    port map (
            O => \N__33459\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0_cascade_\
        );

    \I__5574\ : InMux
    port map (
            O => \N__33456\,
            I => \N__33453\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33450\
        );

    \I__5572\ : Span4Mux_v
    port map (
            O => \N__33450\,
            I => \N__33447\
        );

    \I__5571\ : Sp12to4
    port map (
            O => \N__33447\,
            I => \N__33444\
        );

    \I__5570\ : Odrv12
    port map (
            O => \N__33444\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_7\
        );

    \I__5569\ : CascadeMux
    port map (
            O => \N__33441\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_15_cascade_\
        );

    \I__5568\ : InMux
    port map (
            O => \N__33438\,
            I => \N__33435\
        );

    \I__5567\ : LocalMux
    port map (
            O => \N__33435\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_19\
        );

    \I__5566\ : InMux
    port map (
            O => \N__33432\,
            I => \N__33428\
        );

    \I__5565\ : InMux
    port map (
            O => \N__33431\,
            I => \N__33425\
        );

    \I__5564\ : LocalMux
    port map (
            O => \N__33428\,
            I => \N__33422\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__33425\,
            I => \N__33419\
        );

    \I__5562\ : Span12Mux_v
    port map (
            O => \N__33422\,
            I => \N__33416\
        );

    \I__5561\ : Span12Mux_v
    port map (
            O => \N__33419\,
            I => \N__33413\
        );

    \I__5560\ : Odrv12
    port map (
            O => \N__33416\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable
        );

    \I__5559\ : Odrv12
    port map (
            O => \N__33413\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable
        );

    \I__5558\ : InMux
    port map (
            O => \N__33408\,
            I => \N__33405\
        );

    \I__5557\ : LocalMux
    port map (
            O => \N__33405\,
            I => \N__33402\
        );

    \I__5556\ : Span4Mux_v
    port map (
            O => \N__33402\,
            I => \N__33399\
        );

    \I__5555\ : Sp12to4
    port map (
            O => \N__33399\,
            I => \N__33396\
        );

    \I__5554\ : Odrv12
    port map (
            O => \N__33396\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_0
        );

    \I__5553\ : InMux
    port map (
            O => \N__33393\,
            I => \N__33390\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__33390\,
            I => \N__33387\
        );

    \I__5551\ : Span4Mux_v
    port map (
            O => \N__33387\,
            I => \N__33384\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__33384\,
            I => \N__33381\
        );

    \I__5549\ : Sp12to4
    port map (
            O => \N__33381\,
            I => \N__33378\
        );

    \I__5548\ : Odrv12
    port map (
            O => \N__33378\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_0
        );

    \I__5547\ : CascadeMux
    port map (
            O => \N__33375\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319_cascade_\
        );

    \I__5546\ : CascadeMux
    port map (
            O => \N__33372\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_0_cascade_\
        );

    \I__5545\ : CascadeMux
    port map (
            O => \N__33369\,
            I => \N__33366\
        );

    \I__5544\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33362\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__33365\,
            I => \N__33359\
        );

    \I__5542\ : LocalMux
    port map (
            O => \N__33362\,
            I => \N__33356\
        );

    \I__5541\ : InMux
    port map (
            O => \N__33359\,
            I => \N__33353\
        );

    \I__5540\ : Span4Mux_h
    port map (
            O => \N__33356\,
            I => \N__33350\
        );

    \I__5539\ : LocalMux
    port map (
            O => \N__33353\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_21
        );

    \I__5538\ : Odrv4
    port map (
            O => \N__33350\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_21
        );

    \I__5537\ : CascadeMux
    port map (
            O => \N__33345\,
            I => \N__33342\
        );

    \I__5536\ : InMux
    port map (
            O => \N__33342\,
            I => \N__33339\
        );

    \I__5535\ : LocalMux
    port map (
            O => \N__33339\,
            I => \N__33336\
        );

    \I__5534\ : Span4Mux_h
    port map (
            O => \N__33336\,
            I => \N__33333\
        );

    \I__5533\ : Span4Mux_v
    port map (
            O => \N__33333\,
            I => \N__33330\
        );

    \I__5532\ : Span4Mux_h
    port map (
            O => \N__33330\,
            I => \N__33327\
        );

    \I__5531\ : Odrv4
    port map (
            O => \N__33327\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_22
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__33324\,
            I => \N__33321\
        );

    \I__5529\ : InMux
    port map (
            O => \N__33321\,
            I => \N__33318\
        );

    \I__5528\ : LocalMux
    port map (
            O => \N__33318\,
            I => \N__33315\
        );

    \I__5527\ : Odrv4
    port map (
            O => \N__33315\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_698\
        );

    \I__5526\ : InMux
    port map (
            O => \N__33312\,
            I => \N__33309\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__33309\,
            I => \N__33306\
        );

    \I__5524\ : Sp12to4
    port map (
            O => \N__33306\,
            I => \N__33303\
        );

    \I__5523\ : Span12Mux_s11_v
    port map (
            O => \N__33303\,
            I => \N__33300\
        );

    \I__5522\ : Odrv12
    port map (
            O => \N__33300\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_23
        );

    \I__5521\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33294\
        );

    \I__5520\ : LocalMux
    port map (
            O => \N__33294\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_2\
        );

    \I__5519\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33288\
        );

    \I__5518\ : LocalMux
    port map (
            O => \N__33288\,
            I => \N__33285\
        );

    \I__5517\ : Span4Mux_h
    port map (
            O => \N__33285\,
            I => \N__33282\
        );

    \I__5516\ : Span4Mux_h
    port map (
            O => \N__33282\,
            I => \N__33279\
        );

    \I__5515\ : Span4Mux_h
    port map (
            O => \N__33279\,
            I => \N__33276\
        );

    \I__5514\ : Odrv4
    port map (
            O => \N__33276\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_25
        );

    \I__5513\ : CascadeMux
    port map (
            O => \N__33273\,
            I => \N__33270\
        );

    \I__5512\ : InMux
    port map (
            O => \N__33270\,
            I => \N__33267\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__33267\,
            I => \N__33264\
        );

    \I__5510\ : Span4Mux_v
    port map (
            O => \N__33264\,
            I => \N__33261\
        );

    \I__5509\ : Span4Mux_h
    port map (
            O => \N__33261\,
            I => \N__33258\
        );

    \I__5508\ : Odrv4
    port map (
            O => \N__33258\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_27
        );

    \I__5507\ : InMux
    port map (
            O => \N__33255\,
            I => \N__33252\
        );

    \I__5506\ : LocalMux
    port map (
            O => \N__33252\,
            I => \N__33249\
        );

    \I__5505\ : Span4Mux_v
    port map (
            O => \N__33249\,
            I => \N__33246\
        );

    \I__5504\ : Span4Mux_h
    port map (
            O => \N__33246\,
            I => \N__33243\
        );

    \I__5503\ : Span4Mux_h
    port map (
            O => \N__33243\,
            I => \N__33240\
        );

    \I__5502\ : Odrv4
    port map (
            O => \N__33240\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_19
        );

    \I__5501\ : CascadeMux
    port map (
            O => \N__33237\,
            I => \N__33234\
        );

    \I__5500\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33231\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__33231\,
            I => \N__33228\
        );

    \I__5498\ : Span4Mux_v
    port map (
            O => \N__33228\,
            I => \N__33225\
        );

    \I__5497\ : Span4Mux_h
    port map (
            O => \N__33225\,
            I => \N__33222\
        );

    \I__5496\ : Span4Mux_h
    port map (
            O => \N__33222\,
            I => \N__33219\
        );

    \I__5495\ : Odrv4
    port map (
            O => \N__33219\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_19
        );

    \I__5494\ : InMux
    port map (
            O => \N__33216\,
            I => \N__33213\
        );

    \I__5493\ : LocalMux
    port map (
            O => \N__33213\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_731\
        );

    \I__5492\ : InMux
    port map (
            O => \N__33210\,
            I => \N__33207\
        );

    \I__5491\ : LocalMux
    port map (
            O => \N__33207\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_19\
        );

    \I__5490\ : CascadeMux
    port map (
            O => \N__33204\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_19_cascade_\
        );

    \I__5489\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33198\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__33198\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_19\
        );

    \I__5487\ : InMux
    port map (
            O => \N__33195\,
            I => \N__33192\
        );

    \I__5486\ : LocalMux
    port map (
            O => \N__33192\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_19\
        );

    \I__5485\ : InMux
    port map (
            O => \N__33189\,
            I => \N__33186\
        );

    \I__5484\ : LocalMux
    port map (
            O => \N__33186\,
            I => \serializer_mod_inst.shift_regZ0Z_37\
        );

    \I__5483\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33180\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__33180\,
            I => \serializer_mod_inst.shift_regZ0Z_38\
        );

    \I__5481\ : InMux
    port map (
            O => \N__33177\,
            I => \N__33174\
        );

    \I__5480\ : LocalMux
    port map (
            O => \N__33174\,
            I => \serializer_mod_inst.shift_regZ0Z_33\
        );

    \I__5479\ : InMux
    port map (
            O => \N__33171\,
            I => \N__33168\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__33168\,
            I => \serializer_mod_inst.shift_regZ0Z_34\
        );

    \I__5477\ : InMux
    port map (
            O => \N__33165\,
            I => \N__33162\
        );

    \I__5476\ : LocalMux
    port map (
            O => \N__33162\,
            I => \serializer_mod_inst.shift_regZ0Z_35\
        );

    \I__5475\ : InMux
    port map (
            O => \N__33159\,
            I => \N__33156\
        );

    \I__5474\ : LocalMux
    port map (
            O => \N__33156\,
            I => \serializer_mod_inst.shift_regZ0Z_76\
        );

    \I__5473\ : InMux
    port map (
            O => \N__33153\,
            I => \N__33150\
        );

    \I__5472\ : LocalMux
    port map (
            O => \N__33150\,
            I => \N__33147\
        );

    \I__5471\ : Span4Mux_h
    port map (
            O => \N__33147\,
            I => \N__33144\
        );

    \I__5470\ : Span4Mux_v
    port map (
            O => \N__33144\,
            I => \N__33141\
        );

    \I__5469\ : Sp12to4
    port map (
            O => \N__33141\,
            I => \N__33138\
        );

    \I__5468\ : Odrv12
    port map (
            O => \N__33138\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_17
        );

    \I__5467\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33132\
        );

    \I__5466\ : LocalMux
    port map (
            O => \N__33132\,
            I => \N__33129\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__33129\,
            I => \N__33126\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__33126\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_753\
        );

    \I__5463\ : CascadeMux
    port map (
            O => \N__33123\,
            I => \N__33120\
        );

    \I__5462\ : InMux
    port map (
            O => \N__33120\,
            I => \N__33117\
        );

    \I__5461\ : LocalMux
    port map (
            O => \N__33117\,
            I => \N__33114\
        );

    \I__5460\ : Span4Mux_h
    port map (
            O => \N__33114\,
            I => \N__33111\
        );

    \I__5459\ : Span4Mux_v
    port map (
            O => \N__33111\,
            I => \N__33108\
        );

    \I__5458\ : Span4Mux_h
    port map (
            O => \N__33108\,
            I => \N__33105\
        );

    \I__5457\ : Odrv4
    port map (
            O => \N__33105\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_19
        );

    \I__5456\ : InMux
    port map (
            O => \N__33102\,
            I => \N__33099\
        );

    \I__5455\ : LocalMux
    port map (
            O => \N__33099\,
            I => \N__33096\
        );

    \I__5454\ : Span4Mux_v
    port map (
            O => \N__33096\,
            I => \N__33093\
        );

    \I__5453\ : Span4Mux_h
    port map (
            O => \N__33093\,
            I => \N__33090\
        );

    \I__5452\ : Odrv4
    port map (
            O => \N__33090\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_2
        );

    \I__5451\ : InMux
    port map (
            O => \N__33087\,
            I => \N__33084\
        );

    \I__5450\ : LocalMux
    port map (
            O => \N__33084\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_918\
        );

    \I__5449\ : CascadeMux
    port map (
            O => \N__33081\,
            I => \N__33078\
        );

    \I__5448\ : InMux
    port map (
            O => \N__33078\,
            I => \N__33075\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__33075\,
            I => \N__33072\
        );

    \I__5446\ : Span4Mux_v
    port map (
            O => \N__33072\,
            I => \N__33069\
        );

    \I__5445\ : Span4Mux_v
    port map (
            O => \N__33069\,
            I => \N__33066\
        );

    \I__5444\ : Span4Mux_h
    port map (
            O => \N__33066\,
            I => \N__33063\
        );

    \I__5443\ : Odrv4
    port map (
            O => \N__33063\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_4\
        );

    \I__5442\ : InMux
    port map (
            O => \N__33060\,
            I => \N__33057\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__33057\,
            I => \N__33054\
        );

    \I__5440\ : Odrv4
    port map (
            O => \N__33054\,
            I => \serializer_mod_inst.shift_regZ0Z_111\
        );

    \I__5439\ : InMux
    port map (
            O => \N__33051\,
            I => \N__33048\
        );

    \I__5438\ : LocalMux
    port map (
            O => \N__33048\,
            I => \serializer_mod_inst.shift_regZ0Z_119\
        );

    \I__5437\ : InMux
    port map (
            O => \N__33045\,
            I => \N__33042\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__33042\,
            I => \serializer_mod_inst.shift_regZ0Z_120\
        );

    \I__5435\ : InMux
    port map (
            O => \N__33039\,
            I => \N__33036\
        );

    \I__5434\ : LocalMux
    port map (
            O => \N__33036\,
            I => \serializer_mod_inst.shift_regZ0Z_36\
        );

    \I__5433\ : InMux
    port map (
            O => \N__33033\,
            I => \N__33030\
        );

    \I__5432\ : LocalMux
    port map (
            O => \N__33030\,
            I => \serializer_mod_inst.shift_regZ0Z_118\
        );

    \I__5431\ : CascadeMux
    port map (
            O => \N__33027\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_2_cascade_\
        );

    \I__5430\ : InMux
    port map (
            O => \N__33024\,
            I => \N__33021\
        );

    \I__5429\ : LocalMux
    port map (
            O => \N__33021\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1950\
        );

    \I__5428\ : CascadeMux
    port map (
            O => \N__33018\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1949_cascade_\
        );

    \I__5427\ : IoInMux
    port map (
            O => \N__33015\,
            I => \N__33012\
        );

    \I__5426\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__33009\
        );

    \I__5425\ : IoSpan4Mux
    port map (
            O => \N__33009\,
            I => \N__33006\
        );

    \I__5424\ : Sp12to4
    port map (
            O => \N__33006\,
            I => \N__33003\
        );

    \I__5423\ : Span12Mux_h
    port map (
            O => \N__33003\,
            I => \N__33000\
        );

    \I__5422\ : Odrv12
    port map (
            O => \N__33000\,
            I => stop_fpga2_c
        );

    \I__5421\ : InMux
    port map (
            O => \N__32997\,
            I => \N__32994\
        );

    \I__5420\ : LocalMux
    port map (
            O => \N__32994\,
            I => \N__32989\
        );

    \I__5419\ : InMux
    port map (
            O => \N__32993\,
            I => \N__32986\
        );

    \I__5418\ : InMux
    port map (
            O => \N__32992\,
            I => \N__32983\
        );

    \I__5417\ : Span4Mux_v
    port map (
            O => \N__32989\,
            I => \N__32977\
        );

    \I__5416\ : LocalMux
    port map (
            O => \N__32986\,
            I => \N__32977\
        );

    \I__5415\ : LocalMux
    port map (
            O => \N__32983\,
            I => \N__32974\
        );

    \I__5414\ : InMux
    port map (
            O => \N__32982\,
            I => \N__32970\
        );

    \I__5413\ : Span4Mux_h
    port map (
            O => \N__32977\,
            I => \N__32967\
        );

    \I__5412\ : Span4Mux_h
    port map (
            O => \N__32974\,
            I => \N__32964\
        );

    \I__5411\ : InMux
    port map (
            O => \N__32973\,
            I => \N__32961\
        );

    \I__5410\ : LocalMux
    port map (
            O => \N__32970\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_b\
        );

    \I__5409\ : Odrv4
    port map (
            O => \N__32967\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_b\
        );

    \I__5408\ : Odrv4
    port map (
            O => \N__32964\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_b\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__32961\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_b\
        );

    \I__5406\ : InMux
    port map (
            O => \N__32952\,
            I => \N__32946\
        );

    \I__5405\ : InMux
    port map (
            O => \N__32951\,
            I => \N__32943\
        );

    \I__5404\ : InMux
    port map (
            O => \N__32950\,
            I => \N__32938\
        );

    \I__5403\ : InMux
    port map (
            O => \N__32949\,
            I => \N__32938\
        );

    \I__5402\ : LocalMux
    port map (
            O => \N__32946\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847\
        );

    \I__5401\ : LocalMux
    port map (
            O => \N__32943\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__32938\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847\
        );

    \I__5399\ : InMux
    port map (
            O => \N__32931\,
            I => \N__32928\
        );

    \I__5398\ : LocalMux
    port map (
            O => \N__32928\,
            I => \serializer_mod_inst.shift_regZ0Z_112\
        );

    \I__5397\ : CascadeMux
    port map (
            O => \N__32925\,
            I => \N__32922\
        );

    \I__5396\ : InMux
    port map (
            O => \N__32922\,
            I => \N__32919\
        );

    \I__5395\ : LocalMux
    port map (
            O => \N__32919\,
            I => \N__32916\
        );

    \I__5394\ : Span4Mux_v
    port map (
            O => \N__32916\,
            I => \N__32913\
        );

    \I__5393\ : Span4Mux_v
    port map (
            O => \N__32913\,
            I => \N__32910\
        );

    \I__5392\ : Span4Mux_v
    port map (
            O => \N__32910\,
            I => \N__32907\
        );

    \I__5391\ : Odrv4
    port map (
            O => \N__32907\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_2\
        );

    \I__5390\ : InMux
    port map (
            O => \N__32904\,
            I => \N__32896\
        );

    \I__5389\ : InMux
    port map (
            O => \N__32903\,
            I => \N__32885\
        );

    \I__5388\ : InMux
    port map (
            O => \N__32902\,
            I => \N__32885\
        );

    \I__5387\ : InMux
    port map (
            O => \N__32901\,
            I => \N__32885\
        );

    \I__5386\ : InMux
    port map (
            O => \N__32900\,
            I => \N__32885\
        );

    \I__5385\ : InMux
    port map (
            O => \N__32899\,
            I => \N__32885\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__32896\,
            I => \N__32878\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__32885\,
            I => \N__32878\
        );

    \I__5382\ : InMux
    port map (
            O => \N__32884\,
            I => \N__32875\
        );

    \I__5381\ : InMux
    port map (
            O => \N__32883\,
            I => \N__32872\
        );

    \I__5380\ : Odrv4
    port map (
            O => \N__32878\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_a\
        );

    \I__5379\ : LocalMux
    port map (
            O => \N__32875\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_a\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__32872\,
            I => \cemf_module_64ch_ctrl_inst1.end_conf_a\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__32865\,
            I => \cemf_module_64ch_ctrl_inst1.N_1817_0_cascade_\
        );

    \I__5376\ : CascadeMux
    port map (
            O => \N__32862\,
            I => \N__32859\
        );

    \I__5375\ : InMux
    port map (
            O => \N__32859\,
            I => \N__32852\
        );

    \I__5374\ : InMux
    port map (
            O => \N__32858\,
            I => \N__32843\
        );

    \I__5373\ : InMux
    port map (
            O => \N__32857\,
            I => \N__32843\
        );

    \I__5372\ : InMux
    port map (
            O => \N__32856\,
            I => \N__32843\
        );

    \I__5371\ : InMux
    port map (
            O => \N__32855\,
            I => \N__32843\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__32852\,
            I => \cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2\
        );

    \I__5369\ : LocalMux
    port map (
            O => \N__32843\,
            I => \cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2\
        );

    \I__5368\ : InMux
    port map (
            O => \N__32838\,
            I => \N__32835\
        );

    \I__5367\ : LocalMux
    port map (
            O => \N__32835\,
            I => \N__32832\
        );

    \I__5366\ : Span4Mux_v
    port map (
            O => \N__32832\,
            I => \N__32829\
        );

    \I__5365\ : Odrv4
    port map (
            O => \N__32829\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2_8\
        );

    \I__5364\ : CascadeMux
    port map (
            O => \N__32826\,
            I => \N__32822\
        );

    \I__5363\ : InMux
    port map (
            O => \N__32825\,
            I => \N__32819\
        );

    \I__5362\ : InMux
    port map (
            O => \N__32822\,
            I => \N__32814\
        );

    \I__5361\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32811\
        );

    \I__5360\ : InMux
    port map (
            O => \N__32818\,
            I => \N__32806\
        );

    \I__5359\ : InMux
    port map (
            O => \N__32817\,
            I => \N__32806\
        );

    \I__5358\ : LocalMux
    port map (
            O => \N__32814\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845\
        );

    \I__5357\ : Odrv4
    port map (
            O => \N__32811\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845\
        );

    \I__5356\ : LocalMux
    port map (
            O => \N__32806\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845\
        );

    \I__5355\ : CascadeMux
    port map (
            O => \N__32799\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_0_1_cascade_\
        );

    \I__5354\ : InMux
    port map (
            O => \N__32796\,
            I => \N__32793\
        );

    \I__5353\ : LocalMux
    port map (
            O => \N__32793\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1873_0\
        );

    \I__5352\ : InMux
    port map (
            O => \N__32790\,
            I => \N__32787\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__32787\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1874_0\
        );

    \I__5350\ : InMux
    port map (
            O => \N__32784\,
            I => \N__32777\
        );

    \I__5349\ : InMux
    port map (
            O => \N__32783\,
            I => \N__32777\
        );

    \I__5348\ : InMux
    port map (
            O => \N__32782\,
            I => \N__32774\
        );

    \I__5347\ : LocalMux
    port map (
            O => \N__32777\,
            I => \N__32771\
        );

    \I__5346\ : LocalMux
    port map (
            O => \N__32774\,
            I => \N__32767\
        );

    \I__5345\ : Span4Mux_v
    port map (
            O => \N__32771\,
            I => \N__32764\
        );

    \I__5344\ : InMux
    port map (
            O => \N__32770\,
            I => \N__32761\
        );

    \I__5343\ : Span4Mux_v
    port map (
            O => \N__32767\,
            I => \N__32758\
        );

    \I__5342\ : Odrv4
    port map (
            O => \N__32764\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0\
        );

    \I__5341\ : LocalMux
    port map (
            O => \N__32761\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0\
        );

    \I__5340\ : Odrv4
    port map (
            O => \N__32758\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0\
        );

    \I__5339\ : InMux
    port map (
            O => \N__32751\,
            I => \N__32745\
        );

    \I__5338\ : InMux
    port map (
            O => \N__32750\,
            I => \N__32745\
        );

    \I__5337\ : LocalMux
    port map (
            O => \N__32745\,
            I => \N__32740\
        );

    \I__5336\ : ClkMux
    port map (
            O => \N__32744\,
            I => \N__32733\
        );

    \I__5335\ : ClkMux
    port map (
            O => \N__32743\,
            I => \N__32733\
        );

    \I__5334\ : Glb2LocalMux
    port map (
            O => \N__32740\,
            I => \N__32733\
        );

    \I__5333\ : GlobalMux
    port map (
            O => \N__32733\,
            I => \N__32730\
        );

    \I__5332\ : gio2CtrlBuf
    port map (
            O => \N__32730\,
            I => s_sda_i_g
        );

    \I__5331\ : InMux
    port map (
            O => \N__32727\,
            I => \N__32724\
        );

    \I__5330\ : LocalMux
    port map (
            O => \N__32724\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1392\
        );

    \I__5329\ : CascadeMux
    port map (
            O => \N__32721\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1381_0_cascade_\
        );

    \I__5328\ : CascadeMux
    port map (
            O => \N__32718\,
            I => \N__32715\
        );

    \I__5327\ : InMux
    port map (
            O => \N__32715\,
            I => \N__32712\
        );

    \I__5326\ : LocalMux
    port map (
            O => \N__32712\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392\
        );

    \I__5325\ : InMux
    port map (
            O => \N__32709\,
            I => \N__32706\
        );

    \I__5324\ : LocalMux
    port map (
            O => \N__32706\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_i_2_2\
        );

    \I__5323\ : CascadeMux
    port map (
            O => \N__32703\,
            I => \N__32699\
        );

    \I__5322\ : InMux
    port map (
            O => \N__32702\,
            I => \N__32693\
        );

    \I__5321\ : InMux
    port map (
            O => \N__32699\,
            I => \N__32688\
        );

    \I__5320\ : InMux
    port map (
            O => \N__32698\,
            I => \N__32688\
        );

    \I__5319\ : InMux
    port map (
            O => \N__32697\,
            I => \N__32685\
        );

    \I__5318\ : InMux
    port map (
            O => \N__32696\,
            I => \N__32682\
        );

    \I__5317\ : LocalMux
    port map (
            O => \N__32693\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__5316\ : LocalMux
    port map (
            O => \N__32688\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__5315\ : LocalMux
    port map (
            O => \N__32685\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__5314\ : LocalMux
    port map (
            O => \N__32682\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__5313\ : InMux
    port map (
            O => \N__32673\,
            I => \N__32668\
        );

    \I__5312\ : InMux
    port map (
            O => \N__32672\,
            I => \N__32661\
        );

    \I__5311\ : InMux
    port map (
            O => \N__32671\,
            I => \N__32661\
        );

    \I__5310\ : LocalMux
    port map (
            O => \N__32668\,
            I => \N__32658\
        );

    \I__5309\ : InMux
    port map (
            O => \N__32667\,
            I => \N__32653\
        );

    \I__5308\ : InMux
    port map (
            O => \N__32666\,
            I => \N__32653\
        );

    \I__5307\ : LocalMux
    port map (
            O => \N__32661\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17\
        );

    \I__5306\ : Odrv4
    port map (
            O => \N__32658\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17\
        );

    \I__5305\ : LocalMux
    port map (
            O => \N__32653\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17\
        );

    \I__5304\ : InMux
    port map (
            O => \N__32646\,
            I => \N__32643\
        );

    \I__5303\ : LocalMux
    port map (
            O => \N__32643\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_18\
        );

    \I__5302\ : CascadeMux
    port map (
            O => \N__32640\,
            I => \N__32637\
        );

    \I__5301\ : InMux
    port map (
            O => \N__32637\,
            I => \N__32626\
        );

    \I__5300\ : InMux
    port map (
            O => \N__32636\,
            I => \N__32626\
        );

    \I__5299\ : InMux
    port map (
            O => \N__32635\,
            I => \N__32621\
        );

    \I__5298\ : InMux
    port map (
            O => \N__32634\,
            I => \N__32621\
        );

    \I__5297\ : InMux
    port map (
            O => \N__32633\,
            I => \N__32618\
        );

    \I__5296\ : InMux
    port map (
            O => \N__32632\,
            I => \N__32613\
        );

    \I__5295\ : InMux
    port map (
            O => \N__32631\,
            I => \N__32613\
        );

    \I__5294\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32606\
        );

    \I__5293\ : LocalMux
    port map (
            O => \N__32621\,
            I => \N__32606\
        );

    \I__5292\ : LocalMux
    port map (
            O => \N__32618\,
            I => \N__32606\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__32613\,
            I => \N__32603\
        );

    \I__5290\ : Span4Mux_v
    port map (
            O => \N__32606\,
            I => \N__32599\
        );

    \I__5289\ : Span4Mux_v
    port map (
            O => \N__32603\,
            I => \N__32596\
        );

    \I__5288\ : InMux
    port map (
            O => \N__32602\,
            I => \N__32593\
        );

    \I__5287\ : Span4Mux_h
    port map (
            O => \N__32599\,
            I => \N__32588\
        );

    \I__5286\ : Span4Mux_h
    port map (
            O => \N__32596\,
            I => \N__32585\
        );

    \I__5285\ : LocalMux
    port map (
            O => \N__32593\,
            I => \N__32582\
        );

    \I__5284\ : InMux
    port map (
            O => \N__32592\,
            I => \N__32577\
        );

    \I__5283\ : InMux
    port map (
            O => \N__32591\,
            I => \N__32577\
        );

    \I__5282\ : Odrv4
    port map (
            O => \N__32588\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0\
        );

    \I__5281\ : Odrv4
    port map (
            O => \N__32585\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__32582\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0\
        );

    \I__5279\ : LocalMux
    port map (
            O => \N__32577\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0\
        );

    \I__5278\ : InMux
    port map (
            O => \N__32568\,
            I => \N__32561\
        );

    \I__5277\ : InMux
    port map (
            O => \N__32567\,
            I => \N__32561\
        );

    \I__5276\ : InMux
    port map (
            O => \N__32566\,
            I => \N__32558\
        );

    \I__5275\ : LocalMux
    port map (
            O => \N__32561\,
            I => \N__32552\
        );

    \I__5274\ : LocalMux
    port map (
            O => \N__32558\,
            I => \N__32552\
        );

    \I__5273\ : InMux
    port map (
            O => \N__32557\,
            I => \N__32549\
        );

    \I__5272\ : Span4Mux_v
    port map (
            O => \N__32552\,
            I => \N__32546\
        );

    \I__5271\ : LocalMux
    port map (
            O => \N__32549\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1\
        );

    \I__5270\ : Odrv4
    port map (
            O => \N__32546\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1\
        );

    \I__5269\ : InMux
    port map (
            O => \N__32541\,
            I => \N__32529\
        );

    \I__5268\ : InMux
    port map (
            O => \N__32540\,
            I => \N__32529\
        );

    \I__5267\ : InMux
    port map (
            O => \N__32539\,
            I => \N__32529\
        );

    \I__5266\ : InMux
    port map (
            O => \N__32538\,
            I => \N__32529\
        );

    \I__5265\ : LocalMux
    port map (
            O => \N__32529\,
            I => \N__32526\
        );

    \I__5264\ : Span4Mux_v
    port map (
            O => \N__32526\,
            I => \N__32523\
        );

    \I__5263\ : Odrv4
    port map (
            O => \N__32523\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_11_0_i_0_1\
        );

    \I__5262\ : CascadeMux
    port map (
            O => \N__32520\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_1394_cascade_\
        );

    \I__5261\ : CEMux
    port map (
            O => \N__32517\,
            I => \N__32513\
        );

    \I__5260\ : CEMux
    port map (
            O => \N__32516\,
            I => \N__32509\
        );

    \I__5259\ : LocalMux
    port map (
            O => \N__32513\,
            I => \N__32506\
        );

    \I__5258\ : CEMux
    port map (
            O => \N__32512\,
            I => \N__32503\
        );

    \I__5257\ : LocalMux
    port map (
            O => \N__32509\,
            I => \N__32500\
        );

    \I__5256\ : Span4Mux_v
    port map (
            O => \N__32506\,
            I => \N__32497\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__32503\,
            I => \N__32494\
        );

    \I__5254\ : Span4Mux_h
    port map (
            O => \N__32500\,
            I => \N__32491\
        );

    \I__5253\ : Sp12to4
    port map (
            O => \N__32497\,
            I => \N__32485\
        );

    \I__5252\ : Span4Mux_v
    port map (
            O => \N__32494\,
            I => \N__32482\
        );

    \I__5251\ : Span4Mux_h
    port map (
            O => \N__32491\,
            I => \N__32479\
        );

    \I__5250\ : CEMux
    port map (
            O => \N__32490\,
            I => \N__32476\
        );

    \I__5249\ : CEMux
    port map (
            O => \N__32489\,
            I => \N__32473\
        );

    \I__5248\ : CEMux
    port map (
            O => \N__32488\,
            I => \N__32470\
        );

    \I__5247\ : Span12Mux_h
    port map (
            O => \N__32485\,
            I => \N__32465\
        );

    \I__5246\ : Sp12to4
    port map (
            O => \N__32482\,
            I => \N__32465\
        );

    \I__5245\ : Span4Mux_v
    port map (
            O => \N__32479\,
            I => \N__32462\
        );

    \I__5244\ : LocalMux
    port map (
            O => \N__32476\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__32473\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\
        );

    \I__5242\ : LocalMux
    port map (
            O => \N__32470\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\
        );

    \I__5241\ : Odrv12
    port map (
            O => \N__32465\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\
        );

    \I__5240\ : Odrv4
    port map (
            O => \N__32462\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\
        );

    \I__5239\ : InMux
    port map (
            O => \N__32451\,
            I => \N__32448\
        );

    \I__5238\ : LocalMux
    port map (
            O => \N__32448\,
            I => \N__32445\
        );

    \I__5237\ : Span4Mux_h
    port map (
            O => \N__32445\,
            I => \N__32442\
        );

    \I__5236\ : Span4Mux_h
    port map (
            O => \N__32442\,
            I => \N__32439\
        );

    \I__5235\ : Span4Mux_v
    port map (
            O => \N__32439\,
            I => \N__32436\
        );

    \I__5234\ : Odrv4
    port map (
            O => \N__32436\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_16
        );

    \I__5233\ : CascadeMux
    port map (
            O => \N__32433\,
            I => \N__32430\
        );

    \I__5232\ : InMux
    port map (
            O => \N__32430\,
            I => \N__32427\
        );

    \I__5231\ : LocalMux
    port map (
            O => \N__32427\,
            I => \N__32424\
        );

    \I__5230\ : Span4Mux_v
    port map (
            O => \N__32424\,
            I => \N__32421\
        );

    \I__5229\ : Span4Mux_h
    port map (
            O => \N__32421\,
            I => \N__32418\
        );

    \I__5228\ : Span4Mux_h
    port map (
            O => \N__32418\,
            I => \N__32415\
        );

    \I__5227\ : Odrv4
    port map (
            O => \N__32415\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_18
        );

    \I__5226\ : InMux
    port map (
            O => \N__32412\,
            I => \N__32409\
        );

    \I__5225\ : LocalMux
    port map (
            O => \N__32409\,
            I => \N__32406\
        );

    \I__5224\ : Span4Mux_v
    port map (
            O => \N__32406\,
            I => \N__32403\
        );

    \I__5223\ : Odrv4
    port map (
            O => \N__32403\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1911\
        );

    \I__5222\ : InMux
    port map (
            O => \N__32400\,
            I => \N__32397\
        );

    \I__5221\ : LocalMux
    port map (
            O => \N__32397\,
            I => \N__32394\
        );

    \I__5220\ : Span4Mux_v
    port map (
            O => \N__32394\,
            I => \N__32391\
        );

    \I__5219\ : Span4Mux_h
    port map (
            O => \N__32391\,
            I => \N__32388\
        );

    \I__5218\ : Odrv4
    port map (
            O => \N__32388\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_8
        );

    \I__5217\ : CascadeMux
    port map (
            O => \N__32385\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0_cascade_\
        );

    \I__5216\ : InMux
    port map (
            O => \N__32382\,
            I => \N__32379\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__32379\,
            I => \N__32376\
        );

    \I__5214\ : Span4Mux_h
    port map (
            O => \N__32376\,
            I => \N__32373\
        );

    \I__5213\ : Span4Mux_v
    port map (
            O => \N__32373\,
            I => \N__32370\
        );

    \I__5212\ : Span4Mux_v
    port map (
            O => \N__32370\,
            I => \N__32367\
        );

    \I__5211\ : Odrv4
    port map (
            O => \N__32367\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1920\
        );

    \I__5210\ : InMux
    port map (
            O => \N__32364\,
            I => \N__32357\
        );

    \I__5209\ : InMux
    port map (
            O => \N__32363\,
            I => \N__32350\
        );

    \I__5208\ : InMux
    port map (
            O => \N__32362\,
            I => \N__32350\
        );

    \I__5207\ : InMux
    port map (
            O => \N__32361\,
            I => \N__32350\
        );

    \I__5206\ : InMux
    port map (
            O => \N__32360\,
            I => \N__32347\
        );

    \I__5205\ : LocalMux
    port map (
            O => \N__32357\,
            I => \N__32344\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__32350\,
            I => \N__32341\
        );

    \I__5203\ : LocalMux
    port map (
            O => \N__32347\,
            I => \N__32338\
        );

    \I__5202\ : Span4Mux_h
    port map (
            O => \N__32344\,
            I => \N__32331\
        );

    \I__5201\ : Span4Mux_h
    port map (
            O => \N__32341\,
            I => \N__32331\
        );

    \I__5200\ : Span4Mux_h
    port map (
            O => \N__32338\,
            I => \N__32328\
        );

    \I__5199\ : InMux
    port map (
            O => \N__32337\,
            I => \N__32323\
        );

    \I__5198\ : InMux
    port map (
            O => \N__32336\,
            I => \N__32323\
        );

    \I__5197\ : Span4Mux_v
    port map (
            O => \N__32331\,
            I => \N__32320\
        );

    \I__5196\ : Odrv4
    port map (
            O => \N__32328\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable
        );

    \I__5195\ : LocalMux
    port map (
            O => \N__32323\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable
        );

    \I__5194\ : Odrv4
    port map (
            O => \N__32320\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable
        );

    \I__5193\ : InMux
    port map (
            O => \N__32313\,
            I => \N__32306\
        );

    \I__5192\ : InMux
    port map (
            O => \N__32312\,
            I => \N__32306\
        );

    \I__5191\ : InMux
    port map (
            O => \N__32311\,
            I => \N__32303\
        );

    \I__5190\ : LocalMux
    port map (
            O => \N__32306\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0\
        );

    \I__5189\ : LocalMux
    port map (
            O => \N__32303\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0\
        );

    \I__5188\ : InMux
    port map (
            O => \N__32298\,
            I => \N__32294\
        );

    \I__5187\ : InMux
    port map (
            O => \N__32297\,
            I => \N__32291\
        );

    \I__5186\ : LocalMux
    port map (
            O => \N__32294\,
            I => \N__32288\
        );

    \I__5185\ : LocalMux
    port map (
            O => \N__32291\,
            I => \N__32285\
        );

    \I__5184\ : Span4Mux_h
    port map (
            O => \N__32288\,
            I => \N__32280\
        );

    \I__5183\ : Span4Mux_v
    port map (
            O => \N__32285\,
            I => \N__32280\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__32280\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m20_0_a2_4_1\
        );

    \I__5181\ : CascadeMux
    port map (
            O => \N__32277\,
            I => \N__32273\
        );

    \I__5180\ : CascadeMux
    port map (
            O => \N__32276\,
            I => \N__32268\
        );

    \I__5179\ : InMux
    port map (
            O => \N__32273\,
            I => \N__32265\
        );

    \I__5178\ : InMux
    port map (
            O => \N__32272\,
            I => \N__32260\
        );

    \I__5177\ : InMux
    port map (
            O => \N__32271\,
            I => \N__32260\
        );

    \I__5176\ : InMux
    port map (
            O => \N__32268\,
            I => \N__32257\
        );

    \I__5175\ : LocalMux
    port map (
            O => \N__32265\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__32260\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13\
        );

    \I__5173\ : LocalMux
    port map (
            O => \N__32257\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13\
        );

    \I__5172\ : IoInMux
    port map (
            O => \N__32250\,
            I => \N__32247\
        );

    \I__5171\ : LocalMux
    port map (
            O => \N__32247\,
            I => \N__32244\
        );

    \I__5170\ : Span4Mux_s2_h
    port map (
            O => \N__32244\,
            I => \N__32241\
        );

    \I__5169\ : Span4Mux_h
    port map (
            O => \N__32241\,
            I => \N__32238\
        );

    \I__5168\ : Span4Mux_h
    port map (
            O => \N__32238\,
            I => \N__32235\
        );

    \I__5167\ : Span4Mux_h
    port map (
            O => \N__32235\,
            I => \N__32232\
        );

    \I__5166\ : Odrv4
    port map (
            O => \N__32232\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa\
        );

    \I__5165\ : CascadeMux
    port map (
            O => \N__32229\,
            I => \N__32226\
        );

    \I__5164\ : InMux
    port map (
            O => \N__32226\,
            I => \N__32223\
        );

    \I__5163\ : LocalMux
    port map (
            O => \N__32223\,
            I => \N__32219\
        );

    \I__5162\ : InMux
    port map (
            O => \N__32222\,
            I => \N__32216\
        );

    \I__5161\ : Span12Mux_h
    port map (
            O => \N__32219\,
            I => \N__32213\
        );

    \I__5160\ : LocalMux
    port map (
            O => \N__32216\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_5
        );

    \I__5159\ : Odrv12
    port map (
            O => \N__32213\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_5
        );

    \I__5158\ : CascadeMux
    port map (
            O => \N__32208\,
            I => \N__32204\
        );

    \I__5157\ : InMux
    port map (
            O => \N__32207\,
            I => \N__32201\
        );

    \I__5156\ : InMux
    port map (
            O => \N__32204\,
            I => \N__32198\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__32201\,
            I => \N__32194\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__32198\,
            I => \N__32191\
        );

    \I__5153\ : InMux
    port map (
            O => \N__32197\,
            I => \N__32188\
        );

    \I__5152\ : Span4Mux_v
    port map (
            O => \N__32194\,
            I => \N__32185\
        );

    \I__5151\ : Span12Mux_v
    port map (
            O => \N__32191\,
            I => \N__32182\
        );

    \I__5150\ : LocalMux
    port map (
            O => \N__32188\,
            I => \N__32177\
        );

    \I__5149\ : Span4Mux_h
    port map (
            O => \N__32185\,
            I => \N__32177\
        );

    \I__5148\ : Odrv12
    port map (
            O => \N__32182\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_5
        );

    \I__5147\ : Odrv4
    port map (
            O => \N__32177\,
            I => cemf_module_64ch_ctrl_inst1_data_interrupts_5
        );

    \I__5146\ : CascadeMux
    port map (
            O => \N__32172\,
            I => \N__32167\
        );

    \I__5145\ : InMux
    port map (
            O => \N__32171\,
            I => \N__32164\
        );

    \I__5144\ : InMux
    port map (
            O => \N__32170\,
            I => \N__32161\
        );

    \I__5143\ : InMux
    port map (
            O => \N__32167\,
            I => \N__32158\
        );

    \I__5142\ : LocalMux
    port map (
            O => \N__32164\,
            I => \N__32155\
        );

    \I__5141\ : LocalMux
    port map (
            O => \N__32161\,
            I => \N__32152\
        );

    \I__5140\ : LocalMux
    port map (
            O => \N__32158\,
            I => \N__32149\
        );

    \I__5139\ : Odrv12
    port map (
            O => \N__32155\,
            I => cemf_module_64ch_ctrl_inst1_data_config_5
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__32152\,
            I => cemf_module_64ch_ctrl_inst1_data_config_5
        );

    \I__5137\ : Odrv4
    port map (
            O => \N__32149\,
            I => cemf_module_64ch_ctrl_inst1_data_config_5
        );

    \I__5136\ : CascadeMux
    port map (
            O => \N__32142\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_5_cascade_\
        );

    \I__5135\ : InMux
    port map (
            O => \N__32139\,
            I => \N__32136\
        );

    \I__5134\ : LocalMux
    port map (
            O => \N__32136\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRLZ0Z7\
        );

    \I__5133\ : InMux
    port map (
            O => \N__32133\,
            I => \N__32130\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__32130\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_5\
        );

    \I__5131\ : InMux
    port map (
            O => \N__32127\,
            I => \N__32124\
        );

    \I__5130\ : LocalMux
    port map (
            O => \N__32124\,
            I => \N__32120\
        );

    \I__5129\ : InMux
    port map (
            O => \N__32123\,
            I => \N__32117\
        );

    \I__5128\ : Span4Mux_h
    port map (
            O => \N__32120\,
            I => \N__32114\
        );

    \I__5127\ : LocalMux
    port map (
            O => \N__32117\,
            I => \N__32111\
        );

    \I__5126\ : Span4Mux_h
    port map (
            O => \N__32114\,
            I => \N__32105\
        );

    \I__5125\ : Span4Mux_h
    port map (
            O => \N__32111\,
            I => \N__32105\
        );

    \I__5124\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32102\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__32105\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_5
        );

    \I__5122\ : LocalMux
    port map (
            O => \N__32102\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_5
        );

    \I__5121\ : InMux
    port map (
            O => \N__32097\,
            I => \N__32094\
        );

    \I__5120\ : LocalMux
    port map (
            O => \N__32094\,
            I => \N__32091\
        );

    \I__5119\ : Span4Mux_v
    port map (
            O => \N__32091\,
            I => \N__32088\
        );

    \I__5118\ : Span4Mux_h
    port map (
            O => \N__32088\,
            I => \N__32085\
        );

    \I__5117\ : Sp12to4
    port map (
            O => \N__32085\,
            I => \N__32082\
        );

    \I__5116\ : Span12Mux_h
    port map (
            O => \N__32082\,
            I => \N__32077\
        );

    \I__5115\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32072\
        );

    \I__5114\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32072\
        );

    \I__5113\ : Odrv12
    port map (
            O => \N__32077\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_14
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__32072\,
            I => cemf_module_64ch_ctrl_inst1_data_clkctrovf_14
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__32067\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_242_cascade_\
        );

    \I__5110\ : InMux
    port map (
            O => \N__32064\,
            I => \N__32061\
        );

    \I__5109\ : LocalMux
    port map (
            O => \N__32061\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_6\
        );

    \I__5108\ : InMux
    port map (
            O => \N__32058\,
            I => \N__32052\
        );

    \I__5107\ : InMux
    port map (
            O => \N__32057\,
            I => \N__32052\
        );

    \I__5106\ : LocalMux
    port map (
            O => \N__32052\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_7\
        );

    \I__5105\ : InMux
    port map (
            O => \N__32049\,
            I => \N__32046\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__32046\,
            I => \N__32043\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__32043\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_6\
        );

    \I__5102\ : CascadeMux
    port map (
            O => \N__32040\,
            I => \N__32036\
        );

    \I__5101\ : InMux
    port map (
            O => \N__32039\,
            I => \N__32031\
        );

    \I__5100\ : InMux
    port map (
            O => \N__32036\,
            I => \N__32031\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__32031\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_6
        );

    \I__5098\ : InMux
    port map (
            O => \N__32028\,
            I => \N__32025\
        );

    \I__5097\ : LocalMux
    port map (
            O => \N__32025\,
            I => \N__32022\
        );

    \I__5096\ : Span4Mux_h
    port map (
            O => \N__32022\,
            I => \N__32019\
        );

    \I__5095\ : Span4Mux_v
    port map (
            O => \N__32019\,
            I => \N__32016\
        );

    \I__5094\ : Odrv4
    port map (
            O => \N__32016\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_283\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__32013\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_20_cascade_\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__32010\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_20_cascade_\
        );

    \I__5091\ : InMux
    port map (
            O => \N__32007\,
            I => \N__32004\
        );

    \I__5090\ : LocalMux
    port map (
            O => \N__32004\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_20\
        );

    \I__5089\ : InMux
    port map (
            O => \N__32001\,
            I => \N__31998\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__31998\,
            I => \N__31995\
        );

    \I__5087\ : Span4Mux_v
    port map (
            O => \N__31995\,
            I => \N__31992\
        );

    \I__5086\ : Odrv4
    port map (
            O => \N__31992\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_6\
        );

    \I__5085\ : InMux
    port map (
            O => \N__31989\,
            I => \N__31986\
        );

    \I__5084\ : LocalMux
    port map (
            O => \N__31986\,
            I => \N__31982\
        );

    \I__5083\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31978\
        );

    \I__5082\ : Span4Mux_h
    port map (
            O => \N__31982\,
            I => \N__31975\
        );

    \I__5081\ : InMux
    port map (
            O => \N__31981\,
            I => \N__31972\
        );

    \I__5080\ : LocalMux
    port map (
            O => \N__31978\,
            I => cemf_module_64ch_ctrl_inst1_data_config_6
        );

    \I__5079\ : Odrv4
    port map (
            O => \N__31975\,
            I => cemf_module_64ch_ctrl_inst1_data_config_6
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__31972\,
            I => cemf_module_64ch_ctrl_inst1_data_config_6
        );

    \I__5077\ : CascadeMux
    port map (
            O => \N__31965\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_6_cascade_\
        );

    \I__5076\ : CascadeMux
    port map (
            O => \N__31962\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SLZ0Z7_cascade_\
        );

    \I__5075\ : InMux
    port map (
            O => \N__31959\,
            I => \N__31956\
        );

    \I__5074\ : LocalMux
    port map (
            O => \N__31956\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRLZ0Z7\
        );

    \I__5073\ : InMux
    port map (
            O => \N__31953\,
            I => \N__31950\
        );

    \I__5072\ : LocalMux
    port map (
            O => \N__31950\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6\
        );

    \I__5071\ : InMux
    port map (
            O => \N__31947\,
            I => \N__31944\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__31944\,
            I => \N__31941\
        );

    \I__5069\ : Odrv4
    port map (
            O => \N__31941\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_5\
        );

    \I__5068\ : CascadeMux
    port map (
            O => \N__31938\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6_cascade_\
        );

    \I__5067\ : InMux
    port map (
            O => \N__31935\,
            I => \N__31932\
        );

    \I__5066\ : LocalMux
    port map (
            O => \N__31932\,
            I => \N__31929\
        );

    \I__5065\ : Span4Mux_v
    port map (
            O => \N__31929\,
            I => \N__31926\
        );

    \I__5064\ : Span4Mux_h
    port map (
            O => \N__31926\,
            I => \N__31923\
        );

    \I__5063\ : Span4Mux_h
    port map (
            O => \N__31923\,
            I => \N__31920\
        );

    \I__5062\ : Span4Mux_v
    port map (
            O => \N__31920\,
            I => \N__31917\
        );

    \I__5061\ : Odrv4
    port map (
            O => \N__31917\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_11
        );

    \I__5060\ : CascadeMux
    port map (
            O => \N__31914\,
            I => \N__31911\
        );

    \I__5059\ : InMux
    port map (
            O => \N__31911\,
            I => \N__31908\
        );

    \I__5058\ : LocalMux
    port map (
            O => \N__31908\,
            I => \N__31905\
        );

    \I__5057\ : Span4Mux_v
    port map (
            O => \N__31905\,
            I => \N__31902\
        );

    \I__5056\ : Span4Mux_v
    port map (
            O => \N__31902\,
            I => \N__31899\
        );

    \I__5055\ : Sp12to4
    port map (
            O => \N__31899\,
            I => \N__31896\
        );

    \I__5054\ : Odrv12
    port map (
            O => \N__31896\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_11
        );

    \I__5053\ : CascadeMux
    port map (
            O => \N__31893\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_11_cascade_\
        );

    \I__5052\ : InMux
    port map (
            O => \N__31890\,
            I => \N__31887\
        );

    \I__5051\ : LocalMux
    port map (
            O => \N__31887\,
            I => \N__31884\
        );

    \I__5050\ : Span4Mux_v
    port map (
            O => \N__31884\,
            I => \N__31881\
        );

    \I__5049\ : Span4Mux_h
    port map (
            O => \N__31881\,
            I => \N__31878\
        );

    \I__5048\ : Span4Mux_h
    port map (
            O => \N__31878\,
            I => \N__31875\
        );

    \I__5047\ : Odrv4
    port map (
            O => \N__31875\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_11
        );

    \I__5046\ : InMux
    port map (
            O => \N__31872\,
            I => \N__31869\
        );

    \I__5045\ : LocalMux
    port map (
            O => \N__31869\,
            I => \N__31866\
        );

    \I__5044\ : Span4Mux_v
    port map (
            O => \N__31866\,
            I => \N__31863\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__31863\,
            I => \N__31860\
        );

    \I__5042\ : Odrv4
    port map (
            O => \N__31860\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_819\
        );

    \I__5041\ : CascadeMux
    port map (
            O => \N__31857\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_11_cascade_\
        );

    \I__5040\ : InMux
    port map (
            O => \N__31854\,
            I => \N__31851\
        );

    \I__5039\ : LocalMux
    port map (
            O => \N__31851\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_11\
        );

    \I__5038\ : InMux
    port map (
            O => \N__31848\,
            I => \N__31845\
        );

    \I__5037\ : LocalMux
    port map (
            O => \N__31845\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_11\
        );

    \I__5036\ : CascadeMux
    port map (
            O => \N__31842\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_11_cascade_\
        );

    \I__5035\ : InMux
    port map (
            O => \N__31839\,
            I => \N__31836\
        );

    \I__5034\ : LocalMux
    port map (
            O => \N__31836\,
            I => \N__31833\
        );

    \I__5033\ : Span4Mux_h
    port map (
            O => \N__31833\,
            I => \N__31830\
        );

    \I__5032\ : Span4Mux_h
    port map (
            O => \N__31830\,
            I => \N__31827\
        );

    \I__5031\ : Span4Mux_v
    port map (
            O => \N__31827\,
            I => \N__31824\
        );

    \I__5030\ : Odrv4
    port map (
            O => \N__31824\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_19
        );

    \I__5029\ : InMux
    port map (
            O => \N__31821\,
            I => \N__31818\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__31818\,
            I => \N__31815\
        );

    \I__5027\ : Span4Mux_h
    port map (
            O => \N__31815\,
            I => \N__31812\
        );

    \I__5026\ : Span4Mux_h
    port map (
            O => \N__31812\,
            I => \N__31809\
        );

    \I__5025\ : Span4Mux_v
    port map (
            O => \N__31809\,
            I => \N__31806\
        );

    \I__5024\ : Odrv4
    port map (
            O => \N__31806\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_20
        );

    \I__5023\ : CascadeMux
    port map (
            O => \N__31803\,
            I => \N__31800\
        );

    \I__5022\ : InMux
    port map (
            O => \N__31800\,
            I => \N__31797\
        );

    \I__5021\ : LocalMux
    port map (
            O => \N__31797\,
            I => \N__31794\
        );

    \I__5020\ : Span4Mux_v
    port map (
            O => \N__31794\,
            I => \N__31791\
        );

    \I__5019\ : Span4Mux_h
    port map (
            O => \N__31791\,
            I => \N__31788\
        );

    \I__5018\ : Odrv4
    port map (
            O => \N__31788\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_20
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__31785\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_20_cascade_\
        );

    \I__5016\ : InMux
    port map (
            O => \N__31782\,
            I => \N__31779\
        );

    \I__5015\ : LocalMux
    port map (
            O => \N__31779\,
            I => \N__31776\
        );

    \I__5014\ : Span4Mux_h
    port map (
            O => \N__31776\,
            I => \N__31773\
        );

    \I__5013\ : Span4Mux_h
    port map (
            O => \N__31773\,
            I => \N__31770\
        );

    \I__5012\ : Span4Mux_h
    port map (
            O => \N__31770\,
            I => \N__31767\
        );

    \I__5011\ : Odrv4
    port map (
            O => \N__31767\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_20
        );

    \I__5010\ : CascadeMux
    port map (
            O => \N__31764\,
            I => \N__31761\
        );

    \I__5009\ : InMux
    port map (
            O => \N__31761\,
            I => \N__31758\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__31758\,
            I => \N__31755\
        );

    \I__5007\ : Span4Mux_h
    port map (
            O => \N__31755\,
            I => \N__31752\
        );

    \I__5006\ : Span4Mux_h
    port map (
            O => \N__31752\,
            I => \N__31749\
        );

    \I__5005\ : Odrv4
    port map (
            O => \N__31749\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_2
        );

    \I__5004\ : CascadeMux
    port map (
            O => \N__31746\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_2_cascade_\
        );

    \I__5003\ : CascadeMux
    port map (
            O => \N__31743\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_2_cascade_\
        );

    \I__5002\ : InMux
    port map (
            O => \N__31740\,
            I => \N__31737\
        );

    \I__5001\ : LocalMux
    port map (
            O => \N__31737\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_2\
        );

    \I__5000\ : InMux
    port map (
            O => \N__31734\,
            I => \N__31731\
        );

    \I__4999\ : LocalMux
    port map (
            O => \N__31731\,
            I => \N__31728\
        );

    \I__4998\ : Span4Mux_h
    port map (
            O => \N__31728\,
            I => \N__31725\
        );

    \I__4997\ : Span4Mux_v
    port map (
            O => \N__31725\,
            I => \N__31722\
        );

    \I__4996\ : Span4Mux_v
    port map (
            O => \N__31722\,
            I => \N__31719\
        );

    \I__4995\ : Odrv4
    port map (
            O => \N__31719\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_10
        );

    \I__4994\ : CascadeMux
    port map (
            O => \N__31716\,
            I => \N__31713\
        );

    \I__4993\ : InMux
    port map (
            O => \N__31713\,
            I => \N__31710\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__31710\,
            I => \N__31707\
        );

    \I__4991\ : Span4Mux_v
    port map (
            O => \N__31707\,
            I => \N__31704\
        );

    \I__4990\ : Span4Mux_h
    port map (
            O => \N__31704\,
            I => \N__31701\
        );

    \I__4989\ : Odrv4
    port map (
            O => \N__31701\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_10
        );

    \I__4988\ : CascadeMux
    port map (
            O => \N__31698\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_10_cascade_\
        );

    \I__4987\ : InMux
    port map (
            O => \N__31695\,
            I => \N__31692\
        );

    \I__4986\ : LocalMux
    port map (
            O => \N__31692\,
            I => \N__31689\
        );

    \I__4985\ : Span4Mux_h
    port map (
            O => \N__31689\,
            I => \N__31686\
        );

    \I__4984\ : Span4Mux_h
    port map (
            O => \N__31686\,
            I => \N__31683\
        );

    \I__4983\ : Span4Mux_v
    port map (
            O => \N__31683\,
            I => \N__31680\
        );

    \I__4982\ : Odrv4
    port map (
            O => \N__31680\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_10
        );

    \I__4981\ : InMux
    port map (
            O => \N__31677\,
            I => \N__31674\
        );

    \I__4980\ : LocalMux
    port map (
            O => \N__31674\,
            I => \N__31671\
        );

    \I__4979\ : Odrv12
    port map (
            O => \N__31671\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_830\
        );

    \I__4978\ : CascadeMux
    port map (
            O => \N__31668\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_10_cascade_\
        );

    \I__4977\ : InMux
    port map (
            O => \N__31665\,
            I => \N__31662\
        );

    \I__4976\ : LocalMux
    port map (
            O => \N__31662\,
            I => \N__31659\
        );

    \I__4975\ : Span4Mux_h
    port map (
            O => \N__31659\,
            I => \N__31656\
        );

    \I__4974\ : Odrv4
    port map (
            O => \N__31656\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_10\
        );

    \I__4973\ : CascadeMux
    port map (
            O => \N__31653\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_10_cascade_\
        );

    \I__4972\ : InMux
    port map (
            O => \N__31650\,
            I => \N__31647\
        );

    \I__4971\ : LocalMux
    port map (
            O => \N__31647\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_10\
        );

    \I__4970\ : InMux
    port map (
            O => \N__31644\,
            I => \N__31641\
        );

    \I__4969\ : LocalMux
    port map (
            O => \N__31641\,
            I => \N__31638\
        );

    \I__4968\ : Span4Mux_v
    port map (
            O => \N__31638\,
            I => \N__31635\
        );

    \I__4967\ : Span4Mux_v
    port map (
            O => \N__31635\,
            I => \N__31632\
        );

    \I__4966\ : Sp12to4
    port map (
            O => \N__31632\,
            I => \N__31629\
        );

    \I__4965\ : Odrv12
    port map (
            O => \N__31629\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_18
        );

    \I__4964\ : CascadeMux
    port map (
            O => \N__31626\,
            I => \N__31623\
        );

    \I__4963\ : InMux
    port map (
            O => \N__31623\,
            I => \N__31620\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__31620\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_18\
        );

    \I__4961\ : InMux
    port map (
            O => \N__31617\,
            I => \N__31614\
        );

    \I__4960\ : LocalMux
    port map (
            O => \N__31614\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_3\
        );

    \I__4959\ : InMux
    port map (
            O => \N__31611\,
            I => \N__31608\
        );

    \I__4958\ : LocalMux
    port map (
            O => \N__31608\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_2\
        );

    \I__4957\ : InMux
    port map (
            O => \N__31605\,
            I => \N__31602\
        );

    \I__4956\ : LocalMux
    port map (
            O => \N__31602\,
            I => \N__31599\
        );

    \I__4955\ : Odrv12
    port map (
            O => \N__31599\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_275_0\
        );

    \I__4954\ : CascadeMux
    port map (
            O => \N__31596\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_275_0_cascade_\
        );

    \I__4953\ : CascadeMux
    port map (
            O => \N__31593\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_2_cascade_\
        );

    \I__4952\ : CascadeMux
    port map (
            O => \N__31590\,
            I => \N__31586\
        );

    \I__4951\ : InMux
    port map (
            O => \N__31589\,
            I => \N__31583\
        );

    \I__4950\ : InMux
    port map (
            O => \N__31586\,
            I => \N__31580\
        );

    \I__4949\ : LocalMux
    port map (
            O => \N__31583\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_59\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__31580\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.N_59\
        );

    \I__4947\ : InMux
    port map (
            O => \N__31575\,
            I => \N__31572\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__31572\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_2\
        );

    \I__4945\ : InMux
    port map (
            O => \N__31569\,
            I => \N__31566\
        );

    \I__4944\ : LocalMux
    port map (
            O => \N__31566\,
            I => \N__31563\
        );

    \I__4943\ : Span4Mux_v
    port map (
            O => \N__31563\,
            I => \N__31560\
        );

    \I__4942\ : Span4Mux_h
    port map (
            O => \N__31560\,
            I => \N__31557\
        );

    \I__4941\ : Span4Mux_h
    port map (
            O => \N__31557\,
            I => \N__31554\
        );

    \I__4940\ : Odrv4
    port map (
            O => \N__31554\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_2
        );

    \I__4939\ : InMux
    port map (
            O => \N__31551\,
            I => \N__31548\
        );

    \I__4938\ : LocalMux
    port map (
            O => \N__31548\,
            I => \N__31545\
        );

    \I__4937\ : Span4Mux_h
    port map (
            O => \N__31545\,
            I => \N__31542\
        );

    \I__4936\ : Odrv4
    port map (
            O => \N__31542\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1945\
        );

    \I__4935\ : CascadeMux
    port map (
            O => \N__31539\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2_cascade_\
        );

    \I__4934\ : InMux
    port map (
            O => \N__31536\,
            I => \N__31533\
        );

    \I__4933\ : LocalMux
    port map (
            O => \N__31533\,
            I => \N__31530\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__31530\,
            I => \N__31527\
        );

    \I__4931\ : Odrv4
    port map (
            O => \N__31527\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1844\
        );

    \I__4930\ : IoInMux
    port map (
            O => \N__31524\,
            I => \N__31521\
        );

    \I__4929\ : LocalMux
    port map (
            O => \N__31521\,
            I => \N__31518\
        );

    \I__4928\ : Span4Mux_s1_h
    port map (
            O => \N__31518\,
            I => \N__31515\
        );

    \I__4927\ : Span4Mux_h
    port map (
            O => \N__31515\,
            I => \N__31512\
        );

    \I__4926\ : Span4Mux_h
    port map (
            O => \N__31512\,
            I => \N__31509\
        );

    \I__4925\ : Span4Mux_h
    port map (
            O => \N__31509\,
            I => \N__31506\
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__31506\,
            I => \N_528_0\
        );

    \I__4923\ : InMux
    port map (
            O => \N__31503\,
            I => \N__31500\
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__31500\,
            I => \N__31497\
        );

    \I__4921\ : Odrv4
    port map (
            O => \N__31497\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_0\
        );

    \I__4920\ : InMux
    port map (
            O => \N__31494\,
            I => \N__31491\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__31491\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_2\
        );

    \I__4918\ : InMux
    port map (
            O => \N__31488\,
            I => \N__31482\
        );

    \I__4917\ : InMux
    port map (
            O => \N__31487\,
            I => \N__31482\
        );

    \I__4916\ : LocalMux
    port map (
            O => \N__31482\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_1\
        );

    \I__4915\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31474\
        );

    \I__4914\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31471\
        );

    \I__4913\ : InMux
    port map (
            O => \N__31477\,
            I => \N__31468\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__31474\,
            I => \N__31465\
        );

    \I__4911\ : LocalMux
    port map (
            O => \N__31471\,
            I => \cemf_module_64ch_ctrl_inst1.n_state41\
        );

    \I__4910\ : LocalMux
    port map (
            O => \N__31468\,
            I => \cemf_module_64ch_ctrl_inst1.n_state41\
        );

    \I__4909\ : Odrv4
    port map (
            O => \N__31465\,
            I => \cemf_module_64ch_ctrl_inst1.n_state41\
        );

    \I__4908\ : CascadeMux
    port map (
            O => \N__31458\,
            I => \N__31452\
        );

    \I__4907\ : CascadeMux
    port map (
            O => \N__31457\,
            I => \N__31448\
        );

    \I__4906\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31445\
        );

    \I__4905\ : CascadeMux
    port map (
            O => \N__31455\,
            I => \N__31442\
        );

    \I__4904\ : InMux
    port map (
            O => \N__31452\,
            I => \N__31439\
        );

    \I__4903\ : InMux
    port map (
            O => \N__31451\,
            I => \N__31436\
        );

    \I__4902\ : InMux
    port map (
            O => \N__31448\,
            I => \N__31433\
        );

    \I__4901\ : LocalMux
    port map (
            O => \N__31445\,
            I => \N__31430\
        );

    \I__4900\ : InMux
    port map (
            O => \N__31442\,
            I => \N__31427\
        );

    \I__4899\ : LocalMux
    port map (
            O => \N__31439\,
            I => \N__31418\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__31436\,
            I => \N__31418\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__31433\,
            I => \N__31418\
        );

    \I__4896\ : Span4Mux_h
    port map (
            O => \N__31430\,
            I => \N__31418\
        );

    \I__4895\ : LocalMux
    port map (
            O => \N__31427\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_19\
        );

    \I__4894\ : Odrv4
    port map (
            O => \N__31418\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_19\
        );

    \I__4893\ : InMux
    port map (
            O => \N__31413\,
            I => \N__31410\
        );

    \I__4892\ : LocalMux
    port map (
            O => \N__31410\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_1\
        );

    \I__4891\ : InMux
    port map (
            O => \N__31407\,
            I => \N__31404\
        );

    \I__4890\ : LocalMux
    port map (
            O => \N__31404\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_0\
        );

    \I__4889\ : InMux
    port map (
            O => \N__31401\,
            I => \N__31398\
        );

    \I__4888\ : LocalMux
    port map (
            O => \N__31398\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_1\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__31395\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1_cascade_\
        );

    \I__4886\ : InMux
    port map (
            O => \N__31392\,
            I => \N__31389\
        );

    \I__4885\ : LocalMux
    port map (
            O => \N__31389\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_1\
        );

    \I__4884\ : InMux
    port map (
            O => \N__31386\,
            I => \N__31378\
        );

    \I__4883\ : InMux
    port map (
            O => \N__31385\,
            I => \N__31378\
        );

    \I__4882\ : InMux
    port map (
            O => \N__31384\,
            I => \N__31375\
        );

    \I__4881\ : InMux
    port map (
            O => \N__31383\,
            I => \N__31372\
        );

    \I__4880\ : LocalMux
    port map (
            O => \N__31378\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3\
        );

    \I__4879\ : LocalMux
    port map (
            O => \N__31375\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__31372\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3\
        );

    \I__4877\ : CascadeMux
    port map (
            O => \N__31365\,
            I => \N__31361\
        );

    \I__4876\ : InMux
    port map (
            O => \N__31364\,
            I => \N__31358\
        );

    \I__4875\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31355\
        );

    \I__4874\ : LocalMux
    port map (
            O => \N__31358\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2\
        );

    \I__4873\ : LocalMux
    port map (
            O => \N__31355\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2\
        );

    \I__4872\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31347\
        );

    \I__4871\ : LocalMux
    port map (
            O => \N__31347\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_4\
        );

    \I__4870\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31340\
        );

    \I__4869\ : CascadeMux
    port map (
            O => \N__31343\,
            I => \N__31337\
        );

    \I__4868\ : LocalMux
    port map (
            O => \N__31340\,
            I => \N__31333\
        );

    \I__4867\ : InMux
    port map (
            O => \N__31337\,
            I => \N__31330\
        );

    \I__4866\ : InMux
    port map (
            O => \N__31336\,
            I => \N__31327\
        );

    \I__4865\ : Odrv12
    port map (
            O => \N__31333\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__31330\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__31327\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967\
        );

    \I__4862\ : CascadeMux
    port map (
            O => \N__31320\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_2_cascade_\
        );

    \I__4861\ : CascadeMux
    port map (
            O => \N__31317\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_3_cascade_\
        );

    \I__4860\ : InMux
    port map (
            O => \N__31314\,
            I => \N__31311\
        );

    \I__4859\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31308\
        );

    \I__4858\ : Span4Mux_v
    port map (
            O => \N__31308\,
            I => \N__31305\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__31305\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2\
        );

    \I__4856\ : CascadeMux
    port map (
            O => \N__31302\,
            I => \N__31298\
        );

    \I__4855\ : InMux
    port map (
            O => \N__31301\,
            I => \N__31293\
        );

    \I__4854\ : InMux
    port map (
            O => \N__31298\,
            I => \N__31293\
        );

    \I__4853\ : LocalMux
    port map (
            O => \N__31293\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_14\
        );

    \I__4852\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31287\
        );

    \I__4851\ : LocalMux
    port map (
            O => \N__31287\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_14\
        );

    \I__4850\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31275\
        );

    \I__4849\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31275\
        );

    \I__4848\ : InMux
    port map (
            O => \N__31282\,
            I => \N__31268\
        );

    \I__4847\ : InMux
    port map (
            O => \N__31281\,
            I => \N__31268\
        );

    \I__4846\ : InMux
    port map (
            O => \N__31280\,
            I => \N__31268\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__31275\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__31268\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12\
        );

    \I__4843\ : InMux
    port map (
            O => \N__31263\,
            I => \N__31248\
        );

    \I__4842\ : InMux
    port map (
            O => \N__31262\,
            I => \N__31248\
        );

    \I__4841\ : InMux
    port map (
            O => \N__31261\,
            I => \N__31248\
        );

    \I__4840\ : InMux
    port map (
            O => \N__31260\,
            I => \N__31241\
        );

    \I__4839\ : InMux
    port map (
            O => \N__31259\,
            I => \N__31241\
        );

    \I__4838\ : InMux
    port map (
            O => \N__31258\,
            I => \N__31241\
        );

    \I__4837\ : InMux
    port map (
            O => \N__31257\,
            I => \N__31234\
        );

    \I__4836\ : InMux
    port map (
            O => \N__31256\,
            I => \N__31234\
        );

    \I__4835\ : InMux
    port map (
            O => \N__31255\,
            I => \N__31234\
        );

    \I__4834\ : LocalMux
    port map (
            O => \N__31248\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987\
        );

    \I__4833\ : LocalMux
    port map (
            O => \N__31241\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__31234\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987\
        );

    \I__4831\ : CascadeMux
    port map (
            O => \N__31227\,
            I => \N__31222\
        );

    \I__4830\ : CascadeMux
    port map (
            O => \N__31226\,
            I => \N__31219\
        );

    \I__4829\ : InMux
    port map (
            O => \N__31225\,
            I => \N__31215\
        );

    \I__4828\ : InMux
    port map (
            O => \N__31222\,
            I => \N__31208\
        );

    \I__4827\ : InMux
    port map (
            O => \N__31219\,
            I => \N__31208\
        );

    \I__4826\ : InMux
    port map (
            O => \N__31218\,
            I => \N__31208\
        );

    \I__4825\ : LocalMux
    port map (
            O => \N__31215\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15\
        );

    \I__4824\ : LocalMux
    port map (
            O => \N__31208\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15\
        );

    \I__4823\ : CascadeMux
    port map (
            O => \N__31203\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967i_cascade_\
        );

    \I__4822\ : InMux
    port map (
            O => \N__31200\,
            I => \N__31197\
        );

    \I__4821\ : LocalMux
    port map (
            O => \N__31197\,
            I => \N__31194\
        );

    \I__4820\ : Odrv4
    port map (
            O => \N__31194\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retZ0Z_13\
        );

    \I__4819\ : InMux
    port map (
            O => \N__31191\,
            I => \N__31188\
        );

    \I__4818\ : LocalMux
    port map (
            O => \N__31188\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_276_reti\
        );

    \I__4817\ : CascadeMux
    port map (
            O => \N__31185\,
            I => \N__31181\
        );

    \I__4816\ : InMux
    port map (
            O => \N__31184\,
            I => \N__31176\
        );

    \I__4815\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31176\
        );

    \I__4814\ : LocalMux
    port map (
            O => \N__31176\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_8_1\
        );

    \I__4813\ : InMux
    port map (
            O => \N__31173\,
            I => \N__31168\
        );

    \I__4812\ : InMux
    port map (
            O => \N__31172\,
            I => \N__31163\
        );

    \I__4811\ : InMux
    port map (
            O => \N__31171\,
            I => \N__31163\
        );

    \I__4810\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31157\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__31163\,
            I => \N__31154\
        );

    \I__4808\ : InMux
    port map (
            O => \N__31162\,
            I => \N__31147\
        );

    \I__4807\ : InMux
    port map (
            O => \N__31161\,
            I => \N__31147\
        );

    \I__4806\ : InMux
    port map (
            O => \N__31160\,
            I => \N__31147\
        );

    \I__4805\ : Odrv4
    port map (
            O => \N__31157\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8\
        );

    \I__4804\ : Odrv4
    port map (
            O => \N__31154\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__31147\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8\
        );

    \I__4802\ : InMux
    port map (
            O => \N__31140\,
            I => \N__31134\
        );

    \I__4801\ : InMux
    port map (
            O => \N__31139\,
            I => \N__31134\
        );

    \I__4800\ : LocalMux
    port map (
            O => \N__31134\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1\
        );

    \I__4799\ : InMux
    port map (
            O => \N__31131\,
            I => \N__31128\
        );

    \I__4798\ : LocalMux
    port map (
            O => \N__31128\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_6\
        );

    \I__4797\ : CascadeMux
    port map (
            O => \N__31125\,
            I => \N__31120\
        );

    \I__4796\ : InMux
    port map (
            O => \N__31124\,
            I => \N__31116\
        );

    \I__4795\ : InMux
    port map (
            O => \N__31123\,
            I => \N__31113\
        );

    \I__4794\ : InMux
    port map (
            O => \N__31120\,
            I => \N__31108\
        );

    \I__4793\ : InMux
    port map (
            O => \N__31119\,
            I => \N__31108\
        );

    \I__4792\ : LocalMux
    port map (
            O => \N__31116\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7\
        );

    \I__4791\ : LocalMux
    port map (
            O => \N__31113\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7\
        );

    \I__4790\ : LocalMux
    port map (
            O => \N__31108\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__31101\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.en_count_bits_0_i_a2_0_a2_1_cascade_\
        );

    \I__4788\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31095\
        );

    \I__4787\ : LocalMux
    port map (
            O => \N__31095\,
            I => \N__31092\
        );

    \I__4786\ : Span4Mux_v
    port map (
            O => \N__31092\,
            I => \N__31083\
        );

    \I__4785\ : InMux
    port map (
            O => \N__31091\,
            I => \N__31078\
        );

    \I__4784\ : InMux
    port map (
            O => \N__31090\,
            I => \N__31078\
        );

    \I__4783\ : InMux
    port map (
            O => \N__31089\,
            I => \N__31071\
        );

    \I__4782\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31071\
        );

    \I__4781\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31071\
        );

    \I__4780\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31068\
        );

    \I__4779\ : Span4Mux_h
    port map (
            O => \N__31083\,
            I => \N__31061\
        );

    \I__4778\ : LocalMux
    port map (
            O => \N__31078\,
            I => \N__31061\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__31071\,
            I => \N__31061\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__31068\,
            I => \N__31056\
        );

    \I__4775\ : Span4Mux_h
    port map (
            O => \N__31061\,
            I => \N__31056\
        );

    \I__4774\ : Odrv4
    port map (
            O => \N__31056\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_277_0\
        );

    \I__4773\ : InMux
    port map (
            O => \N__31053\,
            I => \N__31044\
        );

    \I__4772\ : InMux
    port map (
            O => \N__31052\,
            I => \N__31044\
        );

    \I__4771\ : InMux
    port map (
            O => \N__31051\,
            I => \N__31044\
        );

    \I__4770\ : LocalMux
    port map (
            O => \N__31044\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_19\
        );

    \I__4769\ : InMux
    port map (
            O => \N__31041\,
            I => \N__31038\
        );

    \I__4768\ : LocalMux
    port map (
            O => \N__31038\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_18\
        );

    \I__4767\ : InMux
    port map (
            O => \N__31035\,
            I => \N__31032\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__31032\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_13\
        );

    \I__4765\ : InMux
    port map (
            O => \N__31029\,
            I => \N__31023\
        );

    \I__4764\ : InMux
    port map (
            O => \N__31028\,
            I => \N__31020\
        );

    \I__4763\ : InMux
    port map (
            O => \N__31027\,
            I => \N__31017\
        );

    \I__4762\ : InMux
    port map (
            O => \N__31026\,
            I => \N__31014\
        );

    \I__4761\ : LocalMux
    port map (
            O => \N__31023\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11\
        );

    \I__4760\ : LocalMux
    port map (
            O => \N__31020\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__31017\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11\
        );

    \I__4758\ : LocalMux
    port map (
            O => \N__31014\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11\
        );

    \I__4757\ : SRMux
    port map (
            O => \N__31005\,
            I => \N__31002\
        );

    \I__4756\ : LocalMux
    port map (
            O => \N__31002\,
            I => \N__30999\
        );

    \I__4755\ : Span4Mux_v
    port map (
            O => \N__30999\,
            I => \N__30996\
        );

    \I__4754\ : Span4Mux_h
    port map (
            O => \N__30996\,
            I => \N__30993\
        );

    \I__4753\ : Odrv4
    port map (
            O => \N__30993\,
            I => \I2C_top_level_inst1.I2C_Control_StartUp_inst.N_8_i\
        );

    \I__4752\ : InMux
    port map (
            O => \N__30990\,
            I => \N__30986\
        );

    \I__4751\ : InMux
    port map (
            O => \N__30989\,
            I => \N__30983\
        );

    \I__4750\ : LocalMux
    port map (
            O => \N__30986\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1\
        );

    \I__4749\ : LocalMux
    port map (
            O => \N__30983\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1\
        );

    \I__4748\ : InMux
    port map (
            O => \N__30978\,
            I => \N__30975\
        );

    \I__4747\ : LocalMux
    port map (
            O => \N__30975\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0\
        );

    \I__4746\ : CascadeMux
    port map (
            O => \N__30972\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0_cascade_\
        );

    \I__4745\ : InMux
    port map (
            O => \N__30969\,
            I => \N__30966\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__30966\,
            I => \N__30963\
        );

    \I__4743\ : Span4Mux_v
    port map (
            O => \N__30963\,
            I => \N__30959\
        );

    \I__4742\ : InMux
    port map (
            O => \N__30962\,
            I => \N__30956\
        );

    \I__4741\ : Span4Mux_h
    port map (
            O => \N__30959\,
            I => \N__30953\
        );

    \I__4740\ : LocalMux
    port map (
            O => \N__30956\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26\
        );

    \I__4739\ : Odrv4
    port map (
            O => \N__30953\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26\
        );

    \I__4738\ : CascadeMux
    port map (
            O => \N__30948\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3Z0Z_0_cascade_\
        );

    \I__4737\ : CascadeMux
    port map (
            O => \N__30945\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1959_cascade_\
        );

    \I__4736\ : CascadeMux
    port map (
            O => \N__30942\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0_cascade_\
        );

    \I__4735\ : CascadeMux
    port map (
            O => \N__30939\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRLZ0Z7_cascade_\
        );

    \I__4734\ : InMux
    port map (
            O => \N__30936\,
            I => \N__30933\
        );

    \I__4733\ : LocalMux
    port map (
            O => \N__30933\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3\
        );

    \I__4732\ : CascadeMux
    port map (
            O => \N__30930\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3_cascade_\
        );

    \I__4731\ : InMux
    port map (
            O => \N__30927\,
            I => \N__30924\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__30924\,
            I => \N__30921\
        );

    \I__4729\ : Odrv4
    port map (
            O => \N__30921\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5\
        );

    \I__4728\ : CascadeMux
    port map (
            O => \N__30918\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5_cascade_\
        );

    \I__4727\ : InMux
    port map (
            O => \N__30915\,
            I => \N__30912\
        );

    \I__4726\ : LocalMux
    port map (
            O => \N__30912\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_3\
        );

    \I__4725\ : InMux
    port map (
            O => \N__30909\,
            I => \N__30906\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__30906\,
            I => \N__30902\
        );

    \I__4723\ : InMux
    port map (
            O => \N__30905\,
            I => \N__30899\
        );

    \I__4722\ : Span4Mux_h
    port map (
            O => \N__30902\,
            I => \N__30896\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__30899\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4\
        );

    \I__4720\ : Odrv4
    port map (
            O => \N__30896\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4\
        );

    \I__4719\ : InMux
    port map (
            O => \N__30891\,
            I => \N__30888\
        );

    \I__4718\ : LocalMux
    port map (
            O => \N__30888\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_4\
        );

    \I__4717\ : InMux
    port map (
            O => \N__30885\,
            I => \N__30882\
        );

    \I__4716\ : LocalMux
    port map (
            O => \N__30882\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_9\
        );

    \I__4715\ : CascadeMux
    port map (
            O => \N__30879\,
            I => \N__30875\
        );

    \I__4714\ : InMux
    port map (
            O => \N__30878\,
            I => \N__30870\
        );

    \I__4713\ : InMux
    port map (
            O => \N__30875\,
            I => \N__30870\
        );

    \I__4712\ : LocalMux
    port map (
            O => \N__30870\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_9
        );

    \I__4711\ : InMux
    port map (
            O => \N__30867\,
            I => \N__30863\
        );

    \I__4710\ : InMux
    port map (
            O => \N__30866\,
            I => \N__30860\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__30863\,
            I => \N__30857\
        );

    \I__4708\ : LocalMux
    port map (
            O => \N__30860\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_22
        );

    \I__4707\ : Odrv12
    port map (
            O => \N__30857\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_22
        );

    \I__4706\ : CascadeMux
    port map (
            O => \N__30852\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_13_cascade_\
        );

    \I__4705\ : CascadeMux
    port map (
            O => \N__30849\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GHZ0Z5_cascade_\
        );

    \I__4704\ : InMux
    port map (
            O => \N__30846\,
            I => \N__30843\
        );

    \I__4703\ : LocalMux
    port map (
            O => \N__30843\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13\
        );

    \I__4702\ : CascadeMux
    port map (
            O => \N__30840\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13_cascade_\
        );

    \I__4701\ : InMux
    port map (
            O => \N__30837\,
            I => \N__30834\
        );

    \I__4700\ : LocalMux
    port map (
            O => \N__30834\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3QZ0Z5\
        );

    \I__4699\ : InMux
    port map (
            O => \N__30831\,
            I => \N__30828\
        );

    \I__4698\ : LocalMux
    port map (
            O => \N__30828\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4\
        );

    \I__4697\ : CascadeMux
    port map (
            O => \N__30825\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4_cascade_\
        );

    \I__4696\ : InMux
    port map (
            O => \N__30822\,
            I => \N__30819\
        );

    \I__4695\ : LocalMux
    port map (
            O => \N__30819\,
            I => \N__30816\
        );

    \I__4694\ : Odrv4
    port map (
            O => \N__30816\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_4\
        );

    \I__4693\ : InMux
    port map (
            O => \N__30813\,
            I => \N__30810\
        );

    \I__4692\ : LocalMux
    port map (
            O => \N__30810\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_13\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__30807\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_3_cascade_\
        );

    \I__4690\ : InMux
    port map (
            O => \N__30804\,
            I => \N__30801\
        );

    \I__4689\ : LocalMux
    port map (
            O => \N__30801\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_17\
        );

    \I__4688\ : CascadeMux
    port map (
            O => \N__30798\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_18_cascade_\
        );

    \I__4687\ : CascadeMux
    port map (
            O => \N__30795\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_18_cascade_\
        );

    \I__4686\ : InMux
    port map (
            O => \N__30792\,
            I => \N__30789\
        );

    \I__4685\ : LocalMux
    port map (
            O => \N__30789\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_18\
        );

    \I__4684\ : InMux
    port map (
            O => \N__30786\,
            I => \N__30783\
        );

    \I__4683\ : LocalMux
    port map (
            O => \N__30783\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_18\
        );

    \I__4682\ : InMux
    port map (
            O => \N__30780\,
            I => \N__30777\
        );

    \I__4681\ : LocalMux
    port map (
            O => \N__30777\,
            I => \N__30774\
        );

    \I__4680\ : Odrv4
    port map (
            O => \N__30774\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_13\
        );

    \I__4679\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30768\
        );

    \I__4678\ : LocalMux
    port map (
            O => \N__30768\,
            I => \N__30765\
        );

    \I__4677\ : Span4Mux_v
    port map (
            O => \N__30765\,
            I => \N__30762\
        );

    \I__4676\ : Odrv4
    port map (
            O => \N__30762\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_14\
        );

    \I__4675\ : InMux
    port map (
            O => \N__30759\,
            I => \N__30756\
        );

    \I__4674\ : LocalMux
    port map (
            O => \N__30756\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_15\
        );

    \I__4673\ : SRMux
    port map (
            O => \N__30753\,
            I => \N__30750\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__30750\,
            I => \N__30747\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__30747\,
            I => \I2C_top_level_inst1.I2C_Control_StartUp_inst.rst_neg_i\
        );

    \I__4670\ : InMux
    port map (
            O => \N__30744\,
            I => \N__30741\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__30741\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_22\
        );

    \I__4668\ : InMux
    port map (
            O => \N__30738\,
            I => \N__30735\
        );

    \I__4667\ : LocalMux
    port map (
            O => \N__30735\,
            I => \N__30732\
        );

    \I__4666\ : Span4Mux_h
    port map (
            O => \N__30732\,
            I => \N__30729\
        );

    \I__4665\ : Span4Mux_v
    port map (
            O => \N__30729\,
            I => \N__30726\
        );

    \I__4664\ : Span4Mux_h
    port map (
            O => \N__30726\,
            I => \N__30723\
        );

    \I__4663\ : Odrv4
    port map (
            O => \N__30723\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_2
        );

    \I__4662\ : InMux
    port map (
            O => \N__30720\,
            I => \N__30717\
        );

    \I__4661\ : LocalMux
    port map (
            O => \N__30717\,
            I => \N__30714\
        );

    \I__4660\ : Span12Mux_v
    port map (
            O => \N__30714\,
            I => \N__30711\
        );

    \I__4659\ : Odrv12
    port map (
            O => \N__30711\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_13
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__30708\,
            I => \N__30705\
        );

    \I__4657\ : InMux
    port map (
            O => \N__30705\,
            I => \N__30702\
        );

    \I__4656\ : LocalMux
    port map (
            O => \N__30702\,
            I => \N__30699\
        );

    \I__4655\ : Span4Mux_h
    port map (
            O => \N__30699\,
            I => \N__30696\
        );

    \I__4654\ : Span4Mux_v
    port map (
            O => \N__30696\,
            I => \N__30693\
        );

    \I__4653\ : Odrv4
    port map (
            O => \N__30693\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_13
        );

    \I__4652\ : CascadeMux
    port map (
            O => \N__30690\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_13_cascade_\
        );

    \I__4651\ : InMux
    port map (
            O => \N__30687\,
            I => \N__30684\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__30684\,
            I => \N__30681\
        );

    \I__4649\ : Span4Mux_h
    port map (
            O => \N__30681\,
            I => \N__30678\
        );

    \I__4648\ : Span4Mux_h
    port map (
            O => \N__30678\,
            I => \N__30675\
        );

    \I__4647\ : Odrv4
    port map (
            O => \N__30675\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_13
        );

    \I__4646\ : InMux
    port map (
            O => \N__30672\,
            I => \N__30669\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__30669\,
            I => \N__30666\
        );

    \I__4644\ : Span4Mux_v
    port map (
            O => \N__30666\,
            I => \N__30663\
        );

    \I__4643\ : Span4Mux_v
    port map (
            O => \N__30663\,
            I => \N__30660\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__30660\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_797\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__30657\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_13_cascade_\
        );

    \I__4640\ : InMux
    port map (
            O => \N__30654\,
            I => \N__30651\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__30651\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_13\
        );

    \I__4638\ : CascadeMux
    port map (
            O => \N__30648\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_13_cascade_\
        );

    \I__4637\ : InMux
    port map (
            O => \N__30645\,
            I => \N__30642\
        );

    \I__4636\ : LocalMux
    port map (
            O => \N__30642\,
            I => \N__30639\
        );

    \I__4635\ : Span4Mux_h
    port map (
            O => \N__30639\,
            I => \N__30636\
        );

    \I__4634\ : Span4Mux_h
    port map (
            O => \N__30636\,
            I => \N__30633\
        );

    \I__4633\ : Odrv4
    port map (
            O => \N__30633\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_18
        );

    \I__4632\ : CascadeMux
    port map (
            O => \N__30630\,
            I => \N__30627\
        );

    \I__4631\ : InMux
    port map (
            O => \N__30627\,
            I => \N__30624\
        );

    \I__4630\ : LocalMux
    port map (
            O => \N__30624\,
            I => \N__30621\
        );

    \I__4629\ : Span4Mux_h
    port map (
            O => \N__30621\,
            I => \N__30618\
        );

    \I__4628\ : Span4Mux_h
    port map (
            O => \N__30618\,
            I => \N__30615\
        );

    \I__4627\ : Span4Mux_h
    port map (
            O => \N__30615\,
            I => \N__30612\
        );

    \I__4626\ : Odrv4
    port map (
            O => \N__30612\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_18
        );

    \I__4625\ : InMux
    port map (
            O => \N__30609\,
            I => \N__30603\
        );

    \I__4624\ : InMux
    port map (
            O => \N__30608\,
            I => \N__30603\
        );

    \I__4623\ : LocalMux
    port map (
            O => \N__30603\,
            I => \N__30600\
        );

    \I__4622\ : Odrv4
    port map (
            O => \N__30600\,
            I => \cemf_module_64ch_ctrl_inst1.N_410_0\
        );

    \I__4621\ : CascadeMux
    port map (
            O => \N__30597\,
            I => \N__30592\
        );

    \I__4620\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30589\
        );

    \I__4619\ : InMux
    port map (
            O => \N__30595\,
            I => \N__30584\
        );

    \I__4618\ : InMux
    port map (
            O => \N__30592\,
            I => \N__30584\
        );

    \I__4617\ : LocalMux
    port map (
            O => \N__30589\,
            I => \N__30581\
        );

    \I__4616\ : LocalMux
    port map (
            O => \N__30584\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_7\
        );

    \I__4615\ : Odrv4
    port map (
            O => \N__30581\,
            I => \cemf_module_64ch_ctrl_inst1.c_state_7\
        );

    \I__4614\ : InMux
    port map (
            O => \N__30576\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0\
        );

    \I__4613\ : InMux
    port map (
            O => \N__30573\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1\
        );

    \I__4612\ : InMux
    port map (
            O => \N__30570\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_2\
        );

    \I__4611\ : InMux
    port map (
            O => \N__30567\,
            I => \N__30564\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__30564\,
            I => \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetterZ0\
        );

    \I__4609\ : CascadeMux
    port map (
            O => \N__30561\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1_cascade_\
        );

    \I__4608\ : InMux
    port map (
            O => \N__30558\,
            I => \N__30549\
        );

    \I__4607\ : InMux
    port map (
            O => \N__30557\,
            I => \N__30549\
        );

    \I__4606\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30542\
        );

    \I__4605\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30542\
        );

    \I__4604\ : InMux
    port map (
            O => \N__30554\,
            I => \N__30542\
        );

    \I__4603\ : LocalMux
    port map (
            O => \N__30549\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4\
        );

    \I__4602\ : LocalMux
    port map (
            O => \N__30542\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4\
        );

    \I__4601\ : InMux
    port map (
            O => \N__30537\,
            I => \N__30534\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__30534\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1\
        );

    \I__4599\ : CascadeMux
    port map (
            O => \N__30531\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_2_cascade_\
        );

    \I__4598\ : CascadeMux
    port map (
            O => \N__30528\,
            I => \N__30525\
        );

    \I__4597\ : InMux
    port map (
            O => \N__30525\,
            I => \N__30522\
        );

    \I__4596\ : LocalMux
    port map (
            O => \N__30522\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_9\
        );

    \I__4595\ : InMux
    port map (
            O => \N__30519\,
            I => \N__30516\
        );

    \I__4594\ : LocalMux
    port map (
            O => \N__30516\,
            I => \N__30510\
        );

    \I__4593\ : InMux
    port map (
            O => \N__30515\,
            I => \N__30507\
        );

    \I__4592\ : InMux
    port map (
            O => \N__30514\,
            I => \N__30504\
        );

    \I__4591\ : InMux
    port map (
            O => \N__30513\,
            I => \N__30501\
        );

    \I__4590\ : Span4Mux_v
    port map (
            O => \N__30510\,
            I => \N__30498\
        );

    \I__4589\ : LocalMux
    port map (
            O => \N__30507\,
            I => \N__30495\
        );

    \I__4588\ : LocalMux
    port map (
            O => \N__30504\,
            I => \N__30492\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__30501\,
            I => \N__30489\
        );

    \I__4586\ : Span4Mux_h
    port map (
            O => \N__30498\,
            I => \N__30484\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__30495\,
            I => \N__30484\
        );

    \I__4584\ : Odrv4
    port map (
            O => \N__30492\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__30489\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9\
        );

    \I__4582\ : Odrv4
    port map (
            O => \N__30484\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9\
        );

    \I__4581\ : InMux
    port map (
            O => \N__30477\,
            I => \N__30464\
        );

    \I__4580\ : InMux
    port map (
            O => \N__30476\,
            I => \N__30464\
        );

    \I__4579\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30464\
        );

    \I__4578\ : CascadeMux
    port map (
            O => \N__30474\,
            I => \N__30455\
        );

    \I__4577\ : InMux
    port map (
            O => \N__30473\,
            I => \N__30452\
        );

    \I__4576\ : InMux
    port map (
            O => \N__30472\,
            I => \N__30449\
        );

    \I__4575\ : CascadeMux
    port map (
            O => \N__30471\,
            I => \N__30446\
        );

    \I__4574\ : LocalMux
    port map (
            O => \N__30464\,
            I => \N__30443\
        );

    \I__4573\ : InMux
    port map (
            O => \N__30463\,
            I => \N__30430\
        );

    \I__4572\ : InMux
    port map (
            O => \N__30462\,
            I => \N__30430\
        );

    \I__4571\ : InMux
    port map (
            O => \N__30461\,
            I => \N__30430\
        );

    \I__4570\ : InMux
    port map (
            O => \N__30460\,
            I => \N__30430\
        );

    \I__4569\ : InMux
    port map (
            O => \N__30459\,
            I => \N__30430\
        );

    \I__4568\ : InMux
    port map (
            O => \N__30458\,
            I => \N__30430\
        );

    \I__4567\ : InMux
    port map (
            O => \N__30455\,
            I => \N__30427\
        );

    \I__4566\ : LocalMux
    port map (
            O => \N__30452\,
            I => \N__30424\
        );

    \I__4565\ : LocalMux
    port map (
            O => \N__30449\,
            I => \N__30421\
        );

    \I__4564\ : InMux
    port map (
            O => \N__30446\,
            I => \N__30418\
        );

    \I__4563\ : Span4Mux_v
    port map (
            O => \N__30443\,
            I => \N__30413\
        );

    \I__4562\ : LocalMux
    port map (
            O => \N__30430\,
            I => \N__30413\
        );

    \I__4561\ : LocalMux
    port map (
            O => \N__30427\,
            I => \N__30410\
        );

    \I__4560\ : Span4Mux_v
    port map (
            O => \N__30424\,
            I => \N__30405\
        );

    \I__4559\ : Span4Mux_v
    port map (
            O => \N__30421\,
            I => \N__30405\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__30418\,
            I => \N__30402\
        );

    \I__4557\ : Span4Mux_h
    port map (
            O => \N__30413\,
            I => \N__30397\
        );

    \I__4556\ : Span4Mux_v
    port map (
            O => \N__30410\,
            I => \N__30397\
        );

    \I__4555\ : Span4Mux_h
    port map (
            O => \N__30405\,
            I => \N__30394\
        );

    \I__4554\ : Span4Mux_h
    port map (
            O => \N__30402\,
            I => \N__30391\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__30397\,
            I => \N__30388\
        );

    \I__4552\ : Odrv4
    port map (
            O => \N__30394\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10\
        );

    \I__4551\ : Odrv4
    port map (
            O => \N__30391\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10\
        );

    \I__4550\ : Odrv4
    port map (
            O => \N__30388\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10\
        );

    \I__4549\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30374\
        );

    \I__4548\ : InMux
    port map (
            O => \N__30380\,
            I => \N__30374\
        );

    \I__4547\ : InMux
    port map (
            O => \N__30379\,
            I => \N__30371\
        );

    \I__4546\ : LocalMux
    port map (
            O => \N__30374\,
            I => \N__30368\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__30371\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9\
        );

    \I__4544\ : Odrv4
    port map (
            O => \N__30368\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9\
        );

    \I__4543\ : InMux
    port map (
            O => \N__30363\,
            I => \N__30360\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__30360\,
            I => \N__30357\
        );

    \I__4541\ : Odrv4
    port map (
            O => \N__30357\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_10\
        );

    \I__4540\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30351\
        );

    \I__4539\ : LocalMux
    port map (
            O => \N__30351\,
            I => \N__30346\
        );

    \I__4538\ : InMux
    port map (
            O => \N__30350\,
            I => \N__30341\
        );

    \I__4537\ : InMux
    port map (
            O => \N__30349\,
            I => \N__30341\
        );

    \I__4536\ : Odrv12
    port map (
            O => \N__30346\,
            I => \cemf_module_64ch_ctrl_inst1.N_68_0\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__30341\,
            I => \cemf_module_64ch_ctrl_inst1.N_68_0\
        );

    \I__4534\ : InMux
    port map (
            O => \N__30336\,
            I => \N__30332\
        );

    \I__4533\ : InMux
    port map (
            O => \N__30335\,
            I => \N__30329\
        );

    \I__4532\ : LocalMux
    port map (
            O => \N__30332\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4\
        );

    \I__4531\ : LocalMux
    port map (
            O => \N__30329\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4\
        );

    \I__4530\ : InMux
    port map (
            O => \N__30324\,
            I => \N__30320\
        );

    \I__4529\ : InMux
    port map (
            O => \N__30323\,
            I => \N__30317\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__30320\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3\
        );

    \I__4527\ : LocalMux
    port map (
            O => \N__30317\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3\
        );

    \I__4526\ : InMux
    port map (
            O => \N__30312\,
            I => \N__30308\
        );

    \I__4525\ : InMux
    port map (
            O => \N__30311\,
            I => \N__30305\
        );

    \I__4524\ : LocalMux
    port map (
            O => \N__30308\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2\
        );

    \I__4523\ : LocalMux
    port map (
            O => \N__30305\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2\
        );

    \I__4522\ : InMux
    port map (
            O => \N__30300\,
            I => \N__30296\
        );

    \I__4521\ : InMux
    port map (
            O => \N__30299\,
            I => \N__30293\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__30296\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1\
        );

    \I__4519\ : LocalMux
    port map (
            O => \N__30293\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1\
        );

    \I__4518\ : CascadeMux
    port map (
            O => \N__30288\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ns_i_a2_1_1_3_cascade_\
        );

    \I__4517\ : InMux
    port map (
            O => \N__30285\,
            I => \N__30281\
        );

    \I__4516\ : InMux
    port map (
            O => \N__30284\,
            I => \N__30278\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__30281\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__30278\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0\
        );

    \I__4513\ : CascadeMux
    port map (
            O => \N__30273\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987_cascade_\
        );

    \I__4512\ : InMux
    port map (
            O => \N__30270\,
            I => \N__30267\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__30267\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_2\
        );

    \I__4510\ : CascadeMux
    port map (
            O => \N__30264\,
            I => \N__30261\
        );

    \I__4509\ : InMux
    port map (
            O => \N__30261\,
            I => \N__30256\
        );

    \I__4508\ : InMux
    port map (
            O => \N__30260\,
            I => \N__30251\
        );

    \I__4507\ : InMux
    port map (
            O => \N__30259\,
            I => \N__30251\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__30256\,
            I => \N__30246\
        );

    \I__4505\ : LocalMux
    port map (
            O => \N__30251\,
            I => \N__30246\
        );

    \I__4504\ : Odrv4
    port map (
            O => \N__30246\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_0\
        );

    \I__4503\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30239\
        );

    \I__4502\ : InMux
    port map (
            O => \N__30242\,
            I => \N__30235\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__30239\,
            I => \N__30232\
        );

    \I__4500\ : InMux
    port map (
            O => \N__30238\,
            I => \N__30229\
        );

    \I__4499\ : LocalMux
    port map (
            O => \N__30235\,
            I => \N__30226\
        );

    \I__4498\ : Odrv12
    port map (
            O => \N__30232\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__30229\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291\
        );

    \I__4496\ : Odrv4
    port map (
            O => \N__30226\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291\
        );

    \I__4495\ : InMux
    port map (
            O => \N__30219\,
            I => \N__30216\
        );

    \I__4494\ : LocalMux
    port map (
            O => \N__30216\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_5\
        );

    \I__4493\ : CascadeMux
    port map (
            O => \N__30213\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_o3_i_a2_1_1_cascade_\
        );

    \I__4492\ : InMux
    port map (
            O => \N__30210\,
            I => \N__30207\
        );

    \I__4491\ : LocalMux
    port map (
            O => \N__30207\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_6\
        );

    \I__4490\ : InMux
    port map (
            O => \N__30204\,
            I => \N__30195\
        );

    \I__4489\ : InMux
    port map (
            O => \N__30203\,
            I => \N__30195\
        );

    \I__4488\ : InMux
    port map (
            O => \N__30202\,
            I => \N__30195\
        );

    \I__4487\ : LocalMux
    port map (
            O => \N__30195\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_5\
        );

    \I__4486\ : InMux
    port map (
            O => \N__30192\,
            I => \N__30189\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__30189\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_10\
        );

    \I__4484\ : InMux
    port map (
            O => \N__30186\,
            I => \N__30183\
        );

    \I__4483\ : LocalMux
    port map (
            O => \N__30183\,
            I => \N__30180\
        );

    \I__4482\ : Span12Mux_v
    port map (
            O => \N__30180\,
            I => \N__30177\
        );

    \I__4481\ : Odrv12
    port map (
            O => \N__30177\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_4
        );

    \I__4480\ : InMux
    port map (
            O => \N__30174\,
            I => \N__30171\
        );

    \I__4479\ : LocalMux
    port map (
            O => \N__30171\,
            I => \N__30168\
        );

    \I__4478\ : Span4Mux_h
    port map (
            O => \N__30168\,
            I => \N__30165\
        );

    \I__4477\ : Odrv4
    port map (
            O => \N__30165\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_896\
        );

    \I__4476\ : CascadeMux
    port map (
            O => \N__30162\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_291_reti_cascade_\
        );

    \I__4475\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30156\
        );

    \I__4474\ : LocalMux
    port map (
            O => \N__30156\,
            I => \N__30153\
        );

    \I__4473\ : Odrv4
    port map (
            O => \N__30153\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_276i\
        );

    \I__4472\ : InMux
    port map (
            O => \N__30150\,
            I => \N__30147\
        );

    \I__4471\ : LocalMux
    port map (
            O => \N__30147\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_retZ0Z_4\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__30144\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_4_0_cascade_\
        );

    \I__4469\ : InMux
    port map (
            O => \N__30141\,
            I => \N__30138\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__30138\,
            I => \N__30134\
        );

    \I__4467\ : InMux
    port map (
            O => \N__30137\,
            I => \N__30131\
        );

    \I__4466\ : Span4Mux_h
    port map (
            O => \N__30134\,
            I => \N__30128\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__30131\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283\
        );

    \I__4464\ : Odrv4
    port map (
            O => \N__30128\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283\
        );

    \I__4463\ : InMux
    port map (
            O => \N__30123\,
            I => \N__30118\
        );

    \I__4462\ : CascadeMux
    port map (
            O => \N__30122\,
            I => \N__30115\
        );

    \I__4461\ : InMux
    port map (
            O => \N__30121\,
            I => \N__30112\
        );

    \I__4460\ : LocalMux
    port map (
            O => \N__30118\,
            I => \N__30109\
        );

    \I__4459\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30106\
        );

    \I__4458\ : LocalMux
    port map (
            O => \N__30112\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10\
        );

    \I__4457\ : Odrv4
    port map (
            O => \N__30109\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__30106\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10\
        );

    \I__4455\ : CascadeMux
    port map (
            O => \N__30099\,
            I => \N__30096\
        );

    \I__4454\ : InMux
    port map (
            O => \N__30096\,
            I => \N__30093\
        );

    \I__4453\ : LocalMux
    port map (
            O => \N__30093\,
            I => \N__30090\
        );

    \I__4452\ : Span4Mux_h
    port map (
            O => \N__30090\,
            I => \N__30087\
        );

    \I__4451\ : Odrv4
    port map (
            O => \N__30087\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__30084\,
            I => \N__30078\
        );

    \I__4449\ : InMux
    port map (
            O => \N__30083\,
            I => \N__30074\
        );

    \I__4448\ : InMux
    port map (
            O => \N__30082\,
            I => \N__30071\
        );

    \I__4447\ : InMux
    port map (
            O => \N__30081\,
            I => \N__30068\
        );

    \I__4446\ : InMux
    port map (
            O => \N__30078\,
            I => \N__30063\
        );

    \I__4445\ : InMux
    port map (
            O => \N__30077\,
            I => \N__30063\
        );

    \I__4444\ : LocalMux
    port map (
            O => \N__30074\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__30071\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__30068\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11\
        );

    \I__4441\ : LocalMux
    port map (
            O => \N__30063\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11\
        );

    \I__4440\ : CascadeMux
    port map (
            O => \N__30054\,
            I => \N__30049\
        );

    \I__4439\ : InMux
    port map (
            O => \N__30053\,
            I => \N__30046\
        );

    \I__4438\ : InMux
    port map (
            O => \N__30052\,
            I => \N__30041\
        );

    \I__4437\ : InMux
    port map (
            O => \N__30049\,
            I => \N__30041\
        );

    \I__4436\ : LocalMux
    port map (
            O => \N__30046\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__30041\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14\
        );

    \I__4434\ : InMux
    port map (
            O => \N__30036\,
            I => \N__30030\
        );

    \I__4433\ : CascadeMux
    port map (
            O => \N__30035\,
            I => \N__30027\
        );

    \I__4432\ : InMux
    port map (
            O => \N__30034\,
            I => \N__30023\
        );

    \I__4431\ : InMux
    port map (
            O => \N__30033\,
            I => \N__30020\
        );

    \I__4430\ : LocalMux
    port map (
            O => \N__30030\,
            I => \N__30017\
        );

    \I__4429\ : InMux
    port map (
            O => \N__30027\,
            I => \N__30012\
        );

    \I__4428\ : InMux
    port map (
            O => \N__30026\,
            I => \N__30012\
        );

    \I__4427\ : LocalMux
    port map (
            O => \N__30023\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15\
        );

    \I__4426\ : LocalMux
    port map (
            O => \N__30020\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15\
        );

    \I__4425\ : Odrv4
    port map (
            O => \N__30017\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15\
        );

    \I__4424\ : LocalMux
    port map (
            O => \N__30012\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15\
        );

    \I__4423\ : CascadeMux
    port map (
            O => \N__30003\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_2_0_cascade_\
        );

    \I__4422\ : InMux
    port map (
            O => \N__30000\,
            I => \N__29996\
        );

    \I__4421\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29993\
        );

    \I__4420\ : LocalMux
    port map (
            O => \N__29996\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286\
        );

    \I__4419\ : LocalMux
    port map (
            O => \N__29993\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286\
        );

    \I__4418\ : CascadeMux
    port map (
            O => \N__29988\,
            I => \N__29983\
        );

    \I__4417\ : InMux
    port map (
            O => \N__29987\,
            I => \N__29976\
        );

    \I__4416\ : InMux
    port map (
            O => \N__29986\,
            I => \N__29976\
        );

    \I__4415\ : InMux
    port map (
            O => \N__29983\,
            I => \N__29976\
        );

    \I__4414\ : LocalMux
    port map (
            O => \N__29976\,
            I => \N__29973\
        );

    \I__4413\ : Odrv4
    port map (
            O => \N__29973\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_0_0\
        );

    \I__4412\ : CascadeMux
    port map (
            O => \N__29970\,
            I => \N__29965\
        );

    \I__4411\ : CascadeMux
    port map (
            O => \N__29969\,
            I => \N__29962\
        );

    \I__4410\ : CascadeMux
    port map (
            O => \N__29968\,
            I => \N__29959\
        );

    \I__4409\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29952\
        );

    \I__4408\ : InMux
    port map (
            O => \N__29962\,
            I => \N__29952\
        );

    \I__4407\ : InMux
    port map (
            O => \N__29959\,
            I => \N__29943\
        );

    \I__4406\ : InMux
    port map (
            O => \N__29958\,
            I => \N__29943\
        );

    \I__4405\ : InMux
    port map (
            O => \N__29957\,
            I => \N__29943\
        );

    \I__4404\ : LocalMux
    port map (
            O => \N__29952\,
            I => \N__29937\
        );

    \I__4403\ : InMux
    port map (
            O => \N__29951\,
            I => \N__29932\
        );

    \I__4402\ : InMux
    port map (
            O => \N__29950\,
            I => \N__29932\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__29943\,
            I => \N__29929\
        );

    \I__4400\ : InMux
    port map (
            O => \N__29942\,
            I => \N__29924\
        );

    \I__4399\ : InMux
    port map (
            O => \N__29941\,
            I => \N__29924\
        );

    \I__4398\ : CascadeMux
    port map (
            O => \N__29940\,
            I => \N__29921\
        );

    \I__4397\ : Span4Mux_v
    port map (
            O => \N__29937\,
            I => \N__29913\
        );

    \I__4396\ : LocalMux
    port map (
            O => \N__29932\,
            I => \N__29913\
        );

    \I__4395\ : Span4Mux_v
    port map (
            O => \N__29929\,
            I => \N__29913\
        );

    \I__4394\ : LocalMux
    port map (
            O => \N__29924\,
            I => \N__29910\
        );

    \I__4393\ : InMux
    port map (
            O => \N__29921\,
            I => \N__29905\
        );

    \I__4392\ : InMux
    port map (
            O => \N__29920\,
            I => \N__29905\
        );

    \I__4391\ : Span4Mux_h
    port map (
            O => \N__29913\,
            I => \N__29900\
        );

    \I__4390\ : Span4Mux_v
    port map (
            O => \N__29910\,
            I => \N__29900\
        );

    \I__4389\ : LocalMux
    port map (
            O => \N__29905\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0\
        );

    \I__4388\ : Odrv4
    port map (
            O => \N__29900\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0\
        );

    \I__4387\ : CascadeMux
    port map (
            O => \N__29895\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_6_cascade_\
        );

    \I__4386\ : CascadeMux
    port map (
            O => \N__29892\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3QZ0Z5_cascade_\
        );

    \I__4385\ : InMux
    port map (
            O => \N__29889\,
            I => \N__29885\
        );

    \I__4384\ : InMux
    port map (
            O => \N__29888\,
            I => \N__29882\
        );

    \I__4383\ : LocalMux
    port map (
            O => \N__29885\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6\
        );

    \I__4382\ : LocalMux
    port map (
            O => \N__29882\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6\
        );

    \I__4381\ : InMux
    port map (
            O => \N__29877\,
            I => \N__29874\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__29874\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3QZ0Z5\
        );

    \I__4379\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29868\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__29868\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5\
        );

    \I__4377\ : CascadeMux
    port map (
            O => \N__29865\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5_cascade_\
        );

    \I__4376\ : InMux
    port map (
            O => \N__29862\,
            I => \N__29859\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__29859\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_5\
        );

    \I__4374\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29852\
        );

    \I__4373\ : InMux
    port map (
            O => \N__29855\,
            I => \N__29849\
        );

    \I__4372\ : LocalMux
    port map (
            O => \N__29852\,
            I => \N__29846\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__29849\,
            I => \cemf_module_64ch_ctrl_inst1.N_1615\
        );

    \I__4370\ : Odrv12
    port map (
            O => \N__29846\,
            I => \cemf_module_64ch_ctrl_inst1.N_1615\
        );

    \I__4369\ : CascadeMux
    port map (
            O => \N__29841\,
            I => \N_1614_cascade_\
        );

    \I__4368\ : InMux
    port map (
            O => \N__29838\,
            I => \N__29835\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29832\
        );

    \I__4366\ : Span4Mux_v
    port map (
            O => \N__29832\,
            I => \N__29829\
        );

    \I__4365\ : Span4Mux_h
    port map (
            O => \N__29829\,
            I => \N__29826\
        );

    \I__4364\ : Odrv4
    port map (
            O => \N__29826\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_28
        );

    \I__4363\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29820\
        );

    \I__4362\ : LocalMux
    port map (
            O => \N__29820\,
            I => \N__29817\
        );

    \I__4361\ : Odrv12
    port map (
            O => \N__29817\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_643\
        );

    \I__4360\ : InMux
    port map (
            O => \N__29814\,
            I => \N__29811\
        );

    \I__4359\ : LocalMux
    port map (
            O => \N__29811\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_5\
        );

    \I__4358\ : InMux
    port map (
            O => \N__29808\,
            I => \N__29805\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__29805\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_6\
        );

    \I__4356\ : InMux
    port map (
            O => \N__29802\,
            I => \N__29799\
        );

    \I__4355\ : LocalMux
    port map (
            O => \N__29799\,
            I => \N__29796\
        );

    \I__4354\ : Span4Mux_v
    port map (
            O => \N__29796\,
            I => \N__29793\
        );

    \I__4353\ : Span4Mux_h
    port map (
            O => \N__29793\,
            I => \N__29790\
        );

    \I__4352\ : Span4Mux_v
    port map (
            O => \N__29790\,
            I => \N__29787\
        );

    \I__4351\ : Span4Mux_v
    port map (
            O => \N__29787\,
            I => \N__29784\
        );

    \I__4350\ : Odrv4
    port map (
            O => \N__29784\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_6
        );

    \I__4349\ : CascadeMux
    port map (
            O => \N__29781\,
            I => \N__29778\
        );

    \I__4348\ : InMux
    port map (
            O => \N__29778\,
            I => \N__29775\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29772\
        );

    \I__4346\ : Span4Mux_v
    port map (
            O => \N__29772\,
            I => \N__29769\
        );

    \I__4345\ : Span4Mux_v
    port map (
            O => \N__29769\,
            I => \N__29766\
        );

    \I__4344\ : Span4Mux_h
    port map (
            O => \N__29766\,
            I => \N__29763\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__29763\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_6
        );

    \I__4342\ : InMux
    port map (
            O => \N__29760\,
            I => \N__29757\
        );

    \I__4341\ : LocalMux
    port map (
            O => \N__29757\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_6\
        );

    \I__4340\ : InMux
    port map (
            O => \N__29754\,
            I => \N__29751\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__29751\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_9\
        );

    \I__4338\ : CascadeMux
    port map (
            O => \N__29748\,
            I => \N__29745\
        );

    \I__4337\ : InMux
    port map (
            O => \N__29745\,
            I => \N__29742\
        );

    \I__4336\ : LocalMux
    port map (
            O => \N__29742\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_841\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__29739\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_9_cascade_\
        );

    \I__4334\ : InMux
    port map (
            O => \N__29736\,
            I => \N__29733\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__29733\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_9\
        );

    \I__4332\ : InMux
    port map (
            O => \N__29730\,
            I => \N__29727\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__29727\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_9\
        );

    \I__4330\ : InMux
    port map (
            O => \N__29724\,
            I => \N__29721\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__29721\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_9\
        );

    \I__4328\ : CascadeMux
    port map (
            O => \N__29718\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_5_cascade_\
        );

    \I__4327\ : CascadeMux
    port map (
            O => \N__29715\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_4_cascade_\
        );

    \I__4326\ : InMux
    port map (
            O => \N__29712\,
            I => \N__29709\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__29709\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_4\
        );

    \I__4324\ : InMux
    port map (
            O => \N__29706\,
            I => \N__29703\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__29703\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_4\
        );

    \I__4322\ : CascadeMux
    port map (
            O => \N__29700\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_4_cascade_\
        );

    \I__4321\ : InMux
    port map (
            O => \N__29697\,
            I => \N__29694\
        );

    \I__4320\ : LocalMux
    port map (
            O => \N__29694\,
            I => \N__29691\
        );

    \I__4319\ : Span4Mux_v
    port map (
            O => \N__29691\,
            I => \N__29686\
        );

    \I__4318\ : InMux
    port map (
            O => \N__29690\,
            I => \N__29681\
        );

    \I__4317\ : InMux
    port map (
            O => \N__29689\,
            I => \N__29681\
        );

    \I__4316\ : Odrv4
    port map (
            O => \N__29686\,
            I => cemf_module_64ch_ctrl_inst1_data_config_4
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__29681\,
            I => cemf_module_64ch_ctrl_inst1_data_config_4
        );

    \I__4314\ : CascadeMux
    port map (
            O => \N__29676\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRLZ0Z7_cascade_\
        );

    \I__4313\ : CascadeMux
    port map (
            O => \N__29673\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_6_cascade_\
        );

    \I__4312\ : InMux
    port map (
            O => \N__29670\,
            I => \N__29667\
        );

    \I__4311\ : LocalMux
    port map (
            O => \N__29667\,
            I => \N__29664\
        );

    \I__4310\ : Odrv12
    port map (
            O => \N__29664\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_6\
        );

    \I__4309\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29658\
        );

    \I__4308\ : LocalMux
    port map (
            O => \N__29658\,
            I => \N__29655\
        );

    \I__4307\ : Span4Mux_v
    port map (
            O => \N__29655\,
            I => \N__29652\
        );

    \I__4306\ : Odrv4
    port map (
            O => \N__29652\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_775\
        );

    \I__4305\ : CascadeMux
    port map (
            O => \N__29649\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_15_cascade_\
        );

    \I__4304\ : CascadeMux
    port map (
            O => \N__29646\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_15_cascade_\
        );

    \I__4303\ : InMux
    port map (
            O => \N__29643\,
            I => \N__29640\
        );

    \I__4302\ : LocalMux
    port map (
            O => \N__29640\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_15\
        );

    \I__4301\ : InMux
    port map (
            O => \N__29637\,
            I => \N__29634\
        );

    \I__4300\ : LocalMux
    port map (
            O => \N__29634\,
            I => \N__29631\
        );

    \I__4299\ : Span4Mux_v
    port map (
            O => \N__29631\,
            I => \N__29628\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__29628\,
            I => \N__29625\
        );

    \I__4297\ : Odrv4
    port map (
            O => \N__29625\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_23
        );

    \I__4296\ : InMux
    port map (
            O => \N__29622\,
            I => \N__29619\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__29619\,
            I => \N__29616\
        );

    \I__4294\ : Span4Mux_h
    port map (
            O => \N__29616\,
            I => \N__29613\
        );

    \I__4293\ : Span4Mux_h
    port map (
            O => \N__29613\,
            I => \N__29610\
        );

    \I__4292\ : Span4Mux_v
    port map (
            O => \N__29610\,
            I => \N__29607\
        );

    \I__4291\ : Odrv4
    port map (
            O => \N__29607\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_17
        );

    \I__4290\ : CascadeMux
    port map (
            O => \N__29604\,
            I => \N__29601\
        );

    \I__4289\ : InMux
    port map (
            O => \N__29601\,
            I => \N__29598\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__29598\,
            I => \N__29595\
        );

    \I__4287\ : Span4Mux_v
    port map (
            O => \N__29595\,
            I => \N__29592\
        );

    \I__4286\ : Sp12to4
    port map (
            O => \N__29592\,
            I => \N__29589\
        );

    \I__4285\ : Odrv12
    port map (
            O => \N__29589\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_17
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__29586\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_17_cascade_\
        );

    \I__4283\ : InMux
    port map (
            O => \N__29583\,
            I => \N__29580\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__29580\,
            I => \N__29577\
        );

    \I__4281\ : Span4Mux_v
    port map (
            O => \N__29577\,
            I => \N__29574\
        );

    \I__4280\ : Span4Mux_h
    port map (
            O => \N__29574\,
            I => \N__29571\
        );

    \I__4279\ : Odrv4
    port map (
            O => \N__29571\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_17
        );

    \I__4278\ : CascadeMux
    port map (
            O => \N__29568\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_17_cascade_\
        );

    \I__4277\ : CascadeMux
    port map (
            O => \N__29565\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_17_cascade_\
        );

    \I__4276\ : InMux
    port map (
            O => \N__29562\,
            I => \N__29559\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__29559\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_17\
        );

    \I__4274\ : InMux
    port map (
            O => \N__29556\,
            I => \N__29553\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__29553\,
            I => \N__29550\
        );

    \I__4272\ : Span4Mux_h
    port map (
            O => \N__29550\,
            I => \N__29547\
        );

    \I__4271\ : Span4Mux_v
    port map (
            O => \N__29547\,
            I => \N__29544\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__29544\,
            I => \N__29541\
        );

    \I__4269\ : Odrv4
    port map (
            O => \N__29541\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_25
        );

    \I__4268\ : InMux
    port map (
            O => \N__29538\,
            I => \N__29535\
        );

    \I__4267\ : LocalMux
    port map (
            O => \N__29535\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_22\
        );

    \I__4266\ : InMux
    port map (
            O => \N__29532\,
            I => \N__29529\
        );

    \I__4265\ : LocalMux
    port map (
            O => \N__29529\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_22\
        );

    \I__4264\ : InMux
    port map (
            O => \N__29526\,
            I => \N__29523\
        );

    \I__4263\ : LocalMux
    port map (
            O => \N__29523\,
            I => \N__29520\
        );

    \I__4262\ : Span12Mux_v
    port map (
            O => \N__29520\,
            I => \N__29517\
        );

    \I__4261\ : Odrv12
    port map (
            O => \N__29517\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_28
        );

    \I__4260\ : CascadeMux
    port map (
            O => \N__29514\,
            I => \N__29511\
        );

    \I__4259\ : InMux
    port map (
            O => \N__29511\,
            I => \N__29508\
        );

    \I__4258\ : LocalMux
    port map (
            O => \N__29508\,
            I => \N__29505\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__29505\,
            I => \N__29502\
        );

    \I__4256\ : Span4Mux_h
    port map (
            O => \N__29502\,
            I => \N__29499\
        );

    \I__4255\ : Odrv4
    port map (
            O => \N__29499\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_28
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__29496\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_28_cascade_\
        );

    \I__4253\ : InMux
    port map (
            O => \N__29493\,
            I => \N__29490\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__29490\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_28\
        );

    \I__4251\ : CascadeMux
    port map (
            O => \N__29487\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_28_cascade_\
        );

    \I__4250\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29481\
        );

    \I__4249\ : LocalMux
    port map (
            O => \N__29481\,
            I => \N__29478\
        );

    \I__4248\ : Span4Mux_h
    port map (
            O => \N__29478\,
            I => \N__29475\
        );

    \I__4247\ : Odrv4
    port map (
            O => \N__29475\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_28\
        );

    \I__4246\ : InMux
    port map (
            O => \N__29472\,
            I => \N__29469\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__29469\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_28\
        );

    \I__4244\ : InMux
    port map (
            O => \N__29466\,
            I => \N__29463\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__29463\,
            I => \N__29460\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__29460\,
            I => \N__29457\
        );

    \I__4241\ : Span4Mux_h
    port map (
            O => \N__29457\,
            I => \N__29454\
        );

    \I__4240\ : Span4Mux_v
    port map (
            O => \N__29454\,
            I => \N__29451\
        );

    \I__4239\ : Odrv4
    port map (
            O => \N__29451\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_15
        );

    \I__4238\ : CascadeMux
    port map (
            O => \N__29448\,
            I => \N__29445\
        );

    \I__4237\ : InMux
    port map (
            O => \N__29445\,
            I => \N__29442\
        );

    \I__4236\ : LocalMux
    port map (
            O => \N__29442\,
            I => \N__29439\
        );

    \I__4235\ : Span4Mux_v
    port map (
            O => \N__29439\,
            I => \N__29436\
        );

    \I__4234\ : Span4Mux_h
    port map (
            O => \N__29436\,
            I => \N__29433\
        );

    \I__4233\ : Odrv4
    port map (
            O => \N__29433\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_15
        );

    \I__4232\ : CascadeMux
    port map (
            O => \N__29430\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_15_cascade_\
        );

    \I__4231\ : InMux
    port map (
            O => \N__29427\,
            I => \N__29424\
        );

    \I__4230\ : LocalMux
    port map (
            O => \N__29424\,
            I => \N__29421\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__29421\,
            I => \N__29418\
        );

    \I__4228\ : Span4Mux_h
    port map (
            O => \N__29418\,
            I => \N__29415\
        );

    \I__4227\ : Odrv4
    port map (
            O => \N__29415\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_15
        );

    \I__4226\ : InMux
    port map (
            O => \N__29412\,
            I => \N__29409\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__29409\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un40_0_a2_4_a2_0\
        );

    \I__4224\ : InMux
    port map (
            O => \N__29406\,
            I => \N__29402\
        );

    \I__4223\ : InMux
    port map (
            O => \N__29405\,
            I => \N__29399\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__29402\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__29399\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0\
        );

    \I__4220\ : InMux
    port map (
            O => \N__29394\,
            I => \N__29382\
        );

    \I__4219\ : InMux
    port map (
            O => \N__29393\,
            I => \N__29382\
        );

    \I__4218\ : InMux
    port map (
            O => \N__29392\,
            I => \N__29382\
        );

    \I__4217\ : InMux
    port map (
            O => \N__29391\,
            I => \N__29377\
        );

    \I__4216\ : InMux
    port map (
            O => \N__29390\,
            I => \N__29377\
        );

    \I__4215\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29374\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__29382\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17\
        );

    \I__4213\ : LocalMux
    port map (
            O => \N__29377\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17\
        );

    \I__4212\ : LocalMux
    port map (
            O => \N__29374\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17\
        );

    \I__4211\ : InMux
    port map (
            O => \N__29367\,
            I => \N__29360\
        );

    \I__4210\ : InMux
    port map (
            O => \N__29366\,
            I => \N__29353\
        );

    \I__4209\ : InMux
    port map (
            O => \N__29365\,
            I => \N__29353\
        );

    \I__4208\ : InMux
    port map (
            O => \N__29364\,
            I => \N__29353\
        );

    \I__4207\ : InMux
    port map (
            O => \N__29363\,
            I => \N__29350\
        );

    \I__4206\ : LocalMux
    port map (
            O => \N__29360\,
            I => \N__29347\
        );

    \I__4205\ : LocalMux
    port map (
            O => \N__29353\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16\
        );

    \I__4204\ : LocalMux
    port map (
            O => \N__29350\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16\
        );

    \I__4203\ : Odrv4
    port map (
            O => \N__29347\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16\
        );

    \I__4202\ : IoInMux
    port map (
            O => \N__29340\,
            I => \N__29337\
        );

    \I__4201\ : LocalMux
    port map (
            O => \N__29337\,
            I => \N__29334\
        );

    \I__4200\ : IoSpan4Mux
    port map (
            O => \N__29334\,
            I => \N__29331\
        );

    \I__4199\ : Span4Mux_s3_h
    port map (
            O => \N__29331\,
            I => \N__29328\
        );

    \I__4198\ : Span4Mux_h
    port map (
            O => \N__29328\,
            I => \N__29325\
        );

    \I__4197\ : Span4Mux_h
    port map (
            O => \N__29325\,
            I => \N__29322\
        );

    \I__4196\ : Odrv4
    port map (
            O => \N__29322\,
            I => sda_o
        );

    \I__4195\ : CascadeMux
    port map (
            O => \N__29319\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_22_cascade_\
        );

    \I__4194\ : InMux
    port map (
            O => \N__29316\,
            I => \N__29313\
        );

    \I__4193\ : LocalMux
    port map (
            O => \N__29313\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_22\
        );

    \I__4192\ : InMux
    port map (
            O => \N__29310\,
            I => \N__29307\
        );

    \I__4191\ : LocalMux
    port map (
            O => \N__29307\,
            I => \N__29304\
        );

    \I__4190\ : Span4Mux_v
    port map (
            O => \N__29304\,
            I => \N__29301\
        );

    \I__4189\ : Span4Mux_h
    port map (
            O => \N__29301\,
            I => \N__29298\
        );

    \I__4188\ : Odrv4
    port map (
            O => \N__29298\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_22
        );

    \I__4187\ : CascadeMux
    port map (
            O => \N__29295\,
            I => \N__29292\
        );

    \I__4186\ : InMux
    port map (
            O => \N__29292\,
            I => \N__29289\
        );

    \I__4185\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29286\
        );

    \I__4184\ : Span4Mux_v
    port map (
            O => \N__29286\,
            I => \N__29283\
        );

    \I__4183\ : Span4Mux_h
    port map (
            O => \N__29283\,
            I => \N__29280\
        );

    \I__4182\ : Odrv4
    port map (
            O => \N__29280\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_22
        );

    \I__4181\ : InMux
    port map (
            O => \N__29277\,
            I => \N__29274\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__29274\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_22\
        );

    \I__4179\ : InMux
    port map (
            O => \N__29271\,
            I => \bfn_12_20_0_\
        );

    \I__4178\ : InMux
    port map (
            O => \N__29268\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0\
        );

    \I__4177\ : InMux
    port map (
            O => \N__29265\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1\
        );

    \I__4176\ : InMux
    port map (
            O => \N__29262\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2\
        );

    \I__4175\ : InMux
    port map (
            O => \N__29259\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_3\
        );

    \I__4174\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29253\
        );

    \I__4173\ : LocalMux
    port map (
            O => \N__29253\,
            I => \cemf_module_64ch_ctrl_inst1.en_ch_cnt_0_a2_0_a2_1\
        );

    \I__4172\ : InMux
    port map (
            O => \N__29250\,
            I => \N__29247\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__29247\,
            I => \N__29244\
        );

    \I__4170\ : Span4Mux_h
    port map (
            O => \N__29244\,
            I => \N__29241\
        );

    \I__4169\ : Span4Mux_h
    port map (
            O => \N__29241\,
            I => \N__29238\
        );

    \I__4168\ : Odrv4
    port map (
            O => \N__29238\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1867_0\
        );

    \I__4167\ : InMux
    port map (
            O => \N__29235\,
            I => \N__29229\
        );

    \I__4166\ : InMux
    port map (
            O => \N__29234\,
            I => \N__29229\
        );

    \I__4165\ : LocalMux
    port map (
            O => \N__29229\,
            I => \N__29226\
        );

    \I__4164\ : Span4Mux_h
    port map (
            O => \N__29226\,
            I => \N__29216\
        );

    \I__4163\ : InMux
    port map (
            O => \N__29225\,
            I => \N__29209\
        );

    \I__4162\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29209\
        );

    \I__4161\ : InMux
    port map (
            O => \N__29223\,
            I => \N__29209\
        );

    \I__4160\ : InMux
    port map (
            O => \N__29222\,
            I => \N__29204\
        );

    \I__4159\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29204\
        );

    \I__4158\ : InMux
    port map (
            O => \N__29220\,
            I => \N__29199\
        );

    \I__4157\ : InMux
    port map (
            O => \N__29219\,
            I => \N__29199\
        );

    \I__4156\ : Odrv4
    port map (
            O => \N__29216\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996\
        );

    \I__4155\ : LocalMux
    port map (
            O => \N__29209\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996\
        );

    \I__4154\ : LocalMux
    port map (
            O => \N__29204\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__29199\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996\
        );

    \I__4152\ : InMux
    port map (
            O => \N__29190\,
            I => \N__29186\
        );

    \I__4151\ : InMux
    port map (
            O => \N__29189\,
            I => \N__29183\
        );

    \I__4150\ : LocalMux
    port map (
            O => \N__29186\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1\
        );

    \I__4149\ : LocalMux
    port map (
            O => \N__29183\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1\
        );

    \I__4148\ : InMux
    port map (
            O => \N__29178\,
            I => \N__29172\
        );

    \I__4147\ : InMux
    port map (
            O => \N__29177\,
            I => \N__29172\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__29172\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_13\
        );

    \I__4145\ : InMux
    port map (
            O => \N__29169\,
            I => \N__29157\
        );

    \I__4144\ : InMux
    port map (
            O => \N__29168\,
            I => \N__29157\
        );

    \I__4143\ : InMux
    port map (
            O => \N__29167\,
            I => \N__29157\
        );

    \I__4142\ : InMux
    port map (
            O => \N__29166\,
            I => \N__29157\
        );

    \I__4141\ : LocalMux
    port map (
            O => \N__29157\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_12\
        );

    \I__4140\ : InMux
    port map (
            O => \N__29154\,
            I => \N__29151\
        );

    \I__4139\ : LocalMux
    port map (
            O => \N__29151\,
            I => \N__29148\
        );

    \I__4138\ : Span4Mux_v
    port map (
            O => \N__29148\,
            I => \N__29142\
        );

    \I__4137\ : InMux
    port map (
            O => \N__29147\,
            I => \N__29135\
        );

    \I__4136\ : InMux
    port map (
            O => \N__29146\,
            I => \N__29135\
        );

    \I__4135\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29135\
        );

    \I__4134\ : Odrv4
    port map (
            O => \N__29142\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4\
        );

    \I__4133\ : LocalMux
    port map (
            O => \N__29135\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4\
        );

    \I__4132\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29126\
        );

    \I__4131\ : InMux
    port map (
            O => \N__29129\,
            I => \N__29123\
        );

    \I__4130\ : LocalMux
    port map (
            O => \N__29126\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__29123\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4\
        );

    \I__4128\ : InMux
    port map (
            O => \N__29118\,
            I => \N__29114\
        );

    \I__4127\ : InMux
    port map (
            O => \N__29117\,
            I => \N__29111\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__29114\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3\
        );

    \I__4125\ : LocalMux
    port map (
            O => \N__29111\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3\
        );

    \I__4124\ : InMux
    port map (
            O => \N__29106\,
            I => \N__29103\
        );

    \I__4123\ : LocalMux
    port map (
            O => \N__29103\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_i_a2_1_1_3\
        );

    \I__4122\ : InMux
    port map (
            O => \N__29100\,
            I => \N__29096\
        );

    \I__4121\ : InMux
    port map (
            O => \N__29099\,
            I => \N__29092\
        );

    \I__4120\ : LocalMux
    port map (
            O => \N__29096\,
            I => \N__29089\
        );

    \I__4119\ : InMux
    port map (
            O => \N__29095\,
            I => \N__29086\
        );

    \I__4118\ : LocalMux
    port map (
            O => \N__29092\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__4117\ : Odrv4
    port map (
            O => \N__29089\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__4116\ : LocalMux
    port map (
            O => \N__29086\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16\
        );

    \I__4115\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29076\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29071\
        );

    \I__4113\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29066\
        );

    \I__4112\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29066\
        );

    \I__4111\ : Odrv4
    port map (
            O => \N__29071\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__29066\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8\
        );

    \I__4109\ : InMux
    port map (
            O => \N__29061\,
            I => \N__29057\
        );

    \I__4108\ : InMux
    port map (
            O => \N__29060\,
            I => \N__29054\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__29057\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__29054\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1\
        );

    \I__4105\ : InMux
    port map (
            O => \N__29049\,
            I => \N__29045\
        );

    \I__4104\ : InMux
    port map (
            O => \N__29048\,
            I => \N__29042\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__29045\,
            I => \N__29038\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__29042\,
            I => \N__29034\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__29041\,
            I => \N__29030\
        );

    \I__4100\ : Span4Mux_h
    port map (
            O => \N__29038\,
            I => \N__29027\
        );

    \I__4099\ : InMux
    port map (
            O => \N__29037\,
            I => \N__29024\
        );

    \I__4098\ : Span4Mux_h
    port map (
            O => \N__29034\,
            I => \N__29021\
        );

    \I__4097\ : InMux
    port map (
            O => \N__29033\,
            I => \N__29016\
        );

    \I__4096\ : InMux
    port map (
            O => \N__29030\,
            I => \N__29016\
        );

    \I__4095\ : Odrv4
    port map (
            O => \N__29027\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__29024\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17\
        );

    \I__4093\ : Odrv4
    port map (
            O => \N__29021\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__29016\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17\
        );

    \I__4091\ : CascadeMux
    port map (
            O => \N__29007\,
            I => \N__29003\
        );

    \I__4090\ : CascadeMux
    port map (
            O => \N__29006\,
            I => \N__29000\
        );

    \I__4089\ : InMux
    port map (
            O => \N__29003\,
            I => \N__28996\
        );

    \I__4088\ : InMux
    port map (
            O => \N__29000\,
            I => \N__28992\
        );

    \I__4087\ : InMux
    port map (
            O => \N__28999\,
            I => \N__28989\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__28996\,
            I => \N__28986\
        );

    \I__4085\ : InMux
    port map (
            O => \N__28995\,
            I => \N__28983\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__28992\,
            I => \N__28980\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__28989\,
            I => \N__28977\
        );

    \I__4082\ : Span12Mux_v
    port map (
            O => \N__28986\,
            I => \N__28974\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__28983\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5\
        );

    \I__4080\ : Odrv4
    port map (
            O => \N__28980\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5\
        );

    \I__4079\ : Odrv4
    port map (
            O => \N__28977\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5\
        );

    \I__4078\ : Odrv12
    port map (
            O => \N__28974\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5\
        );

    \I__4077\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28962\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__28962\,
            I => \N__28959\
        );

    \I__4075\ : Span4Mux_h
    port map (
            O => \N__28959\,
            I => \N__28953\
        );

    \I__4074\ : InMux
    port map (
            O => \N__28958\,
            I => \N__28946\
        );

    \I__4073\ : InMux
    port map (
            O => \N__28957\,
            I => \N__28946\
        );

    \I__4072\ : InMux
    port map (
            O => \N__28956\,
            I => \N__28946\
        );

    \I__4071\ : Odrv4
    port map (
            O => \N__28953\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9\
        );

    \I__4070\ : LocalMux
    port map (
            O => \N__28946\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9\
        );

    \I__4069\ : InMux
    port map (
            O => \N__28941\,
            I => \N__28938\
        );

    \I__4068\ : LocalMux
    port map (
            O => \N__28938\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_18\
        );

    \I__4067\ : InMux
    port map (
            O => \N__28935\,
            I => \N__28932\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__28932\,
            I => \N__28929\
        );

    \I__4065\ : Span4Mux_v
    port map (
            O => \N__28929\,
            I => \N__28926\
        );

    \I__4064\ : Span4Mux_h
    port map (
            O => \N__28926\,
            I => \N__28923\
        );

    \I__4063\ : Odrv4
    port map (
            O => \N__28923\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_18\
        );

    \I__4062\ : CascadeMux
    port map (
            O => \N__28920\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286_cascade_\
        );

    \I__4061\ : InMux
    port map (
            O => \N__28917\,
            I => \N__28914\
        );

    \I__4060\ : LocalMux
    port map (
            O => \N__28914\,
            I => \N__28911\
        );

    \I__4059\ : Span4Mux_h
    port map (
            O => \N__28911\,
            I => \N__28905\
        );

    \I__4058\ : InMux
    port map (
            O => \N__28910\,
            I => \N__28902\
        );

    \I__4057\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28897\
        );

    \I__4056\ : InMux
    port map (
            O => \N__28908\,
            I => \N__28897\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__28905\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3\
        );

    \I__4054\ : LocalMux
    port map (
            O => \N__28902\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3\
        );

    \I__4053\ : LocalMux
    port map (
            O => \N__28897\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3\
        );

    \I__4052\ : CascadeMux
    port map (
            O => \N__28890\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15Z0Z_0_cascade_\
        );

    \I__4051\ : InMux
    port map (
            O => \N__28887\,
            I => \N__28883\
        );

    \I__4050\ : InMux
    port map (
            O => \N__28886\,
            I => \N__28880\
        );

    \I__4049\ : LocalMux
    port map (
            O => \N__28883\,
            I => \N__28875\
        );

    \I__4048\ : LocalMux
    port map (
            O => \N__28880\,
            I => \N__28875\
        );

    \I__4047\ : Span4Mux_h
    port map (
            O => \N__28875\,
            I => \N__28871\
        );

    \I__4046\ : InMux
    port map (
            O => \N__28874\,
            I => \N__28868\
        );

    \I__4045\ : Odrv4
    port map (
            O => \N__28871\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7\
        );

    \I__4044\ : LocalMux
    port map (
            O => \N__28868\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7\
        );

    \I__4043\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28858\
        );

    \I__4042\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28853\
        );

    \I__4041\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28853\
        );

    \I__4040\ : LocalMux
    port map (
            O => \N__28858\,
            I => \N__28850\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__28853\,
            I => \N__28844\
        );

    \I__4038\ : Span4Mux_h
    port map (
            O => \N__28850\,
            I => \N__28841\
        );

    \I__4037\ : InMux
    port map (
            O => \N__28849\,
            I => \N__28834\
        );

    \I__4036\ : InMux
    port map (
            O => \N__28848\,
            I => \N__28834\
        );

    \I__4035\ : InMux
    port map (
            O => \N__28847\,
            I => \N__28834\
        );

    \I__4034\ : Span4Mux_h
    port map (
            O => \N__28844\,
            I => \N__28831\
        );

    \I__4033\ : Span4Mux_h
    port map (
            O => \N__28841\,
            I => \N__28826\
        );

    \I__4032\ : LocalMux
    port map (
            O => \N__28834\,
            I => \N__28826\
        );

    \I__4031\ : Odrv4
    port map (
            O => \N__28831\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0\
        );

    \I__4030\ : Odrv4
    port map (
            O => \N__28826\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0\
        );

    \I__4029\ : InMux
    port map (
            O => \N__28821\,
            I => \N__28812\
        );

    \I__4028\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28812\
        );

    \I__4027\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28812\
        );

    \I__4026\ : LocalMux
    port map (
            O => \N__28812\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_19\
        );

    \I__4025\ : InMux
    port map (
            O => \N__28809\,
            I => \N__28806\
        );

    \I__4024\ : LocalMux
    port map (
            O => \N__28806\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_13\
        );

    \I__4023\ : CascadeMux
    port map (
            O => \N__28803\,
            I => \N__28800\
        );

    \I__4022\ : InMux
    port map (
            O => \N__28800\,
            I => \N__28797\
        );

    \I__4021\ : LocalMux
    port map (
            O => \N__28797\,
            I => \N__28793\
        );

    \I__4020\ : InMux
    port map (
            O => \N__28796\,
            I => \N__28790\
        );

    \I__4019\ : Span12Mux_s9_v
    port map (
            O => \N__28793\,
            I => \N__28787\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__28790\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_8
        );

    \I__4017\ : Odrv12
    port map (
            O => \N__28787\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_8
        );

    \I__4016\ : CascadeMux
    port map (
            O => \N__28782\,
            I => \N__28779\
        );

    \I__4015\ : InMux
    port map (
            O => \N__28779\,
            I => \N__28776\
        );

    \I__4014\ : LocalMux
    port map (
            O => \N__28776\,
            I => \N__28773\
        );

    \I__4013\ : Span4Mux_v
    port map (
            O => \N__28773\,
            I => \N__28770\
        );

    \I__4012\ : Span4Mux_h
    port map (
            O => \N__28770\,
            I => \N__28767\
        );

    \I__4011\ : Odrv4
    port map (
            O => \N__28767\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_0
        );

    \I__4010\ : CascadeMux
    port map (
            O => \N__28764\,
            I => \N__28761\
        );

    \I__4009\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28758\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__28758\,
            I => \N__28755\
        );

    \I__4007\ : Span12Mux_v
    port map (
            O => \N__28755\,
            I => \N__28752\
        );

    \I__4006\ : Odrv12
    port map (
            O => \N__28752\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_11
        );

    \I__4005\ : InMux
    port map (
            O => \N__28749\,
            I => \N__28746\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__28746\,
            I => \N__28743\
        );

    \I__4003\ : Span4Mux_h
    port map (
            O => \N__28743\,
            I => \N__28740\
        );

    \I__4002\ : Span4Mux_h
    port map (
            O => \N__28740\,
            I => \N__28737\
        );

    \I__4001\ : Span4Mux_v
    port map (
            O => \N__28737\,
            I => \N__28734\
        );

    \I__4000\ : Odrv4
    port map (
            O => \N__28734\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_12
        );

    \I__3999\ : CascadeMux
    port map (
            O => \N__28731\,
            I => \N__28728\
        );

    \I__3998\ : InMux
    port map (
            O => \N__28728\,
            I => \N__28725\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__28725\,
            I => \N__28722\
        );

    \I__3996\ : Span4Mux_v
    port map (
            O => \N__28722\,
            I => \N__28719\
        );

    \I__3995\ : Span4Mux_v
    port map (
            O => \N__28719\,
            I => \N__28716\
        );

    \I__3994\ : Odrv4
    port map (
            O => \N__28716\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_13
        );

    \I__3993\ : InMux
    port map (
            O => \N__28713\,
            I => \N__28710\
        );

    \I__3992\ : LocalMux
    port map (
            O => \N__28710\,
            I => \N__28707\
        );

    \I__3991\ : Span4Mux_v
    port map (
            O => \N__28707\,
            I => \N__28704\
        );

    \I__3990\ : Span4Mux_v
    port map (
            O => \N__28704\,
            I => \N__28701\
        );

    \I__3989\ : Odrv4
    port map (
            O => \N__28701\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_14
        );

    \I__3988\ : InMux
    port map (
            O => \N__28698\,
            I => \N__28695\
        );

    \I__3987\ : LocalMux
    port map (
            O => \N__28695\,
            I => \N__28692\
        );

    \I__3986\ : Span4Mux_v
    port map (
            O => \N__28692\,
            I => \N__28689\
        );

    \I__3985\ : Odrv4
    port map (
            O => \N__28689\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_786\
        );

    \I__3984\ : CascadeMux
    port map (
            O => \N__28686\,
            I => \N__28683\
        );

    \I__3983\ : InMux
    port map (
            O => \N__28683\,
            I => \N__28680\
        );

    \I__3982\ : LocalMux
    port map (
            O => \N__28680\,
            I => \N__28677\
        );

    \I__3981\ : Span4Mux_v
    port map (
            O => \N__28677\,
            I => \N__28674\
        );

    \I__3980\ : Span4Mux_h
    port map (
            O => \N__28674\,
            I => \N__28671\
        );

    \I__3979\ : Span4Mux_v
    port map (
            O => \N__28671\,
            I => \N__28668\
        );

    \I__3978\ : Odrv4
    port map (
            O => \N__28668\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_15
        );

    \I__3977\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28662\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__28662\,
            I => \N__28659\
        );

    \I__3975\ : Odrv12
    port map (
            O => \N__28659\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_20
        );

    \I__3974\ : CascadeMux
    port map (
            O => \N__28656\,
            I => \N__28653\
        );

    \I__3973\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28650\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__28650\,
            I => \N__28647\
        );

    \I__3971\ : Span4Mux_v
    port map (
            O => \N__28647\,
            I => \N__28644\
        );

    \I__3970\ : Span4Mux_h
    port map (
            O => \N__28644\,
            I => \N__28641\
        );

    \I__3969\ : Span4Mux_v
    port map (
            O => \N__28641\,
            I => \N__28638\
        );

    \I__3968\ : Odrv4
    port map (
            O => \N__28638\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_9
        );

    \I__3967\ : InMux
    port map (
            O => \N__28635\,
            I => \N__28632\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__28632\,
            I => \N__28629\
        );

    \I__3965\ : Span12Mux_h
    port map (
            O => \N__28629\,
            I => \N__28626\
        );

    \I__3964\ : Span12Mux_v
    port map (
            O => \N__28626\,
            I => \N__28623\
        );

    \I__3963\ : Odrv12
    port map (
            O => \N__28623\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_4
        );

    \I__3962\ : CascadeMux
    port map (
            O => \N__28620\,
            I => \N__28617\
        );

    \I__3961\ : InMux
    port map (
            O => \N__28617\,
            I => \N__28614\
        );

    \I__3960\ : LocalMux
    port map (
            O => \N__28614\,
            I => \N__28611\
        );

    \I__3959\ : Span4Mux_v
    port map (
            O => \N__28611\,
            I => \N__28608\
        );

    \I__3958\ : Span4Mux_v
    port map (
            O => \N__28608\,
            I => \N__28605\
        );

    \I__3957\ : Odrv4
    port map (
            O => \N__28605\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_4
        );

    \I__3956\ : InMux
    port map (
            O => \N__28602\,
            I => \N__28599\
        );

    \I__3955\ : LocalMux
    port map (
            O => \N__28599\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_4\
        );

    \I__3954\ : InMux
    port map (
            O => \N__28596\,
            I => \N__28593\
        );

    \I__3953\ : LocalMux
    port map (
            O => \N__28593\,
            I => \N__28590\
        );

    \I__3952\ : Span4Mux_h
    port map (
            O => \N__28590\,
            I => \N__28587\
        );

    \I__3951\ : Odrv4
    port map (
            O => \N__28587\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_9
        );

    \I__3950\ : InMux
    port map (
            O => \N__28584\,
            I => \N__28580\
        );

    \I__3949\ : InMux
    port map (
            O => \N__28583\,
            I => \N__28577\
        );

    \I__3948\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28574\
        );

    \I__3947\ : LocalMux
    port map (
            O => \N__28577\,
            I => \N__28569\
        );

    \I__3946\ : Span4Mux_v
    port map (
            O => \N__28574\,
            I => \N__28569\
        );

    \I__3945\ : Odrv4
    port map (
            O => \N__28569\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_30
        );

    \I__3944\ : CascadeMux
    port map (
            O => \N__28566\,
            I => \N__28563\
        );

    \I__3943\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28559\
        );

    \I__3942\ : CascadeMux
    port map (
            O => \N__28562\,
            I => \N__28556\
        );

    \I__3941\ : LocalMux
    port map (
            O => \N__28559\,
            I => \N__28553\
        );

    \I__3940\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28550\
        );

    \I__3939\ : Span4Mux_v
    port map (
            O => \N__28553\,
            I => \N__28547\
        );

    \I__3938\ : LocalMux
    port map (
            O => \N__28550\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_4
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__28547\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_4
        );

    \I__3936\ : InMux
    port map (
            O => \N__28542\,
            I => \N__28539\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__28539\,
            I => \N__28536\
        );

    \I__3934\ : Span4Mux_h
    port map (
            O => \N__28536\,
            I => \N__28533\
        );

    \I__3933\ : Span4Mux_v
    port map (
            O => \N__28533\,
            I => \N__28530\
        );

    \I__3932\ : Odrv4
    port map (
            O => \N__28530\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_9
        );

    \I__3931\ : InMux
    port map (
            O => \N__28527\,
            I => \N__28524\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28521\
        );

    \I__3929\ : Span4Mux_v
    port map (
            O => \N__28521\,
            I => \N__28518\
        );

    \I__3928\ : Span4Mux_h
    port map (
            O => \N__28518\,
            I => \N__28515\
        );

    \I__3927\ : Odrv4
    port map (
            O => \N__28515\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_29
        );

    \I__3926\ : InMux
    port map (
            O => \N__28512\,
            I => \N__28509\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__28509\,
            I => \N__28506\
        );

    \I__3924\ : Span4Mux_h
    port map (
            O => \N__28506\,
            I => \N__28503\
        );

    \I__3923\ : Odrv4
    port map (
            O => \N__28503\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_3
        );

    \I__3922\ : CascadeMux
    port map (
            O => \N__28500\,
            I => \N__28497\
        );

    \I__3921\ : InMux
    port map (
            O => \N__28497\,
            I => \N__28494\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__28494\,
            I => \N__28491\
        );

    \I__3919\ : Odrv4
    port map (
            O => \N__28491\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_907\
        );

    \I__3918\ : CascadeMux
    port map (
            O => \N__28488\,
            I => \N__28485\
        );

    \I__3917\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28482\
        );

    \I__3916\ : LocalMux
    port map (
            O => \N__28482\,
            I => \N__28479\
        );

    \I__3915\ : Span4Mux_h
    port map (
            O => \N__28479\,
            I => \N__28476\
        );

    \I__3914\ : Span4Mux_h
    port map (
            O => \N__28476\,
            I => \N__28473\
        );

    \I__3913\ : Odrv4
    port map (
            O => \N__28473\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_30
        );

    \I__3912\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28467\
        );

    \I__3911\ : LocalMux
    port map (
            O => \N__28467\,
            I => \N__28464\
        );

    \I__3910\ : Odrv4
    port map (
            O => \N__28464\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_621\
        );

    \I__3909\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28458\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__28458\,
            I => \N__28455\
        );

    \I__3907\ : Span4Mux_h
    port map (
            O => \N__28455\,
            I => \N__28452\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__28452\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_31
        );

    \I__3905\ : InMux
    port map (
            O => \N__28449\,
            I => \N__28446\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28443\
        );

    \I__3903\ : Span4Mux_h
    port map (
            O => \N__28443\,
            I => \N__28440\
        );

    \I__3902\ : Odrv4
    port map (
            O => \N__28440\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_610\
        );

    \I__3901\ : CascadeMux
    port map (
            O => \N__28437\,
            I => \N__28434\
        );

    \I__3900\ : InMux
    port map (
            O => \N__28434\,
            I => \N__28431\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__28431\,
            I => \N__28428\
        );

    \I__3898\ : Span4Mux_h
    port map (
            O => \N__28428\,
            I => \N__28425\
        );

    \I__3897\ : Odrv4
    port map (
            O => \N__28425\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_1
        );

    \I__3896\ : InMux
    port map (
            O => \N__28422\,
            I => \N__28419\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__28419\,
            I => \N__28416\
        );

    \I__3894\ : Span4Mux_v
    port map (
            O => \N__28416\,
            I => \N__28413\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__28413\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316\
        );

    \I__3892\ : InMux
    port map (
            O => \N__28410\,
            I => \N__28407\
        );

    \I__3891\ : LocalMux
    port map (
            O => \N__28407\,
            I => \N__28404\
        );

    \I__3890\ : Span4Mux_v
    port map (
            O => \N__28404\,
            I => \N__28401\
        );

    \I__3889\ : Span4Mux_h
    port map (
            O => \N__28401\,
            I => \N__28398\
        );

    \I__3888\ : Sp12to4
    port map (
            O => \N__28398\,
            I => \N__28395\
        );

    \I__3887\ : Odrv12
    port map (
            O => \N__28395\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_5
        );

    \I__3886\ : CascadeMux
    port map (
            O => \N__28392\,
            I => \N__28389\
        );

    \I__3885\ : InMux
    port map (
            O => \N__28389\,
            I => \N__28386\
        );

    \I__3884\ : LocalMux
    port map (
            O => \N__28386\,
            I => \N__28383\
        );

    \I__3883\ : Span4Mux_h
    port map (
            O => \N__28383\,
            I => \N__28380\
        );

    \I__3882\ : Odrv4
    port map (
            O => \N__28380\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_885\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__28377\,
            I => \N__28374\
        );

    \I__3880\ : InMux
    port map (
            O => \N__28374\,
            I => \N__28371\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__28371\,
            I => \N__28368\
        );

    \I__3878\ : Span4Mux_v
    port map (
            O => \N__28368\,
            I => \N__28365\
        );

    \I__3877\ : Span4Mux_h
    port map (
            O => \N__28365\,
            I => \N__28362\
        );

    \I__3876\ : Odrv4
    port map (
            O => \N__28362\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_6
        );

    \I__3875\ : CascadeMux
    port map (
            O => \N__28359\,
            I => \N__28356\
        );

    \I__3874\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28353\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__28353\,
            I => \N__28350\
        );

    \I__3872\ : Odrv4
    port map (
            O => \N__28350\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_874\
        );

    \I__3871\ : InMux
    port map (
            O => \N__28347\,
            I => \N__28344\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__28344\,
            I => \N__28341\
        );

    \I__3869\ : Span4Mux_v
    port map (
            O => \N__28341\,
            I => \N__28338\
        );

    \I__3868\ : Span4Mux_h
    port map (
            O => \N__28338\,
            I => \N__28335\
        );

    \I__3867\ : Span4Mux_v
    port map (
            O => \N__28335\,
            I => \N__28332\
        );

    \I__3866\ : Span4Mux_v
    port map (
            O => \N__28332\,
            I => \N__28329\
        );

    \I__3865\ : Odrv4
    port map (
            O => \N__28329\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_9
        );

    \I__3864\ : CascadeMux
    port map (
            O => \N__28326\,
            I => \N__28322\
        );

    \I__3863\ : InMux
    port map (
            O => \N__28325\,
            I => \N__28314\
        );

    \I__3862\ : InMux
    port map (
            O => \N__28322\,
            I => \N__28314\
        );

    \I__3861\ : InMux
    port map (
            O => \N__28321\,
            I => \N__28314\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__28314\,
            I => cemf_module_64ch_ctrl_inst1_data_clkstopmask_4
        );

    \I__3859\ : InMux
    port map (
            O => \N__28311\,
            I => \N__28308\
        );

    \I__3858\ : LocalMux
    port map (
            O => \N__28308\,
            I => \N__28305\
        );

    \I__3857\ : Span4Mux_v
    port map (
            O => \N__28305\,
            I => \N__28302\
        );

    \I__3856\ : Odrv4
    port map (
            O => \N__28302\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_26
        );

    \I__3855\ : InMux
    port map (
            O => \N__28299\,
            I => \N__28296\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__28296\,
            I => \N__28293\
        );

    \I__3853\ : Span4Mux_v
    port map (
            O => \N__28293\,
            I => \N__28290\
        );

    \I__3852\ : Span4Mux_h
    port map (
            O => \N__28290\,
            I => \N__28287\
        );

    \I__3851\ : Span4Mux_v
    port map (
            O => \N__28287\,
            I => \N__28284\
        );

    \I__3850\ : Odrv4
    port map (
            O => \N__28284\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_26
        );

    \I__3849\ : CascadeMux
    port map (
            O => \N__28281\,
            I => \N__28278\
        );

    \I__3848\ : InMux
    port map (
            O => \N__28278\,
            I => \N__28275\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__28275\,
            I => \N__28272\
        );

    \I__3846\ : Span4Mux_v
    port map (
            O => \N__28272\,
            I => \N__28269\
        );

    \I__3845\ : Span4Mux_h
    port map (
            O => \N__28269\,
            I => \N__28266\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__28266\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_26
        );

    \I__3843\ : InMux
    port map (
            O => \N__28263\,
            I => \N__28260\
        );

    \I__3842\ : LocalMux
    port map (
            O => \N__28260\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_0_26\
        );

    \I__3841\ : CascadeMux
    port map (
            O => \N__28257\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_1_26_cascade_\
        );

    \I__3840\ : InMux
    port map (
            O => \N__28254\,
            I => \N__28251\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__28251\,
            I => \N__28248\
        );

    \I__3838\ : Span12Mux_h
    port map (
            O => \N__28248\,
            I => \N__28245\
        );

    \I__3837\ : Odrv12
    port map (
            O => \N__28245\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_26
        );

    \I__3836\ : InMux
    port map (
            O => \N__28242\,
            I => \N__28239\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__28239\,
            I => \N__28236\
        );

    \I__3834\ : Span4Mux_h
    port map (
            O => \N__28236\,
            I => \N__28233\
        );

    \I__3833\ : Span4Mux_h
    port map (
            O => \N__28233\,
            I => \N__28230\
        );

    \I__3832\ : Odrv4
    port map (
            O => \N__28230\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_21
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__28227\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_30_cascade_\
        );

    \I__3830\ : InMux
    port map (
            O => \N__28224\,
            I => \N__28221\
        );

    \I__3829\ : LocalMux
    port map (
            O => \N__28221\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_30\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__28218\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_30_cascade_\
        );

    \I__3827\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28212\
        );

    \I__3826\ : LocalMux
    port map (
            O => \N__28212\,
            I => \N__28209\
        );

    \I__3825\ : Odrv4
    port map (
            O => \N__28209\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_30\
        );

    \I__3824\ : InMux
    port map (
            O => \N__28206\,
            I => \N__28203\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__28203\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_30\
        );

    \I__3822\ : InMux
    port map (
            O => \N__28200\,
            I => \N__28197\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__28197\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_30\
        );

    \I__3820\ : CascadeMux
    port map (
            O => \N__28194\,
            I => \N__28191\
        );

    \I__3819\ : InMux
    port map (
            O => \N__28191\,
            I => \N__28188\
        );

    \I__3818\ : LocalMux
    port map (
            O => \N__28188\,
            I => \N__28185\
        );

    \I__3817\ : Odrv4
    port map (
            O => \N__28185\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_30\
        );

    \I__3816\ : InMux
    port map (
            O => \N__28182\,
            I => \N__28178\
        );

    \I__3815\ : InMux
    port map (
            O => \N__28181\,
            I => \N__28175\
        );

    \I__3814\ : LocalMux
    port map (
            O => \N__28178\,
            I => \N__28171\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__28175\,
            I => \N__28168\
        );

    \I__3812\ : InMux
    port map (
            O => \N__28174\,
            I => \N__28165\
        );

    \I__3811\ : Span4Mux_v
    port map (
            O => \N__28171\,
            I => \N__28162\
        );

    \I__3810\ : Span12Mux_v
    port map (
            O => \N__28168\,
            I => \N__28159\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__28165\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_31
        );

    \I__3808\ : Odrv4
    port map (
            O => \N__28162\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_31
        );

    \I__3807\ : Odrv12
    port map (
            O => \N__28159\,
            I => cemf_module_64ch_ctrl_inst1_s_data_system_o_31
        );

    \I__3806\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28149\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__28149\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_31\
        );

    \I__3804\ : CascadeMux
    port map (
            O => \N__28146\,
            I => \N__28143\
        );

    \I__3803\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28140\
        );

    \I__3802\ : LocalMux
    port map (
            O => \N__28140\,
            I => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_31\
        );

    \I__3801\ : InMux
    port map (
            O => \N__28137\,
            I => \N__28134\
        );

    \I__3800\ : LocalMux
    port map (
            O => \N__28134\,
            I => \N__28131\
        );

    \I__3799\ : Span4Mux_v
    port map (
            O => \N__28131\,
            I => \N__28128\
        );

    \I__3798\ : Odrv4
    port map (
            O => \N__28128\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_4\
        );

    \I__3797\ : InMux
    port map (
            O => \N__28125\,
            I => \N__28122\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__28122\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_8\
        );

    \I__3795\ : InMux
    port map (
            O => \N__28119\,
            I => \N__28116\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__28116\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_8\
        );

    \I__3793\ : CascadeMux
    port map (
            O => \N__28113\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_8_cascade_\
        );

    \I__3792\ : InMux
    port map (
            O => \N__28110\,
            I => \N__28107\
        );

    \I__3791\ : LocalMux
    port map (
            O => \N__28107\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_8\
        );

    \I__3790\ : InMux
    port map (
            O => \N__28104\,
            I => \N__28101\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__28101\,
            I => \N__28098\
        );

    \I__3788\ : Span4Mux_v
    port map (
            O => \N__28098\,
            I => \N__28095\
        );

    \I__3787\ : Span4Mux_v
    port map (
            O => \N__28095\,
            I => \N__28092\
        );

    \I__3786\ : Odrv4
    port map (
            O => \N__28092\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_14
        );

    \I__3785\ : CascadeMux
    port map (
            O => \N__28089\,
            I => \N__28086\
        );

    \I__3784\ : InMux
    port map (
            O => \N__28086\,
            I => \N__28083\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__28083\,
            I => \N__28080\
        );

    \I__3782\ : Span4Mux_v
    port map (
            O => \N__28080\,
            I => \N__28077\
        );

    \I__3781\ : Span4Mux_h
    port map (
            O => \N__28077\,
            I => \N__28074\
        );

    \I__3780\ : Odrv4
    port map (
            O => \N__28074\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_14
        );

    \I__3779\ : CascadeMux
    port map (
            O => \N__28071\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_14_cascade_\
        );

    \I__3778\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28065\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__28065\,
            I => \N__28062\
        );

    \I__3776\ : Span4Mux_h
    port map (
            O => \N__28062\,
            I => \N__28059\
        );

    \I__3775\ : Span4Mux_v
    port map (
            O => \N__28059\,
            I => \N__28056\
        );

    \I__3774\ : Odrv4
    port map (
            O => \N__28056\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_14
        );

    \I__3773\ : CascadeMux
    port map (
            O => \N__28053\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_14_cascade_\
        );

    \I__3772\ : CascadeMux
    port map (
            O => \N__28050\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_14_cascade_\
        );

    \I__3771\ : InMux
    port map (
            O => \N__28047\,
            I => \N__28044\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__28044\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_14\
        );

    \I__3769\ : InMux
    port map (
            O => \N__28041\,
            I => \N__28038\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__28038\,
            I => \N__28035\
        );

    \I__3767\ : Span4Mux_h
    port map (
            O => \N__28035\,
            I => \N__28032\
        );

    \I__3766\ : Span4Mux_v
    port map (
            O => \N__28032\,
            I => \N__28029\
        );

    \I__3765\ : Odrv4
    port map (
            O => \N__28029\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_22
        );

    \I__3764\ : InMux
    port map (
            O => \N__28026\,
            I => \N__28023\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__28023\,
            I => \N__28020\
        );

    \I__3762\ : Span4Mux_v
    port map (
            O => \N__28020\,
            I => \N__28017\
        );

    \I__3761\ : Span4Mux_v
    port map (
            O => \N__28017\,
            I => \N__28014\
        );

    \I__3760\ : Odrv4
    port map (
            O => \N__28014\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_30
        );

    \I__3759\ : CascadeMux
    port map (
            O => \N__28011\,
            I => \N__28008\
        );

    \I__3758\ : InMux
    port map (
            O => \N__28008\,
            I => \N__28005\
        );

    \I__3757\ : LocalMux
    port map (
            O => \N__28005\,
            I => \N__28002\
        );

    \I__3756\ : Span4Mux_v
    port map (
            O => \N__28002\,
            I => \N__27999\
        );

    \I__3755\ : Odrv4
    port map (
            O => \N__27999\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_30
        );

    \I__3754\ : InMux
    port map (
            O => \N__27996\,
            I => \N__27993\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__27993\,
            I => \N__27990\
        );

    \I__3752\ : Span4Mux_v
    port map (
            O => \N__27990\,
            I => \N__27987\
        );

    \I__3751\ : Span4Mux_v
    port map (
            O => \N__27987\,
            I => \N__27984\
        );

    \I__3750\ : IoSpan4Mux
    port map (
            O => \N__27984\,
            I => \N__27981\
        );

    \I__3749\ : Odrv4
    port map (
            O => \N__27981\,
            I => sync_50hz_c
        );

    \I__3748\ : InMux
    port map (
            O => \N__27978\,
            I => \N__27974\
        );

    \I__3747\ : InMux
    port map (
            O => \N__27977\,
            I => \N__27971\
        );

    \I__3746\ : LocalMux
    port map (
            O => \N__27974\,
            I => \cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0\
        );

    \I__3745\ : LocalMux
    port map (
            O => \N__27971\,
            I => \cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0\
        );

    \I__3744\ : InMux
    port map (
            O => \N__27966\,
            I => \N__27962\
        );

    \I__3743\ : InMux
    port map (
            O => \N__27965\,
            I => \N__27959\
        );

    \I__3742\ : LocalMux
    port map (
            O => \N__27962\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config\
        );

    \I__3741\ : LocalMux
    port map (
            O => \N__27959\,
            I => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__27954\,
            I => \cemf_module_64ch_ctrl_inst1.N_410_0_cascade_\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__27951\,
            I => \cemf_module_64ch_ctrl_inst1.N_68_0_cascade_\
        );

    \I__3738\ : InMux
    port map (
            O => \N__27948\,
            I => \N__27945\
        );

    \I__3737\ : LocalMux
    port map (
            O => \N__27945\,
            I => \N__27942\
        );

    \I__3736\ : Span4Mux_v
    port map (
            O => \N__27942\,
            I => \N__27939\
        );

    \I__3735\ : Span4Mux_h
    port map (
            O => \N__27939\,
            I => \N__27936\
        );

    \I__3734\ : Odrv4
    port map (
            O => \N__27936\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_8
        );

    \I__3733\ : CascadeMux
    port map (
            O => \N__27933\,
            I => \N__27930\
        );

    \I__3732\ : InMux
    port map (
            O => \N__27930\,
            I => \N__27927\
        );

    \I__3731\ : LocalMux
    port map (
            O => \N__27927\,
            I => \N__27924\
        );

    \I__3730\ : Span4Mux_v
    port map (
            O => \N__27924\,
            I => \N__27921\
        );

    \I__3729\ : Span4Mux_h
    port map (
            O => \N__27921\,
            I => \N__27918\
        );

    \I__3728\ : Odrv4
    port map (
            O => \N__27918\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_8
        );

    \I__3727\ : CascadeMux
    port map (
            O => \N__27915\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_8_cascade_\
        );

    \I__3726\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27908\
        );

    \I__3725\ : InMux
    port map (
            O => \N__27911\,
            I => \N__27905\
        );

    \I__3724\ : LocalMux
    port map (
            O => \N__27908\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2\
        );

    \I__3723\ : LocalMux
    port map (
            O => \N__27905\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2\
        );

    \I__3722\ : InMux
    port map (
            O => \N__27900\,
            I => \N__27897\
        );

    \I__3721\ : LocalMux
    port map (
            O => \N__27897\,
            I => \N__27894\
        );

    \I__3720\ : Span4Mux_h
    port map (
            O => \N__27894\,
            I => \N__27891\
        );

    \I__3719\ : Odrv4
    port map (
            O => \N__27891\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_1\
        );

    \I__3718\ : CascadeMux
    port map (
            O => \N__27888\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287_cascade_\
        );

    \I__3717\ : InMux
    port map (
            O => \N__27885\,
            I => \N__27881\
        );

    \I__3716\ : InMux
    port map (
            O => \N__27884\,
            I => \N__27878\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__27881\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0\
        );

    \I__3714\ : LocalMux
    port map (
            O => \N__27878\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0\
        );

    \I__3713\ : InMux
    port map (
            O => \N__27873\,
            I => \bfn_11_19_0_\
        );

    \I__3712\ : InMux
    port map (
            O => \N__27870\,
            I => \N__27866\
        );

    \I__3711\ : InMux
    port map (
            O => \N__27869\,
            I => \N__27863\
        );

    \I__3710\ : LocalMux
    port map (
            O => \N__27866\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1\
        );

    \I__3709\ : LocalMux
    port map (
            O => \N__27863\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1\
        );

    \I__3708\ : InMux
    port map (
            O => \N__27858\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0\
        );

    \I__3707\ : CascadeMux
    port map (
            O => \N__27855\,
            I => \N__27851\
        );

    \I__3706\ : InMux
    port map (
            O => \N__27854\,
            I => \N__27848\
        );

    \I__3705\ : InMux
    port map (
            O => \N__27851\,
            I => \N__27845\
        );

    \I__3704\ : LocalMux
    port map (
            O => \N__27848\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__27845\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2\
        );

    \I__3702\ : InMux
    port map (
            O => \N__27840\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1\
        );

    \I__3701\ : InMux
    port map (
            O => \N__27837\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2\
        );

    \I__3700\ : InMux
    port map (
            O => \N__27834\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_3\
        );

    \I__3699\ : InMux
    port map (
            O => \N__27831\,
            I => \N__27828\
        );

    \I__3698\ : LocalMux
    port map (
            O => \N__27828\,
            I => \N__27824\
        );

    \I__3697\ : CascadeMux
    port map (
            O => \N__27827\,
            I => \N__27818\
        );

    \I__3696\ : Span4Mux_v
    port map (
            O => \N__27824\,
            I => \N__27814\
        );

    \I__3695\ : InMux
    port map (
            O => \N__27823\,
            I => \N__27803\
        );

    \I__3694\ : InMux
    port map (
            O => \N__27822\,
            I => \N__27803\
        );

    \I__3693\ : InMux
    port map (
            O => \N__27821\,
            I => \N__27803\
        );

    \I__3692\ : InMux
    port map (
            O => \N__27818\,
            I => \N__27803\
        );

    \I__3691\ : InMux
    port map (
            O => \N__27817\,
            I => \N__27803\
        );

    \I__3690\ : Odrv4
    port map (
            O => \N__27814\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0\
        );

    \I__3689\ : LocalMux
    port map (
            O => \N__27803\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0\
        );

    \I__3688\ : CascadeMux
    port map (
            O => \N__27798\,
            I => \N__27795\
        );

    \I__3687\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27792\
        );

    \I__3686\ : LocalMux
    port map (
            O => \N__27792\,
            I => \N__27789\
        );

    \I__3685\ : Span4Mux_v
    port map (
            O => \N__27789\,
            I => \N__27765\
        );

    \I__3684\ : InMux
    port map (
            O => \N__27788\,
            I => \N__27762\
        );

    \I__3683\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27745\
        );

    \I__3682\ : InMux
    port map (
            O => \N__27786\,
            I => \N__27745\
        );

    \I__3681\ : InMux
    port map (
            O => \N__27785\,
            I => \N__27745\
        );

    \I__3680\ : InMux
    port map (
            O => \N__27784\,
            I => \N__27745\
        );

    \I__3679\ : InMux
    port map (
            O => \N__27783\,
            I => \N__27745\
        );

    \I__3678\ : InMux
    port map (
            O => \N__27782\,
            I => \N__27745\
        );

    \I__3677\ : InMux
    port map (
            O => \N__27781\,
            I => \N__27745\
        );

    \I__3676\ : InMux
    port map (
            O => \N__27780\,
            I => \N__27745\
        );

    \I__3675\ : InMux
    port map (
            O => \N__27779\,
            I => \N__27728\
        );

    \I__3674\ : InMux
    port map (
            O => \N__27778\,
            I => \N__27728\
        );

    \I__3673\ : InMux
    port map (
            O => \N__27777\,
            I => \N__27728\
        );

    \I__3672\ : InMux
    port map (
            O => \N__27776\,
            I => \N__27728\
        );

    \I__3671\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27728\
        );

    \I__3670\ : InMux
    port map (
            O => \N__27774\,
            I => \N__27728\
        );

    \I__3669\ : InMux
    port map (
            O => \N__27773\,
            I => \N__27728\
        );

    \I__3668\ : InMux
    port map (
            O => \N__27772\,
            I => \N__27728\
        );

    \I__3667\ : InMux
    port map (
            O => \N__27771\,
            I => \N__27719\
        );

    \I__3666\ : InMux
    port map (
            O => \N__27770\,
            I => \N__27719\
        );

    \I__3665\ : InMux
    port map (
            O => \N__27769\,
            I => \N__27719\
        );

    \I__3664\ : InMux
    port map (
            O => \N__27768\,
            I => \N__27719\
        );

    \I__3663\ : Odrv4
    port map (
            O => \N__27765\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\
        );

    \I__3662\ : LocalMux
    port map (
            O => \N__27762\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__27745\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__27728\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__27719\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\
        );

    \I__3658\ : CEMux
    port map (
            O => \N__27708\,
            I => \N__27704\
        );

    \I__3657\ : CEMux
    port map (
            O => \N__27707\,
            I => \N__27701\
        );

    \I__3656\ : LocalMux
    port map (
            O => \N__27704\,
            I => \N__27698\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__27701\,
            I => \N__27695\
        );

    \I__3654\ : Odrv4
    port map (
            O => \N__27698\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i\
        );

    \I__3653\ : Odrv4
    port map (
            O => \N__27695\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i\
        );

    \I__3652\ : CascadeMux
    port map (
            O => \N__27690\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996_cascade_\
        );

    \I__3651\ : InMux
    port map (
            O => \N__27687\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1\
        );

    \I__3650\ : InMux
    port map (
            O => \N__27684\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2\
        );

    \I__3649\ : InMux
    port map (
            O => \N__27681\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_3\
        );

    \I__3648\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27675\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__27675\,
            I => \N__27672\
        );

    \I__3646\ : Span4Mux_h
    port map (
            O => \N__27672\,
            I => \N__27669\
        );

    \I__3645\ : Odrv4
    port map (
            O => \N__27669\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2\
        );

    \I__3644\ : InMux
    port map (
            O => \N__27666\,
            I => \N__27662\
        );

    \I__3643\ : InMux
    port map (
            O => \N__27665\,
            I => \N__27659\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__27662\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__27659\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4\
        );

    \I__3640\ : InMux
    port map (
            O => \N__27654\,
            I => \N__27650\
        );

    \I__3639\ : InMux
    port map (
            O => \N__27653\,
            I => \N__27647\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__27650\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__27647\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2\
        );

    \I__3636\ : CascadeMux
    port map (
            O => \N__27642\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2_cascade_\
        );

    \I__3635\ : InMux
    port map (
            O => \N__27639\,
            I => \N__27635\
        );

    \I__3634\ : InMux
    port map (
            O => \N__27638\,
            I => \N__27632\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__27635\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1\
        );

    \I__3632\ : LocalMux
    port map (
            O => \N__27632\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1\
        );

    \I__3631\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27623\
        );

    \I__3630\ : InMux
    port map (
            O => \N__27626\,
            I => \N__27620\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__27623\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__27620\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3\
        );

    \I__3627\ : CascadeMux
    port map (
            O => \N__27615\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m7_3_cascade_\
        );

    \I__3626\ : InMux
    port map (
            O => \N__27612\,
            I => \N__27608\
        );

    \I__3625\ : InMux
    port map (
            O => \N__27611\,
            I => \N__27605\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__27608\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__27605\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0\
        );

    \I__3622\ : InMux
    port map (
            O => \N__27600\,
            I => \N__27591\
        );

    \I__3621\ : InMux
    port map (
            O => \N__27599\,
            I => \N__27591\
        );

    \I__3620\ : InMux
    port map (
            O => \N__27598\,
            I => \N__27584\
        );

    \I__3619\ : InMux
    port map (
            O => \N__27597\,
            I => \N__27584\
        );

    \I__3618\ : InMux
    port map (
            O => \N__27596\,
            I => \N__27584\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__27591\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2\
        );

    \I__3616\ : LocalMux
    port map (
            O => \N__27584\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2\
        );

    \I__3615\ : InMux
    port map (
            O => \N__27579\,
            I => \N__27573\
        );

    \I__3614\ : InMux
    port map (
            O => \N__27578\,
            I => \N__27573\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__27573\,
            I => \N__27569\
        );

    \I__3612\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27564\
        );

    \I__3611\ : Span4Mux_v
    port map (
            O => \N__27569\,
            I => \N__27561\
        );

    \I__3610\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27556\
        );

    \I__3609\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27556\
        );

    \I__3608\ : LocalMux
    port map (
            O => \N__27564\,
            I => \N__27553\
        );

    \I__3607\ : Sp12to4
    port map (
            O => \N__27561\,
            I => \N__27548\
        );

    \I__3606\ : LocalMux
    port map (
            O => \N__27556\,
            I => \N__27548\
        );

    \I__3605\ : Span4Mux_v
    port map (
            O => \N__27553\,
            I => \N__27545\
        );

    \I__3604\ : Odrv12
    port map (
            O => \N__27548\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__27545\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46\
        );

    \I__3602\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27537\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__27537\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_3\
        );

    \I__3600\ : CascadeMux
    port map (
            O => \N__27534\,
            I => \N__27531\
        );

    \I__3599\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27528\
        );

    \I__3598\ : LocalMux
    port map (
            O => \N__27528\,
            I => \N__27525\
        );

    \I__3597\ : Span4Mux_h
    port map (
            O => \N__27525\,
            I => \N__27522\
        );

    \I__3596\ : Odrv4
    port map (
            O => \N__27522\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_3
        );

    \I__3595\ : InMux
    port map (
            O => \N__27519\,
            I => \N__27516\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__27516\,
            I => \N__27513\
        );

    \I__3593\ : Odrv4
    port map (
            O => \N__27513\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3\
        );

    \I__3592\ : InMux
    port map (
            O => \N__27510\,
            I => \N__27507\
        );

    \I__3591\ : LocalMux
    port map (
            O => \N__27507\,
            I => \N__27504\
        );

    \I__3590\ : Span4Mux_h
    port map (
            O => \N__27504\,
            I => \N__27501\
        );

    \I__3589\ : Odrv4
    port map (
            O => \N__27501\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_4
        );

    \I__3588\ : CascadeMux
    port map (
            O => \N__27498\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_cascade_\
        );

    \I__3587\ : InMux
    port map (
            O => \N__27495\,
            I => \N__27492\
        );

    \I__3586\ : LocalMux
    port map (
            O => \N__27492\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_5\
        );

    \I__3585\ : InMux
    port map (
            O => \N__27489\,
            I => \N__27486\
        );

    \I__3584\ : LocalMux
    port map (
            O => \N__27486\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_4\
        );

    \I__3583\ : CascadeMux
    port map (
            O => \N__27483\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_4_cascade_\
        );

    \I__3582\ : InMux
    port map (
            O => \N__27480\,
            I => \N__27477\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__27477\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_4\
        );

    \I__3580\ : InMux
    port map (
            O => \N__27474\,
            I => \bfn_11_15_0_\
        );

    \I__3579\ : InMux
    port map (
            O => \N__27471\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0\
        );

    \I__3578\ : CascadeMux
    port map (
            O => \N__27468\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_31_cascade_\
        );

    \I__3577\ : InMux
    port map (
            O => \N__27465\,
            I => \N__27462\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__27462\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_31\
        );

    \I__3575\ : CascadeMux
    port map (
            O => \N__27459\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_31_cascade_\
        );

    \I__3574\ : InMux
    port map (
            O => \N__27456\,
            I => \N__27453\
        );

    \I__3573\ : LocalMux
    port map (
            O => \N__27453\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_31\
        );

    \I__3572\ : InMux
    port map (
            O => \N__27450\,
            I => \N__27447\
        );

    \I__3571\ : LocalMux
    port map (
            O => \N__27447\,
            I => \N__27444\
        );

    \I__3570\ : Span4Mux_v
    port map (
            O => \N__27444\,
            I => \N__27441\
        );

    \I__3569\ : Odrv4
    port map (
            O => \N__27441\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_27
        );

    \I__3568\ : InMux
    port map (
            O => \N__27438\,
            I => \N__27435\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__27435\,
            I => \N__27432\
        );

    \I__3566\ : Span4Mux_h
    port map (
            O => \N__27432\,
            I => \N__27429\
        );

    \I__3565\ : Odrv4
    port map (
            O => \N__27429\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_28
        );

    \I__3564\ : InMux
    port map (
            O => \N__27426\,
            I => \N__27423\
        );

    \I__3563\ : LocalMux
    port map (
            O => \N__27423\,
            I => \N__27420\
        );

    \I__3562\ : Span4Mux_h
    port map (
            O => \N__27420\,
            I => \N__27417\
        );

    \I__3561\ : Odrv4
    port map (
            O => \N__27417\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_29
        );

    \I__3560\ : InMux
    port map (
            O => \N__27414\,
            I => \N__27411\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__27411\,
            I => \N__27408\
        );

    \I__3558\ : Span4Mux_v
    port map (
            O => \N__27408\,
            I => \N__27405\
        );

    \I__3557\ : Odrv4
    port map (
            O => \N__27405\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_30
        );

    \I__3556\ : InMux
    port map (
            O => \N__27402\,
            I => \N__27399\
        );

    \I__3555\ : LocalMux
    port map (
            O => \N__27399\,
            I => \N__27396\
        );

    \I__3554\ : Span4Mux_h
    port map (
            O => \N__27396\,
            I => \N__27393\
        );

    \I__3553\ : Odrv4
    port map (
            O => \N__27393\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_31
        );

    \I__3552\ : InMux
    port map (
            O => \N__27390\,
            I => \N__27387\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__27387\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_31\
        );

    \I__3550\ : InMux
    port map (
            O => \N__27384\,
            I => \N__27381\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__27381\,
            I => \N__27378\
        );

    \I__3548\ : Span4Mux_v
    port map (
            O => \N__27378\,
            I => \N__27375\
        );

    \I__3547\ : Odrv4
    port map (
            O => \N__27375\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_1\
        );

    \I__3546\ : CascadeMux
    port map (
            O => \N__27372\,
            I => \N__27369\
        );

    \I__3545\ : InMux
    port map (
            O => \N__27369\,
            I => \N__27366\
        );

    \I__3544\ : LocalMux
    port map (
            O => \N__27366\,
            I => \N__27363\
        );

    \I__3543\ : Odrv4
    port map (
            O => \N__27363\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_10
        );

    \I__3542\ : CascadeMux
    port map (
            O => \N__27360\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_3_cascade_\
        );

    \I__3541\ : InMux
    port map (
            O => \N__27357\,
            I => \N__27354\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__27354\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_3\
        );

    \I__3539\ : InMux
    port map (
            O => \N__27351\,
            I => \N__27348\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__27348\,
            I => \N__27345\
        );

    \I__3537\ : Span4Mux_v
    port map (
            O => \N__27345\,
            I => \N__27342\
        );

    \I__3536\ : Span4Mux_v
    port map (
            O => \N__27342\,
            I => \N__27339\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__27339\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_3
        );

    \I__3534\ : CascadeMux
    port map (
            O => \N__27336\,
            I => \N__27333\
        );

    \I__3533\ : InMux
    port map (
            O => \N__27333\,
            I => \N__27330\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__27330\,
            I => \N__27327\
        );

    \I__3531\ : Span12Mux_h
    port map (
            O => \N__27327\,
            I => \N__27324\
        );

    \I__3530\ : Odrv12
    port map (
            O => \N__27324\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_3
        );

    \I__3529\ : CascadeMux
    port map (
            O => \N__27321\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_3_cascade_\
        );

    \I__3528\ : InMux
    port map (
            O => \N__27318\,
            I => \N__27315\
        );

    \I__3527\ : LocalMux
    port map (
            O => \N__27315\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_3\
        );

    \I__3526\ : InMux
    port map (
            O => \N__27312\,
            I => \N__27309\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__27309\,
            I => \N__27306\
        );

    \I__3524\ : Span12Mux_h
    port map (
            O => \N__27306\,
            I => \N__27303\
        );

    \I__3523\ : Odrv12
    port map (
            O => \N__27303\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_31
        );

    \I__3522\ : CascadeMux
    port map (
            O => \N__27300\,
            I => \N__27297\
        );

    \I__3521\ : InMux
    port map (
            O => \N__27297\,
            I => \N__27294\
        );

    \I__3520\ : LocalMux
    port map (
            O => \N__27294\,
            I => \N__27291\
        );

    \I__3519\ : Span4Mux_v
    port map (
            O => \N__27291\,
            I => \N__27288\
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__27288\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_31
        );

    \I__3517\ : InMux
    port map (
            O => \N__27285\,
            I => \N__27282\
        );

    \I__3516\ : LocalMux
    port map (
            O => \N__27282\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_18\
        );

    \I__3515\ : InMux
    port map (
            O => \N__27279\,
            I => \N__27276\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__27276\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_19\
        );

    \I__3513\ : InMux
    port map (
            O => \N__27273\,
            I => \N__27270\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__27270\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_16\
        );

    \I__3511\ : InMux
    port map (
            O => \N__27267\,
            I => \N__27264\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__27264\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_17\
        );

    \I__3509\ : InMux
    port map (
            O => \N__27261\,
            I => \N__27258\
        );

    \I__3508\ : LocalMux
    port map (
            O => \N__27258\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_11\
        );

    \I__3507\ : InMux
    port map (
            O => \N__27255\,
            I => \N__27252\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__27252\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_8\
        );

    \I__3505\ : InMux
    port map (
            O => \N__27249\,
            I => \N__27246\
        );

    \I__3504\ : LocalMux
    port map (
            O => \N__27246\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_9\
        );

    \I__3503\ : InMux
    port map (
            O => \N__27243\,
            I => \N__27240\
        );

    \I__3502\ : LocalMux
    port map (
            O => \N__27240\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_10\
        );

    \I__3501\ : CEMux
    port map (
            O => \N__27237\,
            I => \N__27232\
        );

    \I__3500\ : CEMux
    port map (
            O => \N__27236\,
            I => \N__27229\
        );

    \I__3499\ : CEMux
    port map (
            O => \N__27235\,
            I => \N__27226\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__27232\,
            I => \N__27223\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__27229\,
            I => \N__27220\
        );

    \I__3496\ : LocalMux
    port map (
            O => \N__27226\,
            I => \N__27217\
        );

    \I__3495\ : Odrv4
    port map (
            O => \N__27223\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i\
        );

    \I__3494\ : Odrv4
    port map (
            O => \N__27220\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i\
        );

    \I__3493\ : Odrv4
    port map (
            O => \N__27217\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i\
        );

    \I__3492\ : InMux
    port map (
            O => \N__27210\,
            I => \N__27204\
        );

    \I__3491\ : InMux
    port map (
            O => \N__27209\,
            I => \N__27199\
        );

    \I__3490\ : InMux
    port map (
            O => \N__27208\,
            I => \N__27199\
        );

    \I__3489\ : InMux
    port map (
            O => \N__27207\,
            I => \N__27196\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__27204\,
            I => \N__27190\
        );

    \I__3487\ : LocalMux
    port map (
            O => \N__27199\,
            I => \N__27187\
        );

    \I__3486\ : LocalMux
    port map (
            O => \N__27196\,
            I => \N__27184\
        );

    \I__3485\ : InMux
    port map (
            O => \N__27195\,
            I => \N__27177\
        );

    \I__3484\ : InMux
    port map (
            O => \N__27194\,
            I => \N__27177\
        );

    \I__3483\ : InMux
    port map (
            O => \N__27193\,
            I => \N__27174\
        );

    \I__3482\ : Span4Mux_v
    port map (
            O => \N__27190\,
            I => \N__27169\
        );

    \I__3481\ : Span4Mux_v
    port map (
            O => \N__27187\,
            I => \N__27169\
        );

    \I__3480\ : Span4Mux_h
    port map (
            O => \N__27184\,
            I => \N__27166\
        );

    \I__3479\ : InMux
    port map (
            O => \N__27183\,
            I => \N__27161\
        );

    \I__3478\ : InMux
    port map (
            O => \N__27182\,
            I => \N__27161\
        );

    \I__3477\ : LocalMux
    port map (
            O => \N__27177\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__27174\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\
        );

    \I__3475\ : Odrv4
    port map (
            O => \N__27169\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\
        );

    \I__3474\ : Odrv4
    port map (
            O => \N__27166\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\
        );

    \I__3473\ : LocalMux
    port map (
            O => \N__27161\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\
        );

    \I__3472\ : CascadeMux
    port map (
            O => \N__27150\,
            I => \N__27128\
        );

    \I__3471\ : InMux
    port map (
            O => \N__27149\,
            I => \N__27125\
        );

    \I__3470\ : InMux
    port map (
            O => \N__27148\,
            I => \N__27114\
        );

    \I__3469\ : InMux
    port map (
            O => \N__27147\,
            I => \N__27114\
        );

    \I__3468\ : InMux
    port map (
            O => \N__27146\,
            I => \N__27114\
        );

    \I__3467\ : InMux
    port map (
            O => \N__27145\,
            I => \N__27114\
        );

    \I__3466\ : InMux
    port map (
            O => \N__27144\,
            I => \N__27114\
        );

    \I__3465\ : InMux
    port map (
            O => \N__27143\,
            I => \N__27111\
        );

    \I__3464\ : InMux
    port map (
            O => \N__27142\,
            I => \N__27108\
        );

    \I__3463\ : InMux
    port map (
            O => \N__27141\,
            I => \N__27098\
        );

    \I__3462\ : InMux
    port map (
            O => \N__27140\,
            I => \N__27098\
        );

    \I__3461\ : InMux
    port map (
            O => \N__27139\,
            I => \N__27098\
        );

    \I__3460\ : InMux
    port map (
            O => \N__27138\,
            I => \N__27098\
        );

    \I__3459\ : InMux
    port map (
            O => \N__27137\,
            I => \N__27083\
        );

    \I__3458\ : InMux
    port map (
            O => \N__27136\,
            I => \N__27083\
        );

    \I__3457\ : InMux
    port map (
            O => \N__27135\,
            I => \N__27083\
        );

    \I__3456\ : InMux
    port map (
            O => \N__27134\,
            I => \N__27083\
        );

    \I__3455\ : InMux
    port map (
            O => \N__27133\,
            I => \N__27083\
        );

    \I__3454\ : InMux
    port map (
            O => \N__27132\,
            I => \N__27083\
        );

    \I__3453\ : InMux
    port map (
            O => \N__27131\,
            I => \N__27083\
        );

    \I__3452\ : InMux
    port map (
            O => \N__27128\,
            I => \N__27080\
        );

    \I__3451\ : LocalMux
    port map (
            O => \N__27125\,
            I => \N__27073\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__27114\,
            I => \N__27073\
        );

    \I__3449\ : LocalMux
    port map (
            O => \N__27111\,
            I => \N__27073\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__27108\,
            I => \N__27070\
        );

    \I__3447\ : InMux
    port map (
            O => \N__27107\,
            I => \N__27065\
        );

    \I__3446\ : LocalMux
    port map (
            O => \N__27098\,
            I => \N__27060\
        );

    \I__3445\ : LocalMux
    port map (
            O => \N__27083\,
            I => \N__27060\
        );

    \I__3444\ : LocalMux
    port map (
            O => \N__27080\,
            I => \N__27055\
        );

    \I__3443\ : Span4Mux_h
    port map (
            O => \N__27073\,
            I => \N__27055\
        );

    \I__3442\ : Span4Mux_h
    port map (
            O => \N__27070\,
            I => \N__27052\
        );

    \I__3441\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27047\
        );

    \I__3440\ : InMux
    port map (
            O => \N__27068\,
            I => \N__27047\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__27065\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\
        );

    \I__3438\ : Odrv12
    port map (
            O => \N__27060\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\
        );

    \I__3437\ : Odrv4
    port map (
            O => \N__27055\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\
        );

    \I__3436\ : Odrv4
    port map (
            O => \N__27052\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\
        );

    \I__3435\ : LocalMux
    port map (
            O => \N__27047\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\
        );

    \I__3434\ : CascadeMux
    port map (
            O => \N__27036\,
            I => \N__27032\
        );

    \I__3433\ : InMux
    port map (
            O => \N__27035\,
            I => \N__27027\
        );

    \I__3432\ : InMux
    port map (
            O => \N__27032\,
            I => \N__27027\
        );

    \I__3431\ : LocalMux
    port map (
            O => \N__27027\,
            I => \N__27024\
        );

    \I__3430\ : Odrv12
    port map (
            O => \N__27024\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_391\
        );

    \I__3429\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27018\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__27018\,
            I => \N__27015\
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__27015\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_8\
        );

    \I__3426\ : InMux
    port map (
            O => \N__27012\,
            I => \N__27009\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__27009\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_11\
        );

    \I__3424\ : InMux
    port map (
            O => \N__27006\,
            I => \N__27003\
        );

    \I__3423\ : LocalMux
    port map (
            O => \N__27003\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_12\
        );

    \I__3422\ : InMux
    port map (
            O => \N__27000\,
            I => \N__26991\
        );

    \I__3421\ : InMux
    port map (
            O => \N__26999\,
            I => \N__26983\
        );

    \I__3420\ : InMux
    port map (
            O => \N__26998\,
            I => \N__26983\
        );

    \I__3419\ : InMux
    port map (
            O => \N__26997\,
            I => \N__26983\
        );

    \I__3418\ : InMux
    port map (
            O => \N__26996\,
            I => \N__26977\
        );

    \I__3417\ : InMux
    port map (
            O => \N__26995\,
            I => \N__26977\
        );

    \I__3416\ : InMux
    port map (
            O => \N__26994\,
            I => \N__26973\
        );

    \I__3415\ : LocalMux
    port map (
            O => \N__26991\,
            I => \N__26970\
        );

    \I__3414\ : InMux
    port map (
            O => \N__26990\,
            I => \N__26967\
        );

    \I__3413\ : LocalMux
    port map (
            O => \N__26983\,
            I => \N__26964\
        );

    \I__3412\ : InMux
    port map (
            O => \N__26982\,
            I => \N__26961\
        );

    \I__3411\ : LocalMux
    port map (
            O => \N__26977\,
            I => \N__26958\
        );

    \I__3410\ : InMux
    port map (
            O => \N__26976\,
            I => \N__26955\
        );

    \I__3409\ : LocalMux
    port map (
            O => \N__26973\,
            I => \N__26948\
        );

    \I__3408\ : Span4Mux_v
    port map (
            O => \N__26970\,
            I => \N__26948\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26948\
        );

    \I__3406\ : Odrv4
    port map (
            O => \N__26964\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\
        );

    \I__3405\ : LocalMux
    port map (
            O => \N__26961\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\
        );

    \I__3404\ : Odrv12
    port map (
            O => \N__26958\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\
        );

    \I__3403\ : LocalMux
    port map (
            O => \N__26955\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\
        );

    \I__3402\ : Odrv4
    port map (
            O => \N__26948\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\
        );

    \I__3401\ : InMux
    port map (
            O => \N__26937\,
            I => \N__26934\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__26934\,
            I => \N__26928\
        );

    \I__3399\ : InMux
    port map (
            O => \N__26933\,
            I => \N__26925\
        );

    \I__3398\ : InMux
    port map (
            O => \N__26932\,
            I => \N__26920\
        );

    \I__3397\ : InMux
    port map (
            O => \N__26931\,
            I => \N__26917\
        );

    \I__3396\ : Span4Mux_h
    port map (
            O => \N__26928\,
            I => \N__26914\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__26925\,
            I => \N__26911\
        );

    \I__3394\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26906\
        );

    \I__3393\ : InMux
    port map (
            O => \N__26923\,
            I => \N__26906\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__26920\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\
        );

    \I__3391\ : LocalMux
    port map (
            O => \N__26917\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\
        );

    \I__3390\ : Odrv4
    port map (
            O => \N__26914\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\
        );

    \I__3389\ : Odrv12
    port map (
            O => \N__26911\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\
        );

    \I__3388\ : LocalMux
    port map (
            O => \N__26906\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\
        );

    \I__3387\ : CascadeMux
    port map (
            O => \N__26895\,
            I => \N__26890\
        );

    \I__3386\ : InMux
    port map (
            O => \N__26894\,
            I => \N__26883\
        );

    \I__3385\ : InMux
    port map (
            O => \N__26893\,
            I => \N__26883\
        );

    \I__3384\ : InMux
    port map (
            O => \N__26890\,
            I => \N__26878\
        );

    \I__3383\ : InMux
    port map (
            O => \N__26889\,
            I => \N__26878\
        );

    \I__3382\ : InMux
    port map (
            O => \N__26888\,
            I => \N__26875\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__26883\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__26878\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i\
        );

    \I__3379\ : LocalMux
    port map (
            O => \N__26875\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i\
        );

    \I__3378\ : InMux
    port map (
            O => \N__26868\,
            I => \N__26865\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__26865\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_12\
        );

    \I__3376\ : InMux
    port map (
            O => \N__26862\,
            I => \N__26859\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__26859\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_13\
        );

    \I__3374\ : InMux
    port map (
            O => \N__26856\,
            I => \N__26853\
        );

    \I__3373\ : LocalMux
    port map (
            O => \N__26853\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_14\
        );

    \I__3372\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26847\
        );

    \I__3371\ : LocalMux
    port map (
            O => \N__26847\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_15\
        );

    \I__3370\ : InMux
    port map (
            O => \N__26844\,
            I => \N__26841\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__26841\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_14\
        );

    \I__3368\ : InMux
    port map (
            O => \N__26838\,
            I => \N__26835\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__26835\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_21\
        );

    \I__3366\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26829\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__26829\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_20\
        );

    \I__3364\ : InMux
    port map (
            O => \N__26826\,
            I => \N__26823\
        );

    \I__3363\ : LocalMux
    port map (
            O => \N__26823\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_9\
        );

    \I__3362\ : InMux
    port map (
            O => \N__26820\,
            I => \N__26817\
        );

    \I__3361\ : LocalMux
    port map (
            O => \N__26817\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_8\
        );

    \I__3360\ : InMux
    port map (
            O => \N__26814\,
            I => \N__26811\
        );

    \I__3359\ : LocalMux
    port map (
            O => \N__26811\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_10\
        );

    \I__3358\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26805\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__26805\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_22\
        );

    \I__3356\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26799\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__26799\,
            I => \N__26796\
        );

    \I__3354\ : Span4Mux_v
    port map (
            O => \N__26796\,
            I => \N__26793\
        );

    \I__3353\ : Odrv4
    port map (
            O => \N__26793\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.dout_op\
        );

    \I__3352\ : InMux
    port map (
            O => \N__26790\,
            I => \N__26787\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__26787\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_18\
        );

    \I__3350\ : InMux
    port map (
            O => \N__26784\,
            I => \N__26781\
        );

    \I__3349\ : LocalMux
    port map (
            O => \N__26781\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_19\
        );

    \I__3348\ : InMux
    port map (
            O => \N__26778\,
            I => \N__26775\
        );

    \I__3347\ : LocalMux
    port map (
            O => \N__26775\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_6\
        );

    \I__3346\ : InMux
    port map (
            O => \N__26772\,
            I => \N__26769\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__26769\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_17\
        );

    \I__3344\ : InMux
    port map (
            O => \N__26766\,
            I => \N__26763\
        );

    \I__3343\ : LocalMux
    port map (
            O => \N__26763\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_16\
        );

    \I__3342\ : InMux
    port map (
            O => \N__26760\,
            I => \N__26757\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__26757\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_15\
        );

    \I__3340\ : InMux
    port map (
            O => \N__26754\,
            I => \N__26751\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__26751\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_13\
        );

    \I__3338\ : CascadeMux
    port map (
            O => \N__26748\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_5_cascade_\
        );

    \I__3337\ : InMux
    port map (
            O => \N__26745\,
            I => \N__26742\
        );

    \I__3336\ : LocalMux
    port map (
            O => \N__26742\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_5\
        );

    \I__3335\ : InMux
    port map (
            O => \N__26739\,
            I => \N__26736\
        );

    \I__3334\ : LocalMux
    port map (
            O => \N__26736\,
            I => \N__26733\
        );

    \I__3333\ : Span4Mux_h
    port map (
            O => \N__26733\,
            I => \N__26730\
        );

    \I__3332\ : Sp12to4
    port map (
            O => \N__26730\,
            I => \N__26727\
        );

    \I__3331\ : Odrv12
    port map (
            O => \N__26727\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_5
        );

    \I__3330\ : CascadeMux
    port map (
            O => \N__26724\,
            I => \N__26721\
        );

    \I__3329\ : InMux
    port map (
            O => \N__26721\,
            I => \N__26718\
        );

    \I__3328\ : LocalMux
    port map (
            O => \N__26718\,
            I => \N__26715\
        );

    \I__3327\ : Span4Mux_v
    port map (
            O => \N__26715\,
            I => \N__26712\
        );

    \I__3326\ : Span4Mux_v
    port map (
            O => \N__26712\,
            I => \N__26709\
        );

    \I__3325\ : Odrv4
    port map (
            O => \N__26709\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_5
        );

    \I__3324\ : CascadeMux
    port map (
            O => \N__26706\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_5_cascade_\
        );

    \I__3323\ : InMux
    port map (
            O => \N__26703\,
            I => \N__26700\
        );

    \I__3322\ : LocalMux
    port map (
            O => \N__26700\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_5\
        );

    \I__3321\ : InMux
    port map (
            O => \N__26697\,
            I => \N__26694\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__26694\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6\
        );

    \I__3319\ : InMux
    port map (
            O => \N__26691\,
            I => \N__26688\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__26688\,
            I => \N__26685\
        );

    \I__3317\ : Odrv12
    port map (
            O => \N__26685\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_6\
        );

    \I__3316\ : InMux
    port map (
            O => \N__26682\,
            I => \N__26679\
        );

    \I__3315\ : LocalMux
    port map (
            O => \N__26679\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_5\
        );

    \I__3314\ : CascadeMux
    port map (
            O => \N__26676\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283_cascade_\
        );

    \I__3313\ : InMux
    port map (
            O => \N__26673\,
            I => \N__26669\
        );

    \I__3312\ : InMux
    port map (
            O => \N__26672\,
            I => \N__26666\
        );

    \I__3311\ : LocalMux
    port map (
            O => \N__26669\,
            I => \N__26662\
        );

    \I__3310\ : LocalMux
    port map (
            O => \N__26666\,
            I => \N__26659\
        );

    \I__3309\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26656\
        );

    \I__3308\ : Span4Mux_s3_v
    port map (
            O => \N__26662\,
            I => \N__26652\
        );

    \I__3307\ : Span4Mux_v
    port map (
            O => \N__26659\,
            I => \N__26647\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__26656\,
            I => \N__26647\
        );

    \I__3305\ : InMux
    port map (
            O => \N__26655\,
            I => \N__26644\
        );

    \I__3304\ : Odrv4
    port map (
            O => \N__26652\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__26647\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__26644\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0\
        );

    \I__3301\ : CEMux
    port map (
            O => \N__26637\,
            I => \N__26633\
        );

    \I__3300\ : CEMux
    port map (
            O => \N__26636\,
            I => \N__26630\
        );

    \I__3299\ : LocalMux
    port map (
            O => \N__26633\,
            I => \N__26627\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__26630\,
            I => \N__26624\
        );

    \I__3297\ : Span4Mux_h
    port map (
            O => \N__26627\,
            I => \N__26621\
        );

    \I__3296\ : Span4Mux_h
    port map (
            O => \N__26624\,
            I => \N__26618\
        );

    \I__3295\ : Odrv4
    port map (
            O => \N__26621\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0\
        );

    \I__3294\ : Odrv4
    port map (
            O => \N__26618\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0\
        );

    \I__3293\ : InMux
    port map (
            O => \N__26613\,
            I => \N__26610\
        );

    \I__3292\ : LocalMux
    port map (
            O => \N__26610\,
            I => \N__26607\
        );

    \I__3291\ : Span12Mux_v
    port map (
            O => \N__26607\,
            I => \N__26604\
        );

    \I__3290\ : Odrv12
    port map (
            O => \N__26604\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_1
        );

    \I__3289\ : CascadeMux
    port map (
            O => \N__26601\,
            I => \N__26598\
        );

    \I__3288\ : InMux
    port map (
            O => \N__26598\,
            I => \N__26595\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__26595\,
            I => \N__26592\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__26592\,
            I => \N__26589\
        );

    \I__3285\ : Odrv4
    port map (
            O => \N__26589\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_1
        );

    \I__3284\ : CascadeMux
    port map (
            O => \N__26586\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_1_cascade_\
        );

    \I__3283\ : InMux
    port map (
            O => \N__26583\,
            I => \N__26580\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__26580\,
            I => \N__26577\
        );

    \I__3281\ : Span4Mux_h
    port map (
            O => \N__26577\,
            I => \N__26574\
        );

    \I__3280\ : Odrv4
    port map (
            O => \N__26574\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_1
        );

    \I__3279\ : CascadeMux
    port map (
            O => \N__26571\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_1_cascade_\
        );

    \I__3278\ : CascadeMux
    port map (
            O => \N__26568\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_1_cascade_\
        );

    \I__3277\ : InMux
    port map (
            O => \N__26565\,
            I => \N__26562\
        );

    \I__3276\ : LocalMux
    port map (
            O => \N__26562\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_1\
        );

    \I__3275\ : InMux
    port map (
            O => \N__26559\,
            I => \N__26556\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__26556\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5\
        );

    \I__3273\ : InMux
    port map (
            O => \N__26553\,
            I => \N__26549\
        );

    \I__3272\ : InMux
    port map (
            O => \N__26552\,
            I => \N__26545\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__26549\,
            I => \N__26542\
        );

    \I__3270\ : InMux
    port map (
            O => \N__26548\,
            I => \N__26539\
        );

    \I__3269\ : LocalMux
    port map (
            O => \N__26545\,
            I => \N__26535\
        );

    \I__3268\ : Span4Mux_v
    port map (
            O => \N__26542\,
            I => \N__26530\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__26539\,
            I => \N__26530\
        );

    \I__3266\ : InMux
    port map (
            O => \N__26538\,
            I => \N__26527\
        );

    \I__3265\ : Span4Mux_h
    port map (
            O => \N__26535\,
            I => \N__26524\
        );

    \I__3264\ : Span4Mux_v
    port map (
            O => \N__26530\,
            I => \N__26519\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__26527\,
            I => \N__26519\
        );

    \I__3262\ : Odrv4
    port map (
            O => \N__26524\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0\
        );

    \I__3261\ : Odrv4
    port map (
            O => \N__26519\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0\
        );

    \I__3260\ : InMux
    port map (
            O => \N__26514\,
            I => \N__26511\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__26511\,
            I => \N__26506\
        );

    \I__3258\ : InMux
    port map (
            O => \N__26510\,
            I => \N__26503\
        );

    \I__3257\ : InMux
    port map (
            O => \N__26509\,
            I => \N__26499\
        );

    \I__3256\ : Span4Mux_h
    port map (
            O => \N__26506\,
            I => \N__26496\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__26503\,
            I => \N__26493\
        );

    \I__3254\ : InMux
    port map (
            O => \N__26502\,
            I => \N__26490\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__26499\,
            I => \N__26487\
        );

    \I__3252\ : Span4Mux_v
    port map (
            O => \N__26496\,
            I => \N__26482\
        );

    \I__3251\ : Span4Mux_h
    port map (
            O => \N__26493\,
            I => \N__26482\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__26490\,
            I => \N__26479\
        );

    \I__3249\ : Span4Mux_h
    port map (
            O => \N__26487\,
            I => \N__26472\
        );

    \I__3248\ : Span4Mux_v
    port map (
            O => \N__26482\,
            I => \N__26472\
        );

    \I__3247\ : Span4Mux_h
    port map (
            O => \N__26479\,
            I => \N__26472\
        );

    \I__3246\ : Odrv4
    port map (
            O => \N__26472\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_455_0\
        );

    \I__3245\ : InMux
    port map (
            O => \N__26469\,
            I => \N__26466\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__26466\,
            I => \N__26461\
        );

    \I__3243\ : InMux
    port map (
            O => \N__26465\,
            I => \N__26458\
        );

    \I__3242\ : InMux
    port map (
            O => \N__26464\,
            I => \N__26454\
        );

    \I__3241\ : Span4Mux_h
    port map (
            O => \N__26461\,
            I => \N__26451\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__26458\,
            I => \N__26448\
        );

    \I__3239\ : InMux
    port map (
            O => \N__26457\,
            I => \N__26445\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__26454\,
            I => \N__26442\
        );

    \I__3237\ : Span4Mux_v
    port map (
            O => \N__26451\,
            I => \N__26437\
        );

    \I__3236\ : Span4Mux_h
    port map (
            O => \N__26448\,
            I => \N__26437\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__26445\,
            I => \N__26434\
        );

    \I__3234\ : Span4Mux_h
    port map (
            O => \N__26442\,
            I => \N__26427\
        );

    \I__3233\ : Span4Mux_v
    port map (
            O => \N__26437\,
            I => \N__26427\
        );

    \I__3232\ : Span4Mux_h
    port map (
            O => \N__26434\,
            I => \N__26427\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__26427\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_454_0\
        );

    \I__3230\ : InMux
    port map (
            O => \N__26424\,
            I => \N__26421\
        );

    \I__3229\ : LocalMux
    port map (
            O => \N__26421\,
            I => \N__26416\
        );

    \I__3228\ : InMux
    port map (
            O => \N__26420\,
            I => \N__26413\
        );

    \I__3227\ : InMux
    port map (
            O => \N__26419\,
            I => \N__26409\
        );

    \I__3226\ : Span4Mux_v
    port map (
            O => \N__26416\,
            I => \N__26404\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__26413\,
            I => \N__26404\
        );

    \I__3224\ : InMux
    port map (
            O => \N__26412\,
            I => \N__26401\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__26409\,
            I => \N__26398\
        );

    \I__3222\ : Span4Mux_v
    port map (
            O => \N__26404\,
            I => \N__26393\
        );

    \I__3221\ : LocalMux
    port map (
            O => \N__26401\,
            I => \N__26393\
        );

    \I__3220\ : Span4Mux_v
    port map (
            O => \N__26398\,
            I => \N__26388\
        );

    \I__3219\ : Span4Mux_v
    port map (
            O => \N__26393\,
            I => \N__26388\
        );

    \I__3218\ : Odrv4
    port map (
            O => \N__26388\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_453_0\
        );

    \I__3217\ : InMux
    port map (
            O => \N__26385\,
            I => \N__26381\
        );

    \I__3216\ : InMux
    port map (
            O => \N__26384\,
            I => \N__26377\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__26381\,
            I => \N__26373\
        );

    \I__3214\ : InMux
    port map (
            O => \N__26380\,
            I => \N__26370\
        );

    \I__3213\ : LocalMux
    port map (
            O => \N__26377\,
            I => \N__26367\
        );

    \I__3212\ : InMux
    port map (
            O => \N__26376\,
            I => \N__26364\
        );

    \I__3211\ : Span4Mux_h
    port map (
            O => \N__26373\,
            I => \N__26361\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__26370\,
            I => \N__26358\
        );

    \I__3209\ : Span4Mux_h
    port map (
            O => \N__26367\,
            I => \N__26355\
        );

    \I__3208\ : LocalMux
    port map (
            O => \N__26364\,
            I => \N__26352\
        );

    \I__3207\ : Span4Mux_v
    port map (
            O => \N__26361\,
            I => \N__26343\
        );

    \I__3206\ : Span4Mux_h
    port map (
            O => \N__26358\,
            I => \N__26343\
        );

    \I__3205\ : Span4Mux_v
    port map (
            O => \N__26355\,
            I => \N__26343\
        );

    \I__3204\ : Span4Mux_h
    port map (
            O => \N__26352\,
            I => \N__26343\
        );

    \I__3203\ : Odrv4
    port map (
            O => \N__26343\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_463_0\
        );

    \I__3202\ : CascadeMux
    port map (
            O => \N__26340\,
            I => \N__26321\
        );

    \I__3201\ : CascadeMux
    port map (
            O => \N__26339\,
            I => \N__26317\
        );

    \I__3200\ : CascadeMux
    port map (
            O => \N__26338\,
            I => \N__26313\
        );

    \I__3199\ : InMux
    port map (
            O => \N__26337\,
            I => \N__26307\
        );

    \I__3198\ : InMux
    port map (
            O => \N__26336\,
            I => \N__26307\
        );

    \I__3197\ : InMux
    port map (
            O => \N__26335\,
            I => \N__26302\
        );

    \I__3196\ : InMux
    port map (
            O => \N__26334\,
            I => \N__26302\
        );

    \I__3195\ : InMux
    port map (
            O => \N__26333\,
            I => \N__26297\
        );

    \I__3194\ : InMux
    port map (
            O => \N__26332\,
            I => \N__26297\
        );

    \I__3193\ : CascadeMux
    port map (
            O => \N__26331\,
            I => \N__26293\
        );

    \I__3192\ : CascadeMux
    port map (
            O => \N__26330\,
            I => \N__26289\
        );

    \I__3191\ : CascadeMux
    port map (
            O => \N__26329\,
            I => \N__26285\
        );

    \I__3190\ : CascadeMux
    port map (
            O => \N__26328\,
            I => \N__26281\
        );

    \I__3189\ : CascadeMux
    port map (
            O => \N__26327\,
            I => \N__26278\
        );

    \I__3188\ : CascadeMux
    port map (
            O => \N__26326\,
            I => \N__26273\
        );

    \I__3187\ : CascadeMux
    port map (
            O => \N__26325\,
            I => \N__26268\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__26324\,
            I => \N__26265\
        );

    \I__3185\ : InMux
    port map (
            O => \N__26321\,
            I => \N__26258\
        );

    \I__3184\ : InMux
    port map (
            O => \N__26320\,
            I => \N__26258\
        );

    \I__3183\ : InMux
    port map (
            O => \N__26317\,
            I => \N__26249\
        );

    \I__3182\ : InMux
    port map (
            O => \N__26316\,
            I => \N__26249\
        );

    \I__3181\ : InMux
    port map (
            O => \N__26313\,
            I => \N__26249\
        );

    \I__3180\ : InMux
    port map (
            O => \N__26312\,
            I => \N__26249\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__26307\,
            I => \N__26246\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__26302\,
            I => \N__26241\
        );

    \I__3177\ : LocalMux
    port map (
            O => \N__26297\,
            I => \N__26241\
        );

    \I__3176\ : InMux
    port map (
            O => \N__26296\,
            I => \N__26230\
        );

    \I__3175\ : InMux
    port map (
            O => \N__26293\,
            I => \N__26230\
        );

    \I__3174\ : InMux
    port map (
            O => \N__26292\,
            I => \N__26230\
        );

    \I__3173\ : InMux
    port map (
            O => \N__26289\,
            I => \N__26230\
        );

    \I__3172\ : InMux
    port map (
            O => \N__26288\,
            I => \N__26230\
        );

    \I__3171\ : InMux
    port map (
            O => \N__26285\,
            I => \N__26213\
        );

    \I__3170\ : InMux
    port map (
            O => \N__26284\,
            I => \N__26213\
        );

    \I__3169\ : InMux
    port map (
            O => \N__26281\,
            I => \N__26213\
        );

    \I__3168\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26213\
        );

    \I__3167\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26213\
        );

    \I__3166\ : InMux
    port map (
            O => \N__26276\,
            I => \N__26213\
        );

    \I__3165\ : InMux
    port map (
            O => \N__26273\,
            I => \N__26213\
        );

    \I__3164\ : InMux
    port map (
            O => \N__26272\,
            I => \N__26213\
        );

    \I__3163\ : InMux
    port map (
            O => \N__26271\,
            I => \N__26202\
        );

    \I__3162\ : InMux
    port map (
            O => \N__26268\,
            I => \N__26202\
        );

    \I__3161\ : InMux
    port map (
            O => \N__26265\,
            I => \N__26202\
        );

    \I__3160\ : InMux
    port map (
            O => \N__26264\,
            I => \N__26202\
        );

    \I__3159\ : InMux
    port map (
            O => \N__26263\,
            I => \N__26202\
        );

    \I__3158\ : LocalMux
    port map (
            O => \N__26258\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__26249\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3156\ : Odrv4
    port map (
            O => \N__26246\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3155\ : Odrv4
    port map (
            O => \N__26241\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__26230\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__26213\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__26202\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\
        );

    \I__3151\ : InMux
    port map (
            O => \N__26187\,
            I => \N__26183\
        );

    \I__3150\ : InMux
    port map (
            O => \N__26186\,
            I => \N__26179\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__26183\,
            I => \N__26176\
        );

    \I__3148\ : InMux
    port map (
            O => \N__26182\,
            I => \N__26173\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__26179\,
            I => \N__26170\
        );

    \I__3146\ : Span4Mux_h
    port map (
            O => \N__26176\,
            I => \N__26166\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__26173\,
            I => \N__26163\
        );

    \I__3144\ : Span4Mux_h
    port map (
            O => \N__26170\,
            I => \N__26160\
        );

    \I__3143\ : InMux
    port map (
            O => \N__26169\,
            I => \N__26157\
        );

    \I__3142\ : Span4Mux_v
    port map (
            O => \N__26166\,
            I => \N__26152\
        );

    \I__3141\ : Span4Mux_h
    port map (
            O => \N__26163\,
            I => \N__26152\
        );

    \I__3140\ : Span4Mux_v
    port map (
            O => \N__26160\,
            I => \N__26147\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__26157\,
            I => \N__26147\
        );

    \I__3138\ : Odrv4
    port map (
            O => \N__26152\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__26147\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0\
        );

    \I__3136\ : InMux
    port map (
            O => \N__26142\,
            I => \N__26139\
        );

    \I__3135\ : LocalMux
    port map (
            O => \N__26139\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_21\
        );

    \I__3134\ : InMux
    port map (
            O => \N__26136\,
            I => \N__26133\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__26133\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_20\
        );

    \I__3132\ : InMux
    port map (
            O => \N__26130\,
            I => \N__26127\
        );

    \I__3131\ : LocalMux
    port map (
            O => \N__26127\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_22\
        );

    \I__3130\ : InMux
    port map (
            O => \N__26124\,
            I => \N__26121\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__26121\,
            I => \N__26118\
        );

    \I__3128\ : Odrv12
    port map (
            O => \N__26118\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_op\
        );

    \I__3127\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26111\
        );

    \I__3126\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26108\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__26111\,
            I => \N__26105\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__26108\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0\
        );

    \I__3123\ : Odrv4
    port map (
            O => \N__26105\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0\
        );

    \I__3122\ : InMux
    port map (
            O => \N__26100\,
            I => \bfn_9_22_0_\
        );

    \I__3121\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26093\
        );

    \I__3120\ : InMux
    port map (
            O => \N__26096\,
            I => \N__26090\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__26093\,
            I => \N__26087\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__26090\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1\
        );

    \I__3117\ : Odrv12
    port map (
            O => \N__26087\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1\
        );

    \I__3116\ : InMux
    port map (
            O => \N__26082\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0\
        );

    \I__3115\ : InMux
    port map (
            O => \N__26079\,
            I => \N__26075\
        );

    \I__3114\ : InMux
    port map (
            O => \N__26078\,
            I => \N__26072\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__26075\,
            I => \N__26069\
        );

    \I__3112\ : LocalMux
    port map (
            O => \N__26072\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2\
        );

    \I__3111\ : Odrv4
    port map (
            O => \N__26069\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2\
        );

    \I__3110\ : InMux
    port map (
            O => \N__26064\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1\
        );

    \I__3109\ : InMux
    port map (
            O => \N__26061\,
            I => \N__26058\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__26058\,
            I => \N__26054\
        );

    \I__3107\ : InMux
    port map (
            O => \N__26057\,
            I => \N__26051\
        );

    \I__3106\ : Span4Mux_h
    port map (
            O => \N__26054\,
            I => \N__26048\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__26051\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__26048\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3\
        );

    \I__3103\ : InMux
    port map (
            O => \N__26043\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2\
        );

    \I__3102\ : InMux
    port map (
            O => \N__26040\,
            I => \N__26029\
        );

    \I__3101\ : InMux
    port map (
            O => \N__26039\,
            I => \N__26029\
        );

    \I__3100\ : InMux
    port map (
            O => \N__26038\,
            I => \N__26029\
        );

    \I__3099\ : InMux
    port map (
            O => \N__26037\,
            I => \N__26024\
        );

    \I__3098\ : InMux
    port map (
            O => \N__26036\,
            I => \N__26024\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__26029\,
            I => \N__26019\
        );

    \I__3096\ : LocalMux
    port map (
            O => \N__26024\,
            I => \N__26019\
        );

    \I__3095\ : Odrv4
    port map (
            O => \N__26019\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_391_i\
        );

    \I__3094\ : InMux
    port map (
            O => \N__26016\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_3\
        );

    \I__3093\ : InMux
    port map (
            O => \N__26013\,
            I => \N__26010\
        );

    \I__3092\ : LocalMux
    port map (
            O => \N__26010\,
            I => \N__26006\
        );

    \I__3091\ : InMux
    port map (
            O => \N__26009\,
            I => \N__26003\
        );

    \I__3090\ : Span4Mux_h
    port map (
            O => \N__26006\,
            I => \N__26000\
        );

    \I__3089\ : LocalMux
    port map (
            O => \N__26003\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4\
        );

    \I__3088\ : Odrv4
    port map (
            O => \N__26000\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4\
        );

    \I__3087\ : InMux
    port map (
            O => \N__25995\,
            I => \N__25992\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__25992\,
            I => \N__25987\
        );

    \I__3085\ : InMux
    port map (
            O => \N__25991\,
            I => \N__25984\
        );

    \I__3084\ : InMux
    port map (
            O => \N__25990\,
            I => \N__25981\
        );

    \I__3083\ : Span4Mux_h
    port map (
            O => \N__25987\,
            I => \N__25978\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__25984\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1\
        );

    \I__3081\ : LocalMux
    port map (
            O => \N__25981\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1\
        );

    \I__3080\ : Odrv4
    port map (
            O => \N__25978\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1\
        );

    \I__3079\ : InMux
    port map (
            O => \N__25971\,
            I => \N__25968\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__25968\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_CO\
        );

    \I__3077\ : InMux
    port map (
            O => \N__25965\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0\
        );

    \I__3076\ : InMux
    port map (
            O => \N__25962\,
            I => \N__25959\
        );

    \I__3075\ : LocalMux
    port map (
            O => \N__25959\,
            I => \N__25954\
        );

    \I__3074\ : InMux
    port map (
            O => \N__25958\,
            I => \N__25951\
        );

    \I__3073\ : InMux
    port map (
            O => \N__25957\,
            I => \N__25948\
        );

    \I__3072\ : Span4Mux_h
    port map (
            O => \N__25954\,
            I => \N__25945\
        );

    \I__3071\ : LocalMux
    port map (
            O => \N__25951\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__25948\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2\
        );

    \I__3069\ : Odrv4
    port map (
            O => \N__25945\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2\
        );

    \I__3068\ : CascadeMux
    port map (
            O => \N__25938\,
            I => \N__25935\
        );

    \I__3067\ : InMux
    port map (
            O => \N__25935\,
            I => \N__25932\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__25932\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_CO\
        );

    \I__3065\ : InMux
    port map (
            O => \N__25929\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1\
        );

    \I__3064\ : InMux
    port map (
            O => \N__25926\,
            I => \N__25922\
        );

    \I__3063\ : CascadeMux
    port map (
            O => \N__25925\,
            I => \N__25919\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__25922\,
            I => \N__25915\
        );

    \I__3061\ : InMux
    port map (
            O => \N__25919\,
            I => \N__25912\
        );

    \I__3060\ : InMux
    port map (
            O => \N__25918\,
            I => \N__25909\
        );

    \I__3059\ : Span4Mux_v
    port map (
            O => \N__25915\,
            I => \N__25906\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__25912\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3\
        );

    \I__3057\ : LocalMux
    port map (
            O => \N__25909\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3\
        );

    \I__3056\ : Odrv4
    port map (
            O => \N__25906\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3\
        );

    \I__3055\ : InMux
    port map (
            O => \N__25899\,
            I => \N__25896\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__25896\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_CO\
        );

    \I__3053\ : InMux
    port map (
            O => \N__25893\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2\
        );

    \I__3052\ : InMux
    port map (
            O => \N__25890\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_3\
        );

    \I__3051\ : CascadeMux
    port map (
            O => \N__25887\,
            I => \N__25884\
        );

    \I__3050\ : InMux
    port map (
            O => \N__25884\,
            I => \N__25880\
        );

    \I__3049\ : InMux
    port map (
            O => \N__25883\,
            I => \N__25877\
        );

    \I__3048\ : LocalMux
    port map (
            O => \N__25880\,
            I => \N__25874\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__25877\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4\
        );

    \I__3046\ : Odrv4
    port map (
            O => \N__25874\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4\
        );

    \I__3045\ : InMux
    port map (
            O => \N__25869\,
            I => \N__25866\
        );

    \I__3044\ : LocalMux
    port map (
            O => \N__25866\,
            I => \N__25863\
        );

    \I__3043\ : Span4Mux_v
    port map (
            O => \N__25863\,
            I => \N__25860\
        );

    \I__3042\ : Odrv4
    port map (
            O => \N__25860\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_a2_1_0\
        );

    \I__3041\ : InMux
    port map (
            O => \N__25857\,
            I => \N__25854\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__25854\,
            I => \N__25851\
        );

    \I__3039\ : Span4Mux_h
    port map (
            O => \N__25851\,
            I => \N__25848\
        );

    \I__3038\ : Odrv4
    port map (
            O => \N__25848\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_3\
        );

    \I__3037\ : CascadeMux
    port map (
            O => \N__25845\,
            I => \N__25841\
        );

    \I__3036\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25835\
        );

    \I__3035\ : InMux
    port map (
            O => \N__25841\,
            I => \N__25832\
        );

    \I__3034\ : InMux
    port map (
            O => \N__25840\,
            I => \N__25829\
        );

    \I__3033\ : InMux
    port map (
            O => \N__25839\,
            I => \N__25824\
        );

    \I__3032\ : InMux
    port map (
            O => \N__25838\,
            I => \N__25824\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__25835\,
            I => \N__25821\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__25832\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__25829\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14\
        );

    \I__3028\ : LocalMux
    port map (
            O => \N__25824\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14\
        );

    \I__3027\ : Odrv12
    port map (
            O => \N__25821\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14\
        );

    \I__3026\ : CascadeMux
    port map (
            O => \N__25812\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_cascade_\
        );

    \I__3025\ : InMux
    port map (
            O => \N__25809\,
            I => \N__25805\
        );

    \I__3024\ : InMux
    port map (
            O => \N__25808\,
            I => \N__25799\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__25805\,
            I => \N__25796\
        );

    \I__3022\ : InMux
    port map (
            O => \N__25804\,
            I => \N__25789\
        );

    \I__3021\ : InMux
    port map (
            O => \N__25803\,
            I => \N__25789\
        );

    \I__3020\ : InMux
    port map (
            O => \N__25802\,
            I => \N__25789\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__25799\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6\
        );

    \I__3018\ : Odrv4
    port map (
            O => \N__25796\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__25789\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6\
        );

    \I__3016\ : CascadeMux
    port map (
            O => \N__25782\,
            I => \N__25775\
        );

    \I__3015\ : InMux
    port map (
            O => \N__25781\,
            I => \N__25766\
        );

    \I__3014\ : InMux
    port map (
            O => \N__25780\,
            I => \N__25766\
        );

    \I__3013\ : InMux
    port map (
            O => \N__25779\,
            I => \N__25766\
        );

    \I__3012\ : InMux
    port map (
            O => \N__25778\,
            I => \N__25766\
        );

    \I__3011\ : InMux
    port map (
            O => \N__25775\,
            I => \N__25763\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__25766\,
            I => \N__25760\
        );

    \I__3009\ : LocalMux
    port map (
            O => \N__25763\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0\
        );

    \I__3008\ : Odrv4
    port map (
            O => \N__25760\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0\
        );

    \I__3007\ : InMux
    port map (
            O => \N__25755\,
            I => \N__25752\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__25752\,
            I => \N__25748\
        );

    \I__3005\ : CascadeMux
    port map (
            O => \N__25751\,
            I => \N__25737\
        );

    \I__3004\ : Span4Mux_v
    port map (
            O => \N__25748\,
            I => \N__25733\
        );

    \I__3003\ : InMux
    port map (
            O => \N__25747\,
            I => \N__25716\
        );

    \I__3002\ : InMux
    port map (
            O => \N__25746\,
            I => \N__25716\
        );

    \I__3001\ : InMux
    port map (
            O => \N__25745\,
            I => \N__25716\
        );

    \I__3000\ : InMux
    port map (
            O => \N__25744\,
            I => \N__25716\
        );

    \I__2999\ : InMux
    port map (
            O => \N__25743\,
            I => \N__25716\
        );

    \I__2998\ : InMux
    port map (
            O => \N__25742\,
            I => \N__25716\
        );

    \I__2997\ : InMux
    port map (
            O => \N__25741\,
            I => \N__25716\
        );

    \I__2996\ : InMux
    port map (
            O => \N__25740\,
            I => \N__25716\
        );

    \I__2995\ : InMux
    port map (
            O => \N__25737\,
            I => \N__25711\
        );

    \I__2994\ : InMux
    port map (
            O => \N__25736\,
            I => \N__25711\
        );

    \I__2993\ : Odrv4
    port map (
            O => \N__25733\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10\
        );

    \I__2992\ : LocalMux
    port map (
            O => \N__25716\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10\
        );

    \I__2991\ : LocalMux
    port map (
            O => \N__25711\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10\
        );

    \I__2990\ : CascadeMux
    port map (
            O => \N__25704\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.csb_u_i_a2_0_0_cascade_\
        );

    \I__2989\ : CascadeMux
    port map (
            O => \N__25701\,
            I => \N__25698\
        );

    \I__2988\ : InMux
    port map (
            O => \N__25698\,
            I => \N__25690\
        );

    \I__2987\ : InMux
    port map (
            O => \N__25697\,
            I => \N__25690\
        );

    \I__2986\ : CascadeMux
    port map (
            O => \N__25696\,
            I => \N__25687\
        );

    \I__2985\ : InMux
    port map (
            O => \N__25695\,
            I => \N__25683\
        );

    \I__2984\ : LocalMux
    port map (
            O => \N__25690\,
            I => \N__25678\
        );

    \I__2983\ : InMux
    port map (
            O => \N__25687\,
            I => \N__25673\
        );

    \I__2982\ : InMux
    port map (
            O => \N__25686\,
            I => \N__25673\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__25683\,
            I => \N__25670\
        );

    \I__2980\ : InMux
    port map (
            O => \N__25682\,
            I => \N__25665\
        );

    \I__2979\ : InMux
    port map (
            O => \N__25681\,
            I => \N__25665\
        );

    \I__2978\ : Span4Mux_v
    port map (
            O => \N__25678\,
            I => \N__25660\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__25673\,
            I => \N__25660\
        );

    \I__2976\ : Odrv4
    port map (
            O => \N__25670\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__25665\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0\
        );

    \I__2974\ : Odrv4
    port map (
            O => \N__25660\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0\
        );

    \I__2973\ : IoInMux
    port map (
            O => \N__25653\,
            I => \N__25650\
        );

    \I__2972\ : LocalMux
    port map (
            O => \N__25650\,
            I => \N__25647\
        );

    \I__2971\ : Span4Mux_s0_h
    port map (
            O => \N__25647\,
            I => \N__25644\
        );

    \I__2970\ : Sp12to4
    port map (
            O => \N__25644\,
            I => \N__25641\
        );

    \I__2969\ : Span12Mux_v
    port map (
            O => \N__25641\,
            I => \N__25638\
        );

    \I__2968\ : Odrv12
    port map (
            O => \N__25638\,
            I => \N_1822_0\
        );

    \I__2967\ : InMux
    port map (
            O => \N__25635\,
            I => \N__25632\
        );

    \I__2966\ : LocalMux
    port map (
            O => \N__25632\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.csb_u_i_a2_0\
        );

    \I__2965\ : InMux
    port map (
            O => \N__25629\,
            I => \N__25623\
        );

    \I__2964\ : InMux
    port map (
            O => \N__25628\,
            I => \N__25618\
        );

    \I__2963\ : InMux
    port map (
            O => \N__25627\,
            I => \N__25618\
        );

    \I__2962\ : InMux
    port map (
            O => \N__25626\,
            I => \N__25613\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__25623\,
            I => \N__25608\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__25618\,
            I => \N__25608\
        );

    \I__2959\ : InMux
    port map (
            O => \N__25617\,
            I => \N__25605\
        );

    \I__2958\ : InMux
    port map (
            O => \N__25616\,
            I => \N__25602\
        );

    \I__2957\ : LocalMux
    port map (
            O => \N__25613\,
            I => \N__25595\
        );

    \I__2956\ : Span4Mux_v
    port map (
            O => \N__25608\,
            I => \N__25595\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__25605\,
            I => \N__25595\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__25602\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0\
        );

    \I__2953\ : Odrv4
    port map (
            O => \N__25595\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0\
        );

    \I__2952\ : InMux
    port map (
            O => \N__25590\,
            I => \N__25587\
        );

    \I__2951\ : LocalMux
    port map (
            O => \N__25587\,
            I => \N__25584\
        );

    \I__2950\ : Span4Mux_h
    port map (
            O => \N__25584\,
            I => \N__25578\
        );

    \I__2949\ : InMux
    port map (
            O => \N__25583\,
            I => \N__25574\
        );

    \I__2948\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25569\
        );

    \I__2947\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25569\
        );

    \I__2946\ : Span4Mux_v
    port map (
            O => \N__25578\,
            I => \N__25566\
        );

    \I__2945\ : InMux
    port map (
            O => \N__25577\,
            I => \N__25563\
        );

    \I__2944\ : LocalMux
    port map (
            O => \N__25574\,
            I => \N__25560\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__25569\,
            I => \N__25557\
        );

    \I__2942\ : Span4Mux_v
    port map (
            O => \N__25566\,
            I => \N__25554\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__25563\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0\
        );

    \I__2940\ : Odrv4
    port map (
            O => \N__25560\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0\
        );

    \I__2939\ : Odrv12
    port map (
            O => \N__25557\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0\
        );

    \I__2938\ : Odrv4
    port map (
            O => \N__25554\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0\
        );

    \I__2937\ : InMux
    port map (
            O => \N__25545\,
            I => \N__25542\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__25542\,
            I => \N__25539\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__25539\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_CO\
        );

    \I__2934\ : InMux
    port map (
            O => \N__25536\,
            I => \N__25531\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__25535\,
            I => \N__25527\
        );

    \I__2932\ : CascadeMux
    port map (
            O => \N__25534\,
            I => \N__25524\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__25531\,
            I => \N__25520\
        );

    \I__2930\ : InMux
    port map (
            O => \N__25530\,
            I => \N__25517\
        );

    \I__2929\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25514\
        );

    \I__2928\ : InMux
    port map (
            O => \N__25524\,
            I => \N__25509\
        );

    \I__2927\ : InMux
    port map (
            O => \N__25523\,
            I => \N__25509\
        );

    \I__2926\ : Sp12to4
    port map (
            O => \N__25520\,
            I => \N__25506\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__25517\,
            I => \N__25503\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__25514\,
            I => \N__25496\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__25509\,
            I => \N__25496\
        );

    \I__2922\ : Span12Mux_v
    port map (
            O => \N__25506\,
            I => \N__25496\
        );

    \I__2921\ : Odrv4
    port map (
            O => \N__25503\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i\
        );

    \I__2920\ : Odrv12
    port map (
            O => \N__25496\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__25491\,
            I => \N__25488\
        );

    \I__2918\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25484\
        );

    \I__2917\ : InMux
    port map (
            O => \N__25487\,
            I => \N__25480\
        );

    \I__2916\ : LocalMux
    port map (
            O => \N__25484\,
            I => \N__25477\
        );

    \I__2915\ : InMux
    port map (
            O => \N__25483\,
            I => \N__25474\
        );

    \I__2914\ : LocalMux
    port map (
            O => \N__25480\,
            I => \N__25471\
        );

    \I__2913\ : Span4Mux_h
    port map (
            O => \N__25477\,
            I => \N__25468\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__25474\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__25471\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1\
        );

    \I__2910\ : Odrv4
    port map (
            O => \N__25468\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1\
        );

    \I__2909\ : InMux
    port map (
            O => \N__25461\,
            I => \N__25453\
        );

    \I__2908\ : InMux
    port map (
            O => \N__25460\,
            I => \N__25453\
        );

    \I__2907\ : InMux
    port map (
            O => \N__25459\,
            I => \N__25448\
        );

    \I__2906\ : InMux
    port map (
            O => \N__25458\,
            I => \N__25448\
        );

    \I__2905\ : LocalMux
    port map (
            O => \N__25453\,
            I => \N__25444\
        );

    \I__2904\ : LocalMux
    port map (
            O => \N__25448\,
            I => \N__25441\
        );

    \I__2903\ : InMux
    port map (
            O => \N__25447\,
            I => \N__25437\
        );

    \I__2902\ : Span4Mux_v
    port map (
            O => \N__25444\,
            I => \N__25432\
        );

    \I__2901\ : Span4Mux_v
    port map (
            O => \N__25441\,
            I => \N__25432\
        );

    \I__2900\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25429\
        );

    \I__2899\ : LocalMux
    port map (
            O => \N__25437\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0\
        );

    \I__2898\ : Odrv4
    port map (
            O => \N__25432\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__25429\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0\
        );

    \I__2896\ : IoInMux
    port map (
            O => \N__25422\,
            I => \N__25419\
        );

    \I__2895\ : LocalMux
    port map (
            O => \N__25419\,
            I => \N__25416\
        );

    \I__2894\ : IoSpan4Mux
    port map (
            O => \N__25416\,
            I => \N__25413\
        );

    \I__2893\ : Span4Mux_s3_h
    port map (
            O => \N__25413\,
            I => \N__25410\
        );

    \I__2892\ : Span4Mux_h
    port map (
            O => \N__25410\,
            I => \N__25407\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__25407\,
            I => \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_iZ0\
        );

    \I__2890\ : CascadeMux
    port map (
            O => \N__25404\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_596_cascade_\
        );

    \I__2889\ : InMux
    port map (
            O => \N__25401\,
            I => \N__25398\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__25398\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_597\
        );

    \I__2887\ : InMux
    port map (
            O => \N__25395\,
            I => \N__25392\
        );

    \I__2886\ : LocalMux
    port map (
            O => \N__25392\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_oZ0Z_26\
        );

    \I__2885\ : CascadeMux
    port map (
            O => \N__25389\,
            I => \cemf_module_64ch_ctrl_inst1.N_1615_cascade_\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__25386\,
            I => \N__25382\
        );

    \I__2883\ : CascadeMux
    port map (
            O => \N__25385\,
            I => \N__25379\
        );

    \I__2882\ : CascadeBuf
    port map (
            O => \N__25382\,
            I => \N__25376\
        );

    \I__2881\ : CascadeBuf
    port map (
            O => \N__25379\,
            I => \N__25373\
        );

    \I__2880\ : CascadeMux
    port map (
            O => \N__25376\,
            I => \N__25370\
        );

    \I__2879\ : CascadeMux
    port map (
            O => \N__25373\,
            I => \N__25367\
        );

    \I__2878\ : CascadeBuf
    port map (
            O => \N__25370\,
            I => \N__25364\
        );

    \I__2877\ : CascadeBuf
    port map (
            O => \N__25367\,
            I => \N__25361\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__25364\,
            I => \N__25358\
        );

    \I__2875\ : CascadeMux
    port map (
            O => \N__25361\,
            I => \N__25355\
        );

    \I__2874\ : CascadeBuf
    port map (
            O => \N__25358\,
            I => \N__25352\
        );

    \I__2873\ : CascadeBuf
    port map (
            O => \N__25355\,
            I => \N__25349\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__25352\,
            I => \N__25346\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__25349\,
            I => \N__25343\
        );

    \I__2870\ : CascadeBuf
    port map (
            O => \N__25346\,
            I => \N__25340\
        );

    \I__2869\ : CascadeBuf
    port map (
            O => \N__25343\,
            I => \N__25337\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__25340\,
            I => \N__25334\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__25337\,
            I => \N__25331\
        );

    \I__2866\ : CascadeBuf
    port map (
            O => \N__25334\,
            I => \N__25328\
        );

    \I__2865\ : CascadeBuf
    port map (
            O => \N__25331\,
            I => \N__25325\
        );

    \I__2864\ : CascadeMux
    port map (
            O => \N__25328\,
            I => \N__25322\
        );

    \I__2863\ : CascadeMux
    port map (
            O => \N__25325\,
            I => \N__25319\
        );

    \I__2862\ : CascadeBuf
    port map (
            O => \N__25322\,
            I => \N__25316\
        );

    \I__2861\ : CascadeBuf
    port map (
            O => \N__25319\,
            I => \N__25313\
        );

    \I__2860\ : CascadeMux
    port map (
            O => \N__25316\,
            I => \N__25310\
        );

    \I__2859\ : CascadeMux
    port map (
            O => \N__25313\,
            I => \N__25307\
        );

    \I__2858\ : CascadeBuf
    port map (
            O => \N__25310\,
            I => \N__25304\
        );

    \I__2857\ : CascadeBuf
    port map (
            O => \N__25307\,
            I => \N__25301\
        );

    \I__2856\ : CascadeMux
    port map (
            O => \N__25304\,
            I => \N__25298\
        );

    \I__2855\ : CascadeMux
    port map (
            O => \N__25301\,
            I => \N__25295\
        );

    \I__2854\ : InMux
    port map (
            O => \N__25298\,
            I => \N__25292\
        );

    \I__2853\ : InMux
    port map (
            O => \N__25295\,
            I => \N__25289\
        );

    \I__2852\ : LocalMux
    port map (
            O => \N__25292\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__25289\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0\
        );

    \I__2850\ : CascadeMux
    port map (
            O => \N__25284\,
            I => \N__25280\
        );

    \I__2849\ : CascadeMux
    port map (
            O => \N__25283\,
            I => \N__25277\
        );

    \I__2848\ : CascadeBuf
    port map (
            O => \N__25280\,
            I => \N__25274\
        );

    \I__2847\ : CascadeBuf
    port map (
            O => \N__25277\,
            I => \N__25271\
        );

    \I__2846\ : CascadeMux
    port map (
            O => \N__25274\,
            I => \N__25268\
        );

    \I__2845\ : CascadeMux
    port map (
            O => \N__25271\,
            I => \N__25265\
        );

    \I__2844\ : CascadeBuf
    port map (
            O => \N__25268\,
            I => \N__25262\
        );

    \I__2843\ : CascadeBuf
    port map (
            O => \N__25265\,
            I => \N__25259\
        );

    \I__2842\ : CascadeMux
    port map (
            O => \N__25262\,
            I => \N__25256\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__25259\,
            I => \N__25253\
        );

    \I__2840\ : CascadeBuf
    port map (
            O => \N__25256\,
            I => \N__25250\
        );

    \I__2839\ : CascadeBuf
    port map (
            O => \N__25253\,
            I => \N__25247\
        );

    \I__2838\ : CascadeMux
    port map (
            O => \N__25250\,
            I => \N__25244\
        );

    \I__2837\ : CascadeMux
    port map (
            O => \N__25247\,
            I => \N__25241\
        );

    \I__2836\ : CascadeBuf
    port map (
            O => \N__25244\,
            I => \N__25238\
        );

    \I__2835\ : CascadeBuf
    port map (
            O => \N__25241\,
            I => \N__25235\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__25238\,
            I => \N__25232\
        );

    \I__2833\ : CascadeMux
    port map (
            O => \N__25235\,
            I => \N__25229\
        );

    \I__2832\ : CascadeBuf
    port map (
            O => \N__25232\,
            I => \N__25226\
        );

    \I__2831\ : CascadeBuf
    port map (
            O => \N__25229\,
            I => \N__25223\
        );

    \I__2830\ : CascadeMux
    port map (
            O => \N__25226\,
            I => \N__25220\
        );

    \I__2829\ : CascadeMux
    port map (
            O => \N__25223\,
            I => \N__25217\
        );

    \I__2828\ : CascadeBuf
    port map (
            O => \N__25220\,
            I => \N__25214\
        );

    \I__2827\ : CascadeBuf
    port map (
            O => \N__25217\,
            I => \N__25211\
        );

    \I__2826\ : CascadeMux
    port map (
            O => \N__25214\,
            I => \N__25208\
        );

    \I__2825\ : CascadeMux
    port map (
            O => \N__25211\,
            I => \N__25205\
        );

    \I__2824\ : CascadeBuf
    port map (
            O => \N__25208\,
            I => \N__25202\
        );

    \I__2823\ : CascadeBuf
    port map (
            O => \N__25205\,
            I => \N__25199\
        );

    \I__2822\ : CascadeMux
    port map (
            O => \N__25202\,
            I => \N__25196\
        );

    \I__2821\ : CascadeMux
    port map (
            O => \N__25199\,
            I => \N__25193\
        );

    \I__2820\ : InMux
    port map (
            O => \N__25196\,
            I => \N__25190\
        );

    \I__2819\ : InMux
    port map (
            O => \N__25193\,
            I => \N__25187\
        );

    \I__2818\ : LocalMux
    port map (
            O => \N__25190\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0\
        );

    \I__2817\ : LocalMux
    port map (
            O => \N__25187\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0\
        );

    \I__2816\ : CascadeMux
    port map (
            O => \N__25182\,
            I => \N__25178\
        );

    \I__2815\ : CascadeMux
    port map (
            O => \N__25181\,
            I => \N__25175\
        );

    \I__2814\ : CascadeBuf
    port map (
            O => \N__25178\,
            I => \N__25172\
        );

    \I__2813\ : CascadeBuf
    port map (
            O => \N__25175\,
            I => \N__25169\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__25172\,
            I => \N__25166\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__25169\,
            I => \N__25163\
        );

    \I__2810\ : CascadeBuf
    port map (
            O => \N__25166\,
            I => \N__25160\
        );

    \I__2809\ : CascadeBuf
    port map (
            O => \N__25163\,
            I => \N__25157\
        );

    \I__2808\ : CascadeMux
    port map (
            O => \N__25160\,
            I => \N__25154\
        );

    \I__2807\ : CascadeMux
    port map (
            O => \N__25157\,
            I => \N__25151\
        );

    \I__2806\ : CascadeBuf
    port map (
            O => \N__25154\,
            I => \N__25148\
        );

    \I__2805\ : CascadeBuf
    port map (
            O => \N__25151\,
            I => \N__25145\
        );

    \I__2804\ : CascadeMux
    port map (
            O => \N__25148\,
            I => \N__25142\
        );

    \I__2803\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \N__25139\
        );

    \I__2802\ : CascadeBuf
    port map (
            O => \N__25142\,
            I => \N__25136\
        );

    \I__2801\ : CascadeBuf
    port map (
            O => \N__25139\,
            I => \N__25133\
        );

    \I__2800\ : CascadeMux
    port map (
            O => \N__25136\,
            I => \N__25130\
        );

    \I__2799\ : CascadeMux
    port map (
            O => \N__25133\,
            I => \N__25127\
        );

    \I__2798\ : CascadeBuf
    port map (
            O => \N__25130\,
            I => \N__25124\
        );

    \I__2797\ : CascadeBuf
    port map (
            O => \N__25127\,
            I => \N__25121\
        );

    \I__2796\ : CascadeMux
    port map (
            O => \N__25124\,
            I => \N__25118\
        );

    \I__2795\ : CascadeMux
    port map (
            O => \N__25121\,
            I => \N__25115\
        );

    \I__2794\ : CascadeBuf
    port map (
            O => \N__25118\,
            I => \N__25112\
        );

    \I__2793\ : CascadeBuf
    port map (
            O => \N__25115\,
            I => \N__25109\
        );

    \I__2792\ : CascadeMux
    port map (
            O => \N__25112\,
            I => \N__25106\
        );

    \I__2791\ : CascadeMux
    port map (
            O => \N__25109\,
            I => \N__25103\
        );

    \I__2790\ : CascadeBuf
    port map (
            O => \N__25106\,
            I => \N__25100\
        );

    \I__2789\ : CascadeBuf
    port map (
            O => \N__25103\,
            I => \N__25097\
        );

    \I__2788\ : CascadeMux
    port map (
            O => \N__25100\,
            I => \N__25094\
        );

    \I__2787\ : CascadeMux
    port map (
            O => \N__25097\,
            I => \N__25091\
        );

    \I__2786\ : InMux
    port map (
            O => \N__25094\,
            I => \N__25088\
        );

    \I__2785\ : InMux
    port map (
            O => \N__25091\,
            I => \N__25085\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__25088\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3\
        );

    \I__2783\ : LocalMux
    port map (
            O => \N__25085\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3\
        );

    \I__2782\ : InMux
    port map (
            O => \N__25080\,
            I => \N__25077\
        );

    \I__2781\ : LocalMux
    port map (
            O => \N__25077\,
            I => \N__25071\
        );

    \I__2780\ : InMux
    port map (
            O => \N__25076\,
            I => \N__25064\
        );

    \I__2779\ : InMux
    port map (
            O => \N__25075\,
            I => \N__25064\
        );

    \I__2778\ : InMux
    port map (
            O => \N__25074\,
            I => \N__25064\
        );

    \I__2777\ : Odrv12
    port map (
            O => \N__25071\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9\
        );

    \I__2776\ : LocalMux
    port map (
            O => \N__25064\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9\
        );

    \I__2775\ : InMux
    port map (
            O => \N__25059\,
            I => \N__25056\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__25056\,
            I => \N__25053\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__25053\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_6
        );

    \I__2772\ : CascadeMux
    port map (
            O => \N__25050\,
            I => \N__25047\
        );

    \I__2771\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25044\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__25044\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_6\
        );

    \I__2769\ : InMux
    port map (
            O => \N__25041\,
            I => \N__25038\
        );

    \I__2768\ : LocalMux
    port map (
            O => \N__25038\,
            I => \N__25035\
        );

    \I__2767\ : Odrv4
    port map (
            O => \N__25035\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_7
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__25032\,
            I => \N__25029\
        );

    \I__2765\ : InMux
    port map (
            O => \N__25029\,
            I => \N__25026\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__25026\,
            I => \N__25023\
        );

    \I__2763\ : Span4Mux_h
    port map (
            O => \N__25023\,
            I => \N__25020\
        );

    \I__2762\ : Span4Mux_h
    port map (
            O => \N__25020\,
            I => \N__25017\
        );

    \I__2761\ : Odrv4
    port map (
            O => \N__25017\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_7\
        );

    \I__2760\ : InMux
    port map (
            O => \N__25014\,
            I => \N__25011\
        );

    \I__2759\ : LocalMux
    port map (
            O => \N__25011\,
            I => \N__25008\
        );

    \I__2758\ : Odrv4
    port map (
            O => \N__25008\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_7\
        );

    \I__2757\ : CascadeMux
    port map (
            O => \N__25005\,
            I => \N__25001\
        );

    \I__2756\ : CascadeMux
    port map (
            O => \N__25004\,
            I => \N__24998\
        );

    \I__2755\ : CascadeBuf
    port map (
            O => \N__25001\,
            I => \N__24995\
        );

    \I__2754\ : CascadeBuf
    port map (
            O => \N__24998\,
            I => \N__24992\
        );

    \I__2753\ : CascadeMux
    port map (
            O => \N__24995\,
            I => \N__24989\
        );

    \I__2752\ : CascadeMux
    port map (
            O => \N__24992\,
            I => \N__24986\
        );

    \I__2751\ : CascadeBuf
    port map (
            O => \N__24989\,
            I => \N__24983\
        );

    \I__2750\ : CascadeBuf
    port map (
            O => \N__24986\,
            I => \N__24980\
        );

    \I__2749\ : CascadeMux
    port map (
            O => \N__24983\,
            I => \N__24977\
        );

    \I__2748\ : CascadeMux
    port map (
            O => \N__24980\,
            I => \N__24974\
        );

    \I__2747\ : CascadeBuf
    port map (
            O => \N__24977\,
            I => \N__24971\
        );

    \I__2746\ : CascadeBuf
    port map (
            O => \N__24974\,
            I => \N__24968\
        );

    \I__2745\ : CascadeMux
    port map (
            O => \N__24971\,
            I => \N__24965\
        );

    \I__2744\ : CascadeMux
    port map (
            O => \N__24968\,
            I => \N__24962\
        );

    \I__2743\ : CascadeBuf
    port map (
            O => \N__24965\,
            I => \N__24959\
        );

    \I__2742\ : CascadeBuf
    port map (
            O => \N__24962\,
            I => \N__24956\
        );

    \I__2741\ : CascadeMux
    port map (
            O => \N__24959\,
            I => \N__24953\
        );

    \I__2740\ : CascadeMux
    port map (
            O => \N__24956\,
            I => \N__24950\
        );

    \I__2739\ : CascadeBuf
    port map (
            O => \N__24953\,
            I => \N__24947\
        );

    \I__2738\ : CascadeBuf
    port map (
            O => \N__24950\,
            I => \N__24944\
        );

    \I__2737\ : CascadeMux
    port map (
            O => \N__24947\,
            I => \N__24941\
        );

    \I__2736\ : CascadeMux
    port map (
            O => \N__24944\,
            I => \N__24938\
        );

    \I__2735\ : CascadeBuf
    port map (
            O => \N__24941\,
            I => \N__24935\
        );

    \I__2734\ : CascadeBuf
    port map (
            O => \N__24938\,
            I => \N__24932\
        );

    \I__2733\ : CascadeMux
    port map (
            O => \N__24935\,
            I => \N__24929\
        );

    \I__2732\ : CascadeMux
    port map (
            O => \N__24932\,
            I => \N__24926\
        );

    \I__2731\ : CascadeBuf
    port map (
            O => \N__24929\,
            I => \N__24923\
        );

    \I__2730\ : CascadeBuf
    port map (
            O => \N__24926\,
            I => \N__24920\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__24923\,
            I => \N__24917\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__24920\,
            I => \N__24914\
        );

    \I__2727\ : InMux
    port map (
            O => \N__24917\,
            I => \N__24911\
        );

    \I__2726\ : InMux
    port map (
            O => \N__24914\,
            I => \N__24908\
        );

    \I__2725\ : LocalMux
    port map (
            O => \N__24911\,
            I => \N__24905\
        );

    \I__2724\ : LocalMux
    port map (
            O => \N__24908\,
            I => \N__24902\
        );

    \I__2723\ : Span4Mux_h
    port map (
            O => \N__24905\,
            I => \N__24899\
        );

    \I__2722\ : Span4Mux_h
    port map (
            O => \N__24902\,
            I => \N__24896\
        );

    \I__2721\ : Odrv4
    port map (
            O => \N__24899\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4\
        );

    \I__2720\ : Odrv4
    port map (
            O => \N__24896\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4\
        );

    \I__2719\ : CEMux
    port map (
            O => \N__24891\,
            I => \N__24888\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__24888\,
            I => \N__24884\
        );

    \I__2717\ : CEMux
    port map (
            O => \N__24887\,
            I => \N__24881\
        );

    \I__2716\ : Span4Mux_h
    port map (
            O => \N__24884\,
            I => \N__24876\
        );

    \I__2715\ : LocalMux
    port map (
            O => \N__24881\,
            I => \N__24876\
        );

    \I__2714\ : Odrv4
    port map (
            O => \N__24876\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1827_0\
        );

    \I__2713\ : CascadeMux
    port map (
            O => \N__24873\,
            I => \N__24870\
        );

    \I__2712\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24867\
        );

    \I__2711\ : LocalMux
    port map (
            O => \N__24867\,
            I => \N__24864\
        );

    \I__2710\ : Span4Mux_h
    port map (
            O => \N__24864\,
            I => \N__24861\
        );

    \I__2709\ : Span4Mux_v
    port map (
            O => \N__24861\,
            I => \N__24858\
        );

    \I__2708\ : Odrv4
    port map (
            O => \N__24858\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_7
        );

    \I__2707\ : CascadeMux
    port map (
            O => \N__24855\,
            I => \N__24852\
        );

    \I__2706\ : InMux
    port map (
            O => \N__24852\,
            I => \N__24849\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__24849\,
            I => \N__24846\
        );

    \I__2704\ : Span4Mux_h
    port map (
            O => \N__24846\,
            I => \N__24843\
        );

    \I__2703\ : Odrv4
    port map (
            O => \N__24843\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.N_863\
        );

    \I__2702\ : IoInMux
    port map (
            O => \N__24840\,
            I => \N__24837\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__24837\,
            I => \N__24833\
        );

    \I__2700\ : IoInMux
    port map (
            O => \N__24836\,
            I => \N__24830\
        );

    \I__2699\ : IoSpan4Mux
    port map (
            O => \N__24833\,
            I => \N__24825\
        );

    \I__2698\ : LocalMux
    port map (
            O => \N__24830\,
            I => \N__24825\
        );

    \I__2697\ : IoSpan4Mux
    port map (
            O => \N__24825\,
            I => \N__24822\
        );

    \I__2696\ : Span4Mux_s3_h
    port map (
            O => \N__24822\,
            I => \N__24819\
        );

    \I__2695\ : Span4Mux_h
    port map (
            O => \N__24819\,
            I => \N__24815\
        );

    \I__2694\ : InMux
    port map (
            O => \N__24818\,
            I => \N__24812\
        );

    \I__2693\ : Odrv4
    port map (
            O => \N__24815\,
            I => s1_c
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__24812\,
            I => s1_c
        );

    \I__2691\ : CascadeMux
    port map (
            O => \N__24807\,
            I => \N__24804\
        );

    \I__2690\ : CascadeBuf
    port map (
            O => \N__24804\,
            I => \N__24800\
        );

    \I__2689\ : CascadeMux
    port map (
            O => \N__24803\,
            I => \N__24797\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__24800\,
            I => \N__24794\
        );

    \I__2687\ : CascadeBuf
    port map (
            O => \N__24797\,
            I => \N__24791\
        );

    \I__2686\ : CascadeBuf
    port map (
            O => \N__24794\,
            I => \N__24788\
        );

    \I__2685\ : CascadeMux
    port map (
            O => \N__24791\,
            I => \N__24785\
        );

    \I__2684\ : CascadeMux
    port map (
            O => \N__24788\,
            I => \N__24782\
        );

    \I__2683\ : CascadeBuf
    port map (
            O => \N__24785\,
            I => \N__24779\
        );

    \I__2682\ : CascadeBuf
    port map (
            O => \N__24782\,
            I => \N__24776\
        );

    \I__2681\ : CascadeMux
    port map (
            O => \N__24779\,
            I => \N__24773\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__24776\,
            I => \N__24770\
        );

    \I__2679\ : CascadeBuf
    port map (
            O => \N__24773\,
            I => \N__24767\
        );

    \I__2678\ : CascadeBuf
    port map (
            O => \N__24770\,
            I => \N__24764\
        );

    \I__2677\ : CascadeMux
    port map (
            O => \N__24767\,
            I => \N__24761\
        );

    \I__2676\ : CascadeMux
    port map (
            O => \N__24764\,
            I => \N__24758\
        );

    \I__2675\ : CascadeBuf
    port map (
            O => \N__24761\,
            I => \N__24755\
        );

    \I__2674\ : CascadeBuf
    port map (
            O => \N__24758\,
            I => \N__24752\
        );

    \I__2673\ : CascadeMux
    port map (
            O => \N__24755\,
            I => \N__24749\
        );

    \I__2672\ : CascadeMux
    port map (
            O => \N__24752\,
            I => \N__24746\
        );

    \I__2671\ : CascadeBuf
    port map (
            O => \N__24749\,
            I => \N__24743\
        );

    \I__2670\ : CascadeBuf
    port map (
            O => \N__24746\,
            I => \N__24740\
        );

    \I__2669\ : CascadeMux
    port map (
            O => \N__24743\,
            I => \N__24737\
        );

    \I__2668\ : CascadeMux
    port map (
            O => \N__24740\,
            I => \N__24734\
        );

    \I__2667\ : CascadeBuf
    port map (
            O => \N__24737\,
            I => \N__24731\
        );

    \I__2666\ : CascadeBuf
    port map (
            O => \N__24734\,
            I => \N__24728\
        );

    \I__2665\ : CascadeMux
    port map (
            O => \N__24731\,
            I => \N__24725\
        );

    \I__2664\ : CascadeMux
    port map (
            O => \N__24728\,
            I => \N__24722\
        );

    \I__2663\ : CascadeBuf
    port map (
            O => \N__24725\,
            I => \N__24719\
        );

    \I__2662\ : InMux
    port map (
            O => \N__24722\,
            I => \N__24716\
        );

    \I__2661\ : CascadeMux
    port map (
            O => \N__24719\,
            I => \N__24713\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__24716\,
            I => \N__24710\
        );

    \I__2659\ : InMux
    port map (
            O => \N__24713\,
            I => \N__24707\
        );

    \I__2658\ : Odrv4
    port map (
            O => \N__24710\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5\
        );

    \I__2657\ : LocalMux
    port map (
            O => \N__24707\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5\
        );

    \I__2656\ : InMux
    port map (
            O => \N__24702\,
            I => \N__24699\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__24699\,
            I => \N__24694\
        );

    \I__2654\ : InMux
    port map (
            O => \N__24698\,
            I => \N__24691\
        );

    \I__2653\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24688\
        );

    \I__2652\ : Span4Mux_s3_v
    port map (
            O => \N__24694\,
            I => \N__24683\
        );

    \I__2651\ : LocalMux
    port map (
            O => \N__24691\,
            I => \N__24683\
        );

    \I__2650\ : LocalMux
    port map (
            O => \N__24688\,
            I => \N__24680\
        );

    \I__2649\ : Span4Mux_v
    port map (
            O => \N__24683\,
            I => \N__24674\
        );

    \I__2648\ : Span4Mux_v
    port map (
            O => \N__24680\,
            I => \N__24674\
        );

    \I__2647\ : InMux
    port map (
            O => \N__24679\,
            I => \N__24671\
        );

    \I__2646\ : Odrv4
    port map (
            O => \N__24674\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__24671\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0\
        );

    \I__2644\ : InMux
    port map (
            O => \N__24666\,
            I => \N__24662\
        );

    \I__2643\ : InMux
    port map (
            O => \N__24665\,
            I => \N__24658\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__24662\,
            I => \N__24654\
        );

    \I__2641\ : InMux
    port map (
            O => \N__24661\,
            I => \N__24651\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__24658\,
            I => \N__24648\
        );

    \I__2639\ : InMux
    port map (
            O => \N__24657\,
            I => \N__24645\
        );

    \I__2638\ : Span4Mux_h
    port map (
            O => \N__24654\,
            I => \N__24642\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__24651\,
            I => \N__24639\
        );

    \I__2636\ : Span4Mux_v
    port map (
            O => \N__24648\,
            I => \N__24634\
        );

    \I__2635\ : LocalMux
    port map (
            O => \N__24645\,
            I => \N__24634\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__24642\,
            I => \N__24629\
        );

    \I__2633\ : Span4Mux_h
    port map (
            O => \N__24639\,
            I => \N__24629\
        );

    \I__2632\ : Odrv4
    port map (
            O => \N__24634\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0\
        );

    \I__2631\ : Odrv4
    port map (
            O => \N__24629\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0\
        );

    \I__2630\ : InMux
    port map (
            O => \N__24624\,
            I => \N__24621\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__24621\,
            I => \N__24616\
        );

    \I__2628\ : InMux
    port map (
            O => \N__24620\,
            I => \N__24613\
        );

    \I__2627\ : InMux
    port map (
            O => \N__24619\,
            I => \N__24610\
        );

    \I__2626\ : Span4Mux_s3_v
    port map (
            O => \N__24616\,
            I => \N__24605\
        );

    \I__2625\ : LocalMux
    port map (
            O => \N__24613\,
            I => \N__24605\
        );

    \I__2624\ : LocalMux
    port map (
            O => \N__24610\,
            I => \N__24602\
        );

    \I__2623\ : Span4Mux_v
    port map (
            O => \N__24605\,
            I => \N__24596\
        );

    \I__2622\ : Span4Mux_v
    port map (
            O => \N__24602\,
            I => \N__24596\
        );

    \I__2621\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24593\
        );

    \I__2620\ : Odrv4
    port map (
            O => \N__24596\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__24593\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0\
        );

    \I__2618\ : InMux
    port map (
            O => \N__24588\,
            I => \N__24585\
        );

    \I__2617\ : LocalMux
    port map (
            O => \N__24585\,
            I => \N__24580\
        );

    \I__2616\ : InMux
    port map (
            O => \N__24584\,
            I => \N__24577\
        );

    \I__2615\ : InMux
    port map (
            O => \N__24583\,
            I => \N__24574\
        );

    \I__2614\ : Span4Mux_s2_v
    port map (
            O => \N__24580\,
            I => \N__24571\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__24577\,
            I => \N__24568\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__24574\,
            I => \N__24565\
        );

    \I__2611\ : Span4Mux_v
    port map (
            O => \N__24571\,
            I => \N__24557\
        );

    \I__2610\ : Span4Mux_v
    port map (
            O => \N__24568\,
            I => \N__24557\
        );

    \I__2609\ : Span4Mux_h
    port map (
            O => \N__24565\,
            I => \N__24557\
        );

    \I__2608\ : InMux
    port map (
            O => \N__24564\,
            I => \N__24554\
        );

    \I__2607\ : Odrv4
    port map (
            O => \N__24557\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__24554\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0\
        );

    \I__2605\ : CEMux
    port map (
            O => \N__24549\,
            I => \N__24545\
        );

    \I__2604\ : CEMux
    port map (
            O => \N__24548\,
            I => \N__24542\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__24545\,
            I => \N__24537\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__24542\,
            I => \N__24537\
        );

    \I__2601\ : Odrv4
    port map (
            O => \N__24537\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1826_0\
        );

    \I__2600\ : InMux
    port map (
            O => \N__24534\,
            I => \N__24529\
        );

    \I__2599\ : InMux
    port map (
            O => \N__24533\,
            I => \N__24526\
        );

    \I__2598\ : InMux
    port map (
            O => \N__24532\,
            I => \N__24523\
        );

    \I__2597\ : LocalMux
    port map (
            O => \N__24529\,
            I => \N__24520\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__24526\,
            I => \N__24517\
        );

    \I__2595\ : LocalMux
    port map (
            O => \N__24523\,
            I => \N__24514\
        );

    \I__2594\ : Span4Mux_v
    port map (
            O => \N__24520\,
            I => \N__24510\
        );

    \I__2593\ : Span4Mux_v
    port map (
            O => \N__24517\,
            I => \N__24505\
        );

    \I__2592\ : Span4Mux_h
    port map (
            O => \N__24514\,
            I => \N__24505\
        );

    \I__2591\ : InMux
    port map (
            O => \N__24513\,
            I => \N__24502\
        );

    \I__2590\ : Odrv4
    port map (
            O => \N__24510\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0\
        );

    \I__2589\ : Odrv4
    port map (
            O => \N__24505\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0\
        );

    \I__2588\ : LocalMux
    port map (
            O => \N__24502\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0\
        );

    \I__2587\ : InMux
    port map (
            O => \N__24495\,
            I => \N__24492\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__24492\,
            I => \N__24488\
        );

    \I__2585\ : InMux
    port map (
            O => \N__24491\,
            I => \N__24485\
        );

    \I__2584\ : Span4Mux_s2_v
    port map (
            O => \N__24488\,
            I => \N__24478\
        );

    \I__2583\ : LocalMux
    port map (
            O => \N__24485\,
            I => \N__24478\
        );

    \I__2582\ : InMux
    port map (
            O => \N__24484\,
            I => \N__24475\
        );

    \I__2581\ : InMux
    port map (
            O => \N__24483\,
            I => \N__24472\
        );

    \I__2580\ : Span4Mux_v
    port map (
            O => \N__24478\,
            I => \N__24467\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__24475\,
            I => \N__24467\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__24472\,
            I => \N__24464\
        );

    \I__2577\ : Odrv4
    port map (
            O => \N__24467\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0\
        );

    \I__2576\ : Odrv4
    port map (
            O => \N__24464\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0\
        );

    \I__2575\ : InMux
    port map (
            O => \N__24459\,
            I => \N__24456\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__24456\,
            I => \N__24453\
        );

    \I__2573\ : Span4Mux_s2_v
    port map (
            O => \N__24453\,
            I => \N__24449\
        );

    \I__2572\ : InMux
    port map (
            O => \N__24452\,
            I => \N__24446\
        );

    \I__2571\ : Span4Mux_v
    port map (
            O => \N__24449\,
            I => \N__24440\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__24446\,
            I => \N__24440\
        );

    \I__2569\ : InMux
    port map (
            O => \N__24445\,
            I => \N__24437\
        );

    \I__2568\ : Span4Mux_h
    port map (
            O => \N__24440\,
            I => \N__24434\
        );

    \I__2567\ : LocalMux
    port map (
            O => \N__24437\,
            I => \N__24431\
        );

    \I__2566\ : Span4Mux_v
    port map (
            O => \N__24434\,
            I => \N__24425\
        );

    \I__2565\ : Span4Mux_v
    port map (
            O => \N__24431\,
            I => \N__24425\
        );

    \I__2564\ : InMux
    port map (
            O => \N__24430\,
            I => \N__24422\
        );

    \I__2563\ : Odrv4
    port map (
            O => \N__24425\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0\
        );

    \I__2562\ : LocalMux
    port map (
            O => \N__24422\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0\
        );

    \I__2561\ : InMux
    port map (
            O => \N__24417\,
            I => \N__24414\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__24414\,
            I => \N__24411\
        );

    \I__2559\ : Odrv4
    port map (
            O => \N__24411\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_1_5
        );

    \I__2558\ : CascadeMux
    port map (
            O => \N__24408\,
            I => \N__24405\
        );

    \I__2557\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24402\
        );

    \I__2556\ : LocalMux
    port map (
            O => \N__24402\,
            I => \N__24399\
        );

    \I__2555\ : Span4Mux_h
    port map (
            O => \N__24399\,
            I => \N__24396\
        );

    \I__2554\ : Odrv4
    port map (
            O => \N__24396\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_5\
        );

    \I__2553\ : InMux
    port map (
            O => \N__24393\,
            I => \N__24388\
        );

    \I__2552\ : InMux
    port map (
            O => \N__24392\,
            I => \N__24384\
        );

    \I__2551\ : InMux
    port map (
            O => \N__24391\,
            I => \N__24381\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__24388\,
            I => \N__24378\
        );

    \I__2549\ : InMux
    port map (
            O => \N__24387\,
            I => \N__24375\
        );

    \I__2548\ : LocalMux
    port map (
            O => \N__24384\,
            I => \N__24372\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__24381\,
            I => \N__24369\
        );

    \I__2546\ : Span4Mux_s3_v
    port map (
            O => \N__24378\,
            I => \N__24364\
        );

    \I__2545\ : LocalMux
    port map (
            O => \N__24375\,
            I => \N__24364\
        );

    \I__2544\ : Span4Mux_v
    port map (
            O => \N__24372\,
            I => \N__24359\
        );

    \I__2543\ : Span4Mux_h
    port map (
            O => \N__24369\,
            I => \N__24359\
        );

    \I__2542\ : Odrv4
    port map (
            O => \N__24364\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__24359\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0\
        );

    \I__2540\ : InMux
    port map (
            O => \N__24354\,
            I => \N__24350\
        );

    \I__2539\ : InMux
    port map (
            O => \N__24353\,
            I => \N__24346\
        );

    \I__2538\ : LocalMux
    port map (
            O => \N__24350\,
            I => \N__24342\
        );

    \I__2537\ : InMux
    port map (
            O => \N__24349\,
            I => \N__24339\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__24346\,
            I => \N__24336\
        );

    \I__2535\ : InMux
    port map (
            O => \N__24345\,
            I => \N__24333\
        );

    \I__2534\ : Span4Mux_s3_v
    port map (
            O => \N__24342\,
            I => \N__24328\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__24339\,
            I => \N__24328\
        );

    \I__2532\ : Span4Mux_v
    port map (
            O => \N__24336\,
            I => \N__24323\
        );

    \I__2531\ : LocalMux
    port map (
            O => \N__24333\,
            I => \N__24323\
        );

    \I__2530\ : Odrv4
    port map (
            O => \N__24328\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0\
        );

    \I__2529\ : Odrv4
    port map (
            O => \N__24323\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0\
        );

    \I__2528\ : InMux
    port map (
            O => \N__24318\,
            I => \N__24314\
        );

    \I__2527\ : InMux
    port map (
            O => \N__24317\,
            I => \N__24311\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__24314\,
            I => \N__24307\
        );

    \I__2525\ : LocalMux
    port map (
            O => \N__24311\,
            I => \N__24304\
        );

    \I__2524\ : InMux
    port map (
            O => \N__24310\,
            I => \N__24301\
        );

    \I__2523\ : Span4Mux_h
    port map (
            O => \N__24307\,
            I => \N__24298\
        );

    \I__2522\ : Span4Mux_v
    port map (
            O => \N__24304\,
            I => \N__24293\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__24301\,
            I => \N__24293\
        );

    \I__2520\ : Span4Mux_v
    port map (
            O => \N__24298\,
            I => \N__24287\
        );

    \I__2519\ : Span4Mux_v
    port map (
            O => \N__24293\,
            I => \N__24287\
        );

    \I__2518\ : InMux
    port map (
            O => \N__24292\,
            I => \N__24284\
        );

    \I__2517\ : Odrv4
    port map (
            O => \N__24287\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0\
        );

    \I__2516\ : LocalMux
    port map (
            O => \N__24284\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0\
        );

    \I__2515\ : InMux
    port map (
            O => \N__24279\,
            I => \N__24276\
        );

    \I__2514\ : LocalMux
    port map (
            O => \N__24276\,
            I => \N__24271\
        );

    \I__2513\ : InMux
    port map (
            O => \N__24275\,
            I => \N__24268\
        );

    \I__2512\ : InMux
    port map (
            O => \N__24274\,
            I => \N__24265\
        );

    \I__2511\ : Span4Mux_s0_v
    port map (
            O => \N__24271\,
            I => \N__24262\
        );

    \I__2510\ : LocalMux
    port map (
            O => \N__24268\,
            I => \N__24259\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__24265\,
            I => \N__24256\
        );

    \I__2508\ : Span4Mux_v
    port map (
            O => \N__24262\,
            I => \N__24248\
        );

    \I__2507\ : Span4Mux_v
    port map (
            O => \N__24259\,
            I => \N__24248\
        );

    \I__2506\ : Span4Mux_h
    port map (
            O => \N__24256\,
            I => \N__24248\
        );

    \I__2505\ : InMux
    port map (
            O => \N__24255\,
            I => \N__24245\
        );

    \I__2504\ : Odrv4
    port map (
            O => \N__24248\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__24245\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0\
        );

    \I__2502\ : InMux
    port map (
            O => \N__24240\,
            I => \N__24236\
        );

    \I__2501\ : InMux
    port map (
            O => \N__24239\,
            I => \N__24232\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__24236\,
            I => \N__24228\
        );

    \I__2499\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24225\
        );

    \I__2498\ : LocalMux
    port map (
            O => \N__24232\,
            I => \N__24222\
        );

    \I__2497\ : InMux
    port map (
            O => \N__24231\,
            I => \N__24219\
        );

    \I__2496\ : Span4Mux_h
    port map (
            O => \N__24228\,
            I => \N__24216\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__24225\,
            I => \N__24213\
        );

    \I__2494\ : Span4Mux_v
    port map (
            O => \N__24222\,
            I => \N__24208\
        );

    \I__2493\ : LocalMux
    port map (
            O => \N__24219\,
            I => \N__24208\
        );

    \I__2492\ : Span4Mux_v
    port map (
            O => \N__24216\,
            I => \N__24203\
        );

    \I__2491\ : Span4Mux_h
    port map (
            O => \N__24213\,
            I => \N__24203\
        );

    \I__2490\ : Odrv4
    port map (
            O => \N__24208\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0\
        );

    \I__2489\ : Odrv4
    port map (
            O => \N__24203\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0\
        );

    \I__2488\ : InMux
    port map (
            O => \N__24198\,
            I => \N__24194\
        );

    \I__2487\ : InMux
    port map (
            O => \N__24197\,
            I => \N__24190\
        );

    \I__2486\ : LocalMux
    port map (
            O => \N__24194\,
            I => \N__24186\
        );

    \I__2485\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24183\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__24190\,
            I => \N__24180\
        );

    \I__2483\ : InMux
    port map (
            O => \N__24189\,
            I => \N__24177\
        );

    \I__2482\ : Span4Mux_v
    port map (
            O => \N__24186\,
            I => \N__24172\
        );

    \I__2481\ : LocalMux
    port map (
            O => \N__24183\,
            I => \N__24172\
        );

    \I__2480\ : Span4Mux_v
    port map (
            O => \N__24180\,
            I => \N__24167\
        );

    \I__2479\ : LocalMux
    port map (
            O => \N__24177\,
            I => \N__24167\
        );

    \I__2478\ : Span4Mux_v
    port map (
            O => \N__24172\,
            I => \N__24164\
        );

    \I__2477\ : Odrv4
    port map (
            O => \N__24167\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0\
        );

    \I__2476\ : Odrv4
    port map (
            O => \N__24164\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0\
        );

    \I__2475\ : InMux
    port map (
            O => \N__24159\,
            I => \N__24155\
        );

    \I__2474\ : InMux
    port map (
            O => \N__24158\,
            I => \N__24151\
        );

    \I__2473\ : LocalMux
    port map (
            O => \N__24155\,
            I => \N__24147\
        );

    \I__2472\ : InMux
    port map (
            O => \N__24154\,
            I => \N__24144\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__24151\,
            I => \N__24141\
        );

    \I__2470\ : InMux
    port map (
            O => \N__24150\,
            I => \N__24138\
        );

    \I__2469\ : Span4Mux_v
    port map (
            O => \N__24147\,
            I => \N__24133\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__24144\,
            I => \N__24133\
        );

    \I__2467\ : Span4Mux_v
    port map (
            O => \N__24141\,
            I => \N__24128\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__24138\,
            I => \N__24128\
        );

    \I__2465\ : Span4Mux_v
    port map (
            O => \N__24133\,
            I => \N__24123\
        );

    \I__2464\ : Span4Mux_v
    port map (
            O => \N__24128\,
            I => \N__24123\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__24123\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_448_0\
        );

    \I__2462\ : InMux
    port map (
            O => \N__24120\,
            I => \N__24114\
        );

    \I__2461\ : InMux
    port map (
            O => \N__24119\,
            I => \N__24111\
        );

    \I__2460\ : InMux
    port map (
            O => \N__24118\,
            I => \N__24108\
        );

    \I__2459\ : InMux
    port map (
            O => \N__24117\,
            I => \N__24105\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__24114\,
            I => \N__24102\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__24111\,
            I => \N__24099\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__24108\,
            I => \N__24096\
        );

    \I__2455\ : LocalMux
    port map (
            O => \N__24105\,
            I => \N__24093\
        );

    \I__2454\ : Span4Mux_v
    port map (
            O => \N__24102\,
            I => \N__24090\
        );

    \I__2453\ : Span4Mux_v
    port map (
            O => \N__24099\,
            I => \N__24083\
        );

    \I__2452\ : Span4Mux_h
    port map (
            O => \N__24096\,
            I => \N__24083\
        );

    \I__2451\ : Span4Mux_h
    port map (
            O => \N__24093\,
            I => \N__24083\
        );

    \I__2450\ : Odrv4
    port map (
            O => \N__24090\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0\
        );

    \I__2449\ : Odrv4
    port map (
            O => \N__24083\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0\
        );

    \I__2448\ : InMux
    port map (
            O => \N__24078\,
            I => \N__24074\
        );

    \I__2447\ : InMux
    port map (
            O => \N__24077\,
            I => \N__24070\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__24074\,
            I => \N__24066\
        );

    \I__2445\ : InMux
    port map (
            O => \N__24073\,
            I => \N__24063\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__24070\,
            I => \N__24060\
        );

    \I__2443\ : InMux
    port map (
            O => \N__24069\,
            I => \N__24057\
        );

    \I__2442\ : Span4Mux_v
    port map (
            O => \N__24066\,
            I => \N__24052\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__24063\,
            I => \N__24052\
        );

    \I__2440\ : Span4Mux_v
    port map (
            O => \N__24060\,
            I => \N__24047\
        );

    \I__2439\ : LocalMux
    port map (
            O => \N__24057\,
            I => \N__24047\
        );

    \I__2438\ : Odrv4
    port map (
            O => \N__24052\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0\
        );

    \I__2437\ : Odrv4
    port map (
            O => \N__24047\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0\
        );

    \I__2436\ : InMux
    port map (
            O => \N__24042\,
            I => \N__24038\
        );

    \I__2435\ : InMux
    port map (
            O => \N__24041\,
            I => \N__24034\
        );

    \I__2434\ : LocalMux
    port map (
            O => \N__24038\,
            I => \N__24030\
        );

    \I__2433\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24027\
        );

    \I__2432\ : LocalMux
    port map (
            O => \N__24034\,
            I => \N__24024\
        );

    \I__2431\ : InMux
    port map (
            O => \N__24033\,
            I => \N__24021\
        );

    \I__2430\ : Span4Mux_v
    port map (
            O => \N__24030\,
            I => \N__24016\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__24027\,
            I => \N__24016\
        );

    \I__2428\ : Span4Mux_s2_v
    port map (
            O => \N__24024\,
            I => \N__24011\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__24021\,
            I => \N__24011\
        );

    \I__2426\ : Odrv4
    port map (
            O => \N__24016\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0\
        );

    \I__2425\ : Odrv4
    port map (
            O => \N__24011\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0\
        );

    \I__2424\ : InMux
    port map (
            O => \N__24006\,
            I => \N__24002\
        );

    \I__2423\ : InMux
    port map (
            O => \N__24005\,
            I => \N__23999\
        );

    \I__2422\ : LocalMux
    port map (
            O => \N__24002\,
            I => \N__23995\
        );

    \I__2421\ : LocalMux
    port map (
            O => \N__23999\,
            I => \N__23992\
        );

    \I__2420\ : InMux
    port map (
            O => \N__23998\,
            I => \N__23988\
        );

    \I__2419\ : Span4Mux_s0_v
    port map (
            O => \N__23995\,
            I => \N__23985\
        );

    \I__2418\ : Span4Mux_h
    port map (
            O => \N__23992\,
            I => \N__23982\
        );

    \I__2417\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23979\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__23988\,
            I => \N__23976\
        );

    \I__2415\ : Span4Mux_v
    port map (
            O => \N__23985\,
            I => \N__23967\
        );

    \I__2414\ : Span4Mux_v
    port map (
            O => \N__23982\,
            I => \N__23967\
        );

    \I__2413\ : LocalMux
    port map (
            O => \N__23979\,
            I => \N__23967\
        );

    \I__2412\ : Span4Mux_h
    port map (
            O => \N__23976\,
            I => \N__23967\
        );

    \I__2411\ : Odrv4
    port map (
            O => \N__23967\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_459_0\
        );

    \I__2410\ : InMux
    port map (
            O => \N__23964\,
            I => \N__23958\
        );

    \I__2409\ : InMux
    port map (
            O => \N__23963\,
            I => \N__23955\
        );

    \I__2408\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23952\
        );

    \I__2407\ : InMux
    port map (
            O => \N__23961\,
            I => \N__23949\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__23958\,
            I => \N__23946\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__23955\,
            I => \N__23943\
        );

    \I__2404\ : LocalMux
    port map (
            O => \N__23952\,
            I => \N__23940\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__23949\,
            I => \N__23937\
        );

    \I__2402\ : Span4Mux_s2_v
    port map (
            O => \N__23946\,
            I => \N__23934\
        );

    \I__2401\ : Span4Mux_v
    port map (
            O => \N__23943\,
            I => \N__23927\
        );

    \I__2400\ : Span4Mux_h
    port map (
            O => \N__23940\,
            I => \N__23927\
        );

    \I__2399\ : Span4Mux_h
    port map (
            O => \N__23937\,
            I => \N__23927\
        );

    \I__2398\ : Odrv4
    port map (
            O => \N__23934\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0\
        );

    \I__2397\ : Odrv4
    port map (
            O => \N__23927\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0\
        );

    \I__2396\ : InMux
    port map (
            O => \N__23922\,
            I => \N__23917\
        );

    \I__2395\ : InMux
    port map (
            O => \N__23921\,
            I => \N__23914\
        );

    \I__2394\ : InMux
    port map (
            O => \N__23920\,
            I => \N__23910\
        );

    \I__2393\ : LocalMux
    port map (
            O => \N__23917\,
            I => \N__23907\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__23914\,
            I => \N__23904\
        );

    \I__2391\ : InMux
    port map (
            O => \N__23913\,
            I => \N__23901\
        );

    \I__2390\ : LocalMux
    port map (
            O => \N__23910\,
            I => \N__23898\
        );

    \I__2389\ : Span4Mux_s3_v
    port map (
            O => \N__23907\,
            I => \N__23895\
        );

    \I__2388\ : Span4Mux_v
    port map (
            O => \N__23904\,
            I => \N__23888\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__23901\,
            I => \N__23888\
        );

    \I__2386\ : Span4Mux_h
    port map (
            O => \N__23898\,
            I => \N__23888\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__23895\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0\
        );

    \I__2384\ : Odrv4
    port map (
            O => \N__23888\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0\
        );

    \I__2383\ : InMux
    port map (
            O => \N__23883\,
            I => \N__23879\
        );

    \I__2382\ : InMux
    port map (
            O => \N__23882\,
            I => \N__23875\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__23879\,
            I => \N__23872\
        );

    \I__2380\ : InMux
    port map (
            O => \N__23878\,
            I => \N__23869\
        );

    \I__2379\ : LocalMux
    port map (
            O => \N__23875\,
            I => \N__23866\
        );

    \I__2378\ : Span4Mux_v
    port map (
            O => \N__23872\,
            I => \N__23861\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__23869\,
            I => \N__23861\
        );

    \I__2376\ : Span4Mux_v
    port map (
            O => \N__23866\,
            I => \N__23855\
        );

    \I__2375\ : Span4Mux_v
    port map (
            O => \N__23861\,
            I => \N__23855\
        );

    \I__2374\ : InMux
    port map (
            O => \N__23860\,
            I => \N__23852\
        );

    \I__2373\ : Odrv4
    port map (
            O => \N__23855\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0\
        );

    \I__2372\ : LocalMux
    port map (
            O => \N__23852\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0\
        );

    \I__2371\ : InMux
    port map (
            O => \N__23847\,
            I => \N__23844\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__23844\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_1_8
        );

    \I__2369\ : InMux
    port map (
            O => \N__23841\,
            I => \N__23837\
        );

    \I__2368\ : InMux
    port map (
            O => \N__23840\,
            I => \N__23833\
        );

    \I__2367\ : LocalMux
    port map (
            O => \N__23837\,
            I => \N__23830\
        );

    \I__2366\ : InMux
    port map (
            O => \N__23836\,
            I => \N__23827\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__23833\,
            I => \N__23824\
        );

    \I__2364\ : Span4Mux_v
    port map (
            O => \N__23830\,
            I => \N__23819\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__23827\,
            I => \N__23819\
        );

    \I__2362\ : Span4Mux_h
    port map (
            O => \N__23824\,
            I => \N__23815\
        );

    \I__2361\ : Span4Mux_v
    port map (
            O => \N__23819\,
            I => \N__23812\
        );

    \I__2360\ : InMux
    port map (
            O => \N__23818\,
            I => \N__23809\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__23815\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__23812\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__23809\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0\
        );

    \I__2356\ : CascadeMux
    port map (
            O => \N__23802\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0_cascade_\
        );

    \I__2355\ : InMux
    port map (
            O => \N__23799\,
            I => \N__23795\
        );

    \I__2354\ : InMux
    port map (
            O => \N__23798\,
            I => \N__23791\
        );

    \I__2353\ : LocalMux
    port map (
            O => \N__23795\,
            I => \N__23787\
        );

    \I__2352\ : InMux
    port map (
            O => \N__23794\,
            I => \N__23784\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__23791\,
            I => \N__23781\
        );

    \I__2350\ : InMux
    port map (
            O => \N__23790\,
            I => \N__23778\
        );

    \I__2349\ : Span4Mux_s3_v
    port map (
            O => \N__23787\,
            I => \N__23773\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__23784\,
            I => \N__23773\
        );

    \I__2347\ : Span4Mux_v
    port map (
            O => \N__23781\,
            I => \N__23768\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__23778\,
            I => \N__23768\
        );

    \I__2345\ : Span4Mux_v
    port map (
            O => \N__23773\,
            I => \N__23763\
        );

    \I__2344\ : Span4Mux_v
    port map (
            O => \N__23768\,
            I => \N__23763\
        );

    \I__2343\ : Odrv4
    port map (
            O => \N__23763\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_466_0\
        );

    \I__2342\ : CascadeMux
    port map (
            O => \N__23760\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.csb_u_i_a2_0_0_cascade_\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__23757\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_331_cascade_\
        );

    \I__2340\ : CascadeMux
    port map (
            O => \N__23754\,
            I => \N__23751\
        );

    \I__2339\ : InMux
    port map (
            O => \N__23751\,
            I => \N__23748\
        );

    \I__2338\ : LocalMux
    port map (
            O => \N__23748\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_0\
        );

    \I__2337\ : InMux
    port map (
            O => \N__23745\,
            I => \N__23742\
        );

    \I__2336\ : LocalMux
    port map (
            O => \N__23742\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.m7_0_a2_3\
        );

    \I__2335\ : CEMux
    port map (
            O => \N__23739\,
            I => \N__23736\
        );

    \I__2334\ : LocalMux
    port map (
            O => \N__23736\,
            I => \N__23733\
        );

    \I__2333\ : Span4Mux_v
    port map (
            O => \N__23733\,
            I => \N__23729\
        );

    \I__2332\ : CEMux
    port map (
            O => \N__23732\,
            I => \N__23726\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__23729\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0\
        );

    \I__2330\ : LocalMux
    port map (
            O => \N__23726\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0\
        );

    \I__2329\ : InMux
    port map (
            O => \N__23721\,
            I => \N__23717\
        );

    \I__2328\ : InMux
    port map (
            O => \N__23720\,
            I => \N__23713\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__23717\,
            I => \N__23710\
        );

    \I__2326\ : InMux
    port map (
            O => \N__23716\,
            I => \N__23707\
        );

    \I__2325\ : LocalMux
    port map (
            O => \N__23713\,
            I => \N__23704\
        );

    \I__2324\ : Span4Mux_v
    port map (
            O => \N__23710\,
            I => \N__23699\
        );

    \I__2323\ : LocalMux
    port map (
            O => \N__23707\,
            I => \N__23699\
        );

    \I__2322\ : Span4Mux_v
    port map (
            O => \N__23704\,
            I => \N__23693\
        );

    \I__2321\ : Span4Mux_v
    port map (
            O => \N__23699\,
            I => \N__23693\
        );

    \I__2320\ : InMux
    port map (
            O => \N__23698\,
            I => \N__23690\
        );

    \I__2319\ : Odrv4
    port map (
            O => \N__23693\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__23690\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0\
        );

    \I__2317\ : InMux
    port map (
            O => \N__23685\,
            I => \N__23681\
        );

    \I__2316\ : InMux
    port map (
            O => \N__23684\,
            I => \N__23678\
        );

    \I__2315\ : LocalMux
    port map (
            O => \N__23681\,
            I => \N__23674\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__23678\,
            I => \N__23671\
        );

    \I__2313\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23668\
        );

    \I__2312\ : Span4Mux_s1_v
    port map (
            O => \N__23674\,
            I => \N__23665\
        );

    \I__2311\ : Span4Mux_v
    port map (
            O => \N__23671\,
            I => \N__23660\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__23668\,
            I => \N__23660\
        );

    \I__2309\ : Span4Mux_v
    port map (
            O => \N__23665\,
            I => \N__23654\
        );

    \I__2308\ : Span4Mux_v
    port map (
            O => \N__23660\,
            I => \N__23654\
        );

    \I__2307\ : InMux
    port map (
            O => \N__23659\,
            I => \N__23651\
        );

    \I__2306\ : Odrv4
    port map (
            O => \N__23654\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0\
        );

    \I__2305\ : LocalMux
    port map (
            O => \N__23651\,
            I => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0\
        );

    \I__2304\ : CascadeMux
    port map (
            O => \N__23646\,
            I => \N__23643\
        );

    \I__2303\ : InMux
    port map (
            O => \N__23643\,
            I => \N__23640\
        );

    \I__2302\ : LocalMux
    port map (
            O => \N__23640\,
            I => \N__23637\
        );

    \I__2301\ : Span4Mux_h
    port map (
            O => \N__23637\,
            I => \N__23634\
        );

    \I__2300\ : Span4Mux_v
    port map (
            O => \N__23634\,
            I => \N__23631\
        );

    \I__2299\ : Span4Mux_v
    port map (
            O => \N__23631\,
            I => \N__23628\
        );

    \I__2298\ : Odrv4
    port map (
            O => \N__23628\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_CO\
        );

    \I__2297\ : InMux
    port map (
            O => \N__23625\,
            I => \N__23622\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__23622\,
            I => \N__23618\
        );

    \I__2295\ : InMux
    port map (
            O => \N__23621\,
            I => \N__23615\
        );

    \I__2294\ : Span4Mux_v
    port map (
            O => \N__23618\,
            I => \N__23610\
        );

    \I__2293\ : LocalMux
    port map (
            O => \N__23615\,
            I => \N__23610\
        );

    \I__2292\ : Span4Mux_h
    port map (
            O => \N__23610\,
            I => \N__23607\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__23607\,
            I => \N__23603\
        );

    \I__2290\ : InMux
    port map (
            O => \N__23606\,
            I => \N__23600\
        );

    \I__2289\ : Span4Mux_v
    port map (
            O => \N__23603\,
            I => \N__23597\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__23600\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__23597\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2\
        );

    \I__2286\ : CascadeMux
    port map (
            O => \N__23592\,
            I => \N__23588\
        );

    \I__2285\ : InMux
    port map (
            O => \N__23591\,
            I => \N__23582\
        );

    \I__2284\ : InMux
    port map (
            O => \N__23588\,
            I => \N__23582\
        );

    \I__2283\ : InMux
    port map (
            O => \N__23587\,
            I => \N__23579\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__23582\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__23579\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15\
        );

    \I__2280\ : InMux
    port map (
            O => \N__23574\,
            I => \N__23568\
        );

    \I__2279\ : InMux
    port map (
            O => \N__23573\,
            I => \N__23568\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__23568\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_13\
        );

    \I__2277\ : InMux
    port map (
            O => \N__23565\,
            I => \N__23560\
        );

    \I__2276\ : InMux
    port map (
            O => \N__23564\,
            I => \N__23557\
        );

    \I__2275\ : InMux
    port map (
            O => \N__23563\,
            I => \N__23554\
        );

    \I__2274\ : LocalMux
    port map (
            O => \N__23560\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__23557\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2\
        );

    \I__2272\ : LocalMux
    port map (
            O => \N__23554\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2\
        );

    \I__2271\ : InMux
    port map (
            O => \N__23547\,
            I => \N__23542\
        );

    \I__2270\ : InMux
    port map (
            O => \N__23546\,
            I => \N__23539\
        );

    \I__2269\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23536\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__23542\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__23539\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__23536\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__23529\,
            I => \N__23524\
        );

    \I__2264\ : InMux
    port map (
            O => \N__23528\,
            I => \N__23521\
        );

    \I__2263\ : InMux
    port map (
            O => \N__23527\,
            I => \N__23518\
        );

    \I__2262\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23515\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__23521\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3\
        );

    \I__2260\ : LocalMux
    port map (
            O => \N__23518\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3\
        );

    \I__2259\ : LocalMux
    port map (
            O => \N__23515\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3\
        );

    \I__2258\ : InMux
    port map (
            O => \N__23508\,
            I => \N__23503\
        );

    \I__2257\ : InMux
    port map (
            O => \N__23507\,
            I => \N__23500\
        );

    \I__2256\ : InMux
    port map (
            O => \N__23506\,
            I => \N__23497\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__23503\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__23500\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__23497\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0\
        );

    \I__2252\ : CascadeMux
    port map (
            O => \N__23490\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383_cascade_\
        );

    \I__2251\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23480\
        );

    \I__2250\ : InMux
    port map (
            O => \N__23486\,
            I => \N__23480\
        );

    \I__2249\ : InMux
    port map (
            O => \N__23485\,
            I => \N__23477\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__23480\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__23477\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0\
        );

    \I__2246\ : CascadeMux
    port map (
            O => \N__23472\,
            I => \N__23468\
        );

    \I__2245\ : InMux
    port map (
            O => \N__23471\,
            I => \N__23463\
        );

    \I__2244\ : InMux
    port map (
            O => \N__23468\,
            I => \N__23463\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__23463\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_16\
        );

    \I__2242\ : CascadeMux
    port map (
            O => \N__23460\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_369_cascade_\
        );

    \I__2241\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23454\
        );

    \I__2240\ : LocalMux
    port map (
            O => \N__23454\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_12\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__23451\,
            I => \N__23443\
        );

    \I__2238\ : InMux
    port map (
            O => \N__23450\,
            I => \N__23438\
        );

    \I__2237\ : InMux
    port map (
            O => \N__23449\,
            I => \N__23433\
        );

    \I__2236\ : InMux
    port map (
            O => \N__23448\,
            I => \N__23433\
        );

    \I__2235\ : InMux
    port map (
            O => \N__23447\,
            I => \N__23428\
        );

    \I__2234\ : InMux
    port map (
            O => \N__23446\,
            I => \N__23428\
        );

    \I__2233\ : InMux
    port map (
            O => \N__23443\,
            I => \N__23425\
        );

    \I__2232\ : InMux
    port map (
            O => \N__23442\,
            I => \N__23422\
        );

    \I__2231\ : InMux
    port map (
            O => \N__23441\,
            I => \N__23419\
        );

    \I__2230\ : LocalMux
    port map (
            O => \N__23438\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__23433\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__23428\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__23425\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__23422\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__23419\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\
        );

    \I__2224\ : InMux
    port map (
            O => \N__23406\,
            I => \N__23395\
        );

    \I__2223\ : InMux
    port map (
            O => \N__23405\,
            I => \N__23395\
        );

    \I__2222\ : InMux
    port map (
            O => \N__23404\,
            I => \N__23395\
        );

    \I__2221\ : InMux
    port map (
            O => \N__23403\,
            I => \N__23390\
        );

    \I__2220\ : InMux
    port map (
            O => \N__23402\,
            I => \N__23390\
        );

    \I__2219\ : LocalMux
    port map (
            O => \N__23395\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__23390\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383\
        );

    \I__2217\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23378\
        );

    \I__2216\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23378\
        );

    \I__2215\ : InMux
    port map (
            O => \N__23383\,
            I => \N__23375\
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__23378\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__23375\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7\
        );

    \I__2212\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23367\
        );

    \I__2211\ : LocalMux
    port map (
            O => \N__23367\,
            I => \N__23363\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__23366\,
            I => \N__23360\
        );

    \I__2209\ : Span4Mux_h
    port map (
            O => \N__23363\,
            I => \N__23357\
        );

    \I__2208\ : InMux
    port map (
            O => \N__23360\,
            I => \N__23354\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__23357\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__23354\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16\
        );

    \I__2205\ : InMux
    port map (
            O => \N__23349\,
            I => \N__23344\
        );

    \I__2204\ : InMux
    port map (
            O => \N__23348\,
            I => \N__23341\
        );

    \I__2203\ : InMux
    port map (
            O => \N__23347\,
            I => \N__23338\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__23344\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__23341\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__23338\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__23331\,
            I => \N__23328\
        );

    \I__2198\ : InMux
    port map (
            O => \N__23328\,
            I => \N__23325\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__23325\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_0\
        );

    \I__2196\ : CascadeMux
    port map (
            O => \N__23322\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0_cascade_\
        );

    \I__2195\ : InMux
    port map (
            O => \N__23319\,
            I => \N__23316\
        );

    \I__2194\ : LocalMux
    port map (
            O => \N__23316\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_4\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__23313\,
            I => \N__23310\
        );

    \I__2192\ : InMux
    port map (
            O => \N__23310\,
            I => \N__23304\
        );

    \I__2191\ : InMux
    port map (
            O => \N__23309\,
            I => \N__23304\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__23304\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_5\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__23301\,
            I => \N__23298\
        );

    \I__2188\ : InMux
    port map (
            O => \N__23298\,
            I => \N__23292\
        );

    \I__2187\ : InMux
    port map (
            O => \N__23297\,
            I => \N__23292\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__23292\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_8\
        );

    \I__2185\ : InMux
    port map (
            O => \N__23289\,
            I => \N__23285\
        );

    \I__2184\ : InMux
    port map (
            O => \N__23288\,
            I => \N__23282\
        );

    \I__2183\ : LocalMux
    port map (
            O => \N__23285\,
            I => \N__23279\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__23282\,
            I => \N__23276\
        );

    \I__2181\ : Span4Mux_h
    port map (
            O => \N__23279\,
            I => \N__23273\
        );

    \I__2180\ : Odrv4
    port map (
            O => \N__23276\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15\
        );

    \I__2179\ : Odrv4
    port map (
            O => \N__23273\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15\
        );

    \I__2178\ : CascadeMux
    port map (
            O => \N__23268\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1Z0Z_23_cascade_\
        );

    \I__2177\ : IoInMux
    port map (
            O => \N__23265\,
            I => \N__23262\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__23262\,
            I => \N__23259\
        );

    \I__2175\ : IoSpan4Mux
    port map (
            O => \N__23259\,
            I => \N__23256\
        );

    \I__2174\ : Span4Mux_s0_v
    port map (
            O => \N__23256\,
            I => \N__23253\
        );

    \I__2173\ : Span4Mux_v
    port map (
            O => \N__23253\,
            I => \N__23250\
        );

    \I__2172\ : Sp12to4
    port map (
            O => \N__23250\,
            I => \N__23247\
        );

    \I__2171\ : Odrv12
    port map (
            O => \N__23247\,
            I => \N_29\
        );

    \I__2170\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23241\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__23241\,
            I => \N__23238\
        );

    \I__2168\ : Span4Mux_h
    port map (
            O => \N__23238\,
            I => \N__23235\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__23235\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_read\
        );

    \I__2166\ : InMux
    port map (
            O => \N__23232\,
            I => \N__23229\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__23229\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01Z0Z_0\
        );

    \I__2164\ : InMux
    port map (
            O => \N__23226\,
            I => \N__23223\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__23223\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_reti_0_1\
        );

    \I__2162\ : InMux
    port map (
            O => \N__23220\,
            I => \N__23217\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__23217\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0\
        );

    \I__2160\ : CascadeMux
    port map (
            O => \N__23214\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0_cascade_\
        );

    \I__2159\ : InMux
    port map (
            O => \N__23211\,
            I => \N__23208\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__23208\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.sclk_u_i_0\
        );

    \I__2157\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23202\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__23202\,
            I => \N__23199\
        );

    \I__2155\ : Sp12to4
    port map (
            O => \N__23199\,
            I => \N__23196\
        );

    \I__2154\ : Span12Mux_v
    port map (
            O => \N__23196\,
            I => \N__23193\
        );

    \I__2153\ : Odrv12
    port map (
            O => \N__23193\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_1_7
        );

    \I__2152\ : CascadeMux
    port map (
            O => \N__23190\,
            I => \N__23187\
        );

    \I__2151\ : InMux
    port map (
            O => \N__23187\,
            I => \N__23184\
        );

    \I__2150\ : LocalMux
    port map (
            O => \N__23184\,
            I => \N__23181\
        );

    \I__2149\ : Span4Mux_h
    port map (
            O => \N__23181\,
            I => \N__23178\
        );

    \I__2148\ : Span4Mux_v
    port map (
            O => \N__23178\,
            I => \N__23175\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__23175\,
            I => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_1_7
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__23172\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_7_cascade_\
        );

    \I__2145\ : InMux
    port map (
            O => \N__23169\,
            I => \N__23166\
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__23166\,
            I => \N__23163\
        );

    \I__2143\ : Span4Mux_h
    port map (
            O => \N__23163\,
            I => \N__23160\
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__23160\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_7\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__23157\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_7_cascade_\
        );

    \I__2140\ : InMux
    port map (
            O => \N__23154\,
            I => \N__23151\
        );

    \I__2139\ : LocalMux
    port map (
            O => \N__23151\,
            I => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_7\
        );

    \I__2138\ : InMux
    port map (
            O => \N__23148\,
            I => \N__23145\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__23145\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.dout_read\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__23142\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_237_cascade_\
        );

    \I__2135\ : IoInMux
    port map (
            O => \N__23139\,
            I => \N__23136\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__23136\,
            I => \N__23133\
        );

    \I__2133\ : Span4Mux_s2_h
    port map (
            O => \N__23133\,
            I => \N__23130\
        );

    \I__2132\ : Span4Mux_v
    port map (
            O => \N__23130\,
            I => \N__23127\
        );

    \I__2131\ : Odrv4
    port map (
            O => \N__23127\,
            I => \N_85_0\
        );

    \I__2130\ : InMux
    port map (
            O => \N__23124\,
            I => \N__23121\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__23121\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_6\
        );

    \I__2128\ : InMux
    port map (
            O => \N__23118\,
            I => \N__23115\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__23115\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_5\
        );

    \I__2126\ : InMux
    port map (
            O => \N__23112\,
            I => \N__23109\
        );

    \I__2125\ : LocalMux
    port map (
            O => \N__23109\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_4\
        );

    \I__2124\ : InMux
    port map (
            O => \N__23106\,
            I => \N__23103\
        );

    \I__2123\ : LocalMux
    port map (
            O => \N__23103\,
            I => \N__23100\
        );

    \I__2122\ : Span4Mux_v
    port map (
            O => \N__23100\,
            I => \N__23097\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__23097\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_2\
        );

    \I__2120\ : InMux
    port map (
            O => \N__23094\,
            I => \N__23091\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__23091\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_3\
        );

    \I__2118\ : CEMux
    port map (
            O => \N__23088\,
            I => \N__23084\
        );

    \I__2117\ : CEMux
    port map (
            O => \N__23087\,
            I => \N__23081\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__23084\,
            I => \N__23078\
        );

    \I__2115\ : LocalMux
    port map (
            O => \N__23081\,
            I => \N__23075\
        );

    \I__2114\ : Span4Mux_v
    port map (
            O => \N__23078\,
            I => \N__23070\
        );

    \I__2113\ : Span4Mux_h
    port map (
            O => \N__23075\,
            I => \N__23070\
        );

    \I__2112\ : Span4Mux_s3_h
    port map (
            O => \N__23070\,
            I => \N__23067\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__23067\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_370_i\
        );

    \I__2110\ : IoInMux
    port map (
            O => \N__23064\,
            I => \N__23061\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__23061\,
            I => \N__23058\
        );

    \I__2108\ : IoSpan4Mux
    port map (
            O => \N__23058\,
            I => \N__23055\
        );

    \I__2107\ : Span4Mux_s2_v
    port map (
            O => \N__23055\,
            I => \N__23052\
        );

    \I__2106\ : Sp12to4
    port map (
            O => \N__23052\,
            I => \N__23049\
        );

    \I__2105\ : Odrv12
    port map (
            O => \N__23049\,
            I => \N_1820_0\
        );

    \I__2104\ : InMux
    port map (
            O => \N__23046\,
            I => \N__23043\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__23043\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_u_i_0\
        );

    \I__2102\ : InMux
    port map (
            O => \N__23040\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2\
        );

    \I__2101\ : InMux
    port map (
            O => \N__23037\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_3\
        );

    \I__2100\ : CascadeMux
    port map (
            O => \N__23034\,
            I => \N__23031\
        );

    \I__2099\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23028\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__23028\,
            I => \N__23025\
        );

    \I__2097\ : Odrv4
    port map (
            O => \N__23025\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_333\
        );

    \I__2096\ : InMux
    port map (
            O => \N__23022\,
            I => \N__23019\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__23019\,
            I => \N__23016\
        );

    \I__2094\ : Span4Mux_h
    port map (
            O => \N__23016\,
            I => \N__23012\
        );

    \I__2093\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23009\
        );

    \I__2092\ : Sp12to4
    port map (
            O => \N__23012\,
            I => \N__23004\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__23009\,
            I => \N__23004\
        );

    \I__2090\ : Odrv12
    port map (
            O => \N__23004\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_376\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__23001\,
            I => \N__22998\
        );

    \I__2088\ : InMux
    port map (
            O => \N__22998\,
            I => \N__22995\
        );

    \I__2087\ : LocalMux
    port map (
            O => \N__22995\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1\
        );

    \I__2086\ : CascadeMux
    port map (
            O => \N__22992\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1_cascade_\
        );

    \I__2085\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22978\
        );

    \I__2084\ : InMux
    port map (
            O => \N__22988\,
            I => \N__22978\
        );

    \I__2083\ : InMux
    port map (
            O => \N__22987\,
            I => \N__22978\
        );

    \I__2082\ : InMux
    port map (
            O => \N__22986\,
            I => \N__22973\
        );

    \I__2081\ : InMux
    port map (
            O => \N__22985\,
            I => \N__22973\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__22978\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__22973\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0\
        );

    \I__2078\ : InMux
    port map (
            O => \N__22968\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0\
        );

    \I__2077\ : InMux
    port map (
            O => \N__22965\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1\
        );

    \I__2076\ : InMux
    port map (
            O => \N__22962\,
            I => \N__22958\
        );

    \I__2075\ : InMux
    port map (
            O => \N__22961\,
            I => \N__22954\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__22958\,
            I => \N__22951\
        );

    \I__2073\ : InMux
    port map (
            O => \N__22957\,
            I => \N__22948\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__22954\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3\
        );

    \I__2071\ : Odrv4
    port map (
            O => \N__22951\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__22948\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3\
        );

    \I__2069\ : CascadeMux
    port map (
            O => \N__22941\,
            I => \N__22938\
        );

    \I__2068\ : InMux
    port map (
            O => \N__22938\,
            I => \N__22935\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__22935\,
            I => \N__22932\
        );

    \I__2066\ : Odrv4
    port map (
            O => \N__22932\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_CO\
        );

    \I__2065\ : InMux
    port map (
            O => \N__22929\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2\
        );

    \I__2064\ : InMux
    port map (
            O => \N__22926\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_3\
        );

    \I__2063\ : InMux
    port map (
            O => \N__22923\,
            I => \N__22919\
        );

    \I__2062\ : InMux
    port map (
            O => \N__22922\,
            I => \N__22916\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__22919\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__22916\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4\
        );

    \I__2059\ : InMux
    port map (
            O => \N__22911\,
            I => \bfn_6_19_0_\
        );

    \I__2058\ : InMux
    port map (
            O => \N__22908\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0\
        );

    \I__2057\ : InMux
    port map (
            O => \N__22905\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1\
        );

    \I__2056\ : CascadeMux
    port map (
            O => \N__22902\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93Z0Z_0_cascade_\
        );

    \I__2055\ : IoInMux
    port map (
            O => \N__22899\,
            I => \N__22896\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__22896\,
            I => \N__22893\
        );

    \I__2053\ : Odrv12
    port map (
            O => \N__22893\,
            I => sclk1_c
        );

    \I__2052\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22887\
        );

    \I__2051\ : LocalMux
    port map (
            O => \N__22887\,
            I => \N__22884\
        );

    \I__2050\ : Span4Mux_v
    port map (
            O => \N__22884\,
            I => \N__22879\
        );

    \I__2049\ : InMux
    port map (
            O => \N__22883\,
            I => \N__22876\
        );

    \I__2048\ : InMux
    port map (
            O => \N__22882\,
            I => \N__22873\
        );

    \I__2047\ : Odrv4
    port map (
            O => \N__22879\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__22876\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__22873\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458\
        );

    \I__2044\ : InMux
    port map (
            O => \N__22866\,
            I => \N__22863\
        );

    \I__2043\ : LocalMux
    port map (
            O => \N__22863\,
            I => \N__22860\
        );

    \I__2042\ : Span4Mux_v
    port map (
            O => \N__22860\,
            I => \N__22852\
        );

    \I__2041\ : InMux
    port map (
            O => \N__22859\,
            I => \N__22847\
        );

    \I__2040\ : InMux
    port map (
            O => \N__22858\,
            I => \N__22847\
        );

    \I__2039\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22840\
        );

    \I__2038\ : InMux
    port map (
            O => \N__22856\,
            I => \N__22840\
        );

    \I__2037\ : InMux
    port map (
            O => \N__22855\,
            I => \N__22840\
        );

    \I__2036\ : Odrv4
    port map (
            O => \N__22852\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i\
        );

    \I__2035\ : LocalMux
    port map (
            O => \N__22847\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i\
        );

    \I__2034\ : LocalMux
    port map (
            O => \N__22840\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i\
        );

    \I__2033\ : InMux
    port map (
            O => \N__22833\,
            I => \N__22830\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__22830\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32Z0Z_0\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__22827\,
            I => \N__22822\
        );

    \I__2030\ : InMux
    port map (
            O => \N__22826\,
            I => \N__22819\
        );

    \I__2029\ : InMux
    port map (
            O => \N__22825\,
            I => \N__22816\
        );

    \I__2028\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22813\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__22819\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__22816\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__22813\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3\
        );

    \I__2024\ : InMux
    port map (
            O => \N__22806\,
            I => \N__22801\
        );

    \I__2023\ : InMux
    port map (
            O => \N__22805\,
            I => \N__22798\
        );

    \I__2022\ : InMux
    port map (
            O => \N__22804\,
            I => \N__22795\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__22801\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__22798\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2\
        );

    \I__2019\ : LocalMux
    port map (
            O => \N__22795\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2\
        );

    \I__2018\ : InMux
    port map (
            O => \N__22788\,
            I => \N__22783\
        );

    \I__2017\ : InMux
    port map (
            O => \N__22787\,
            I => \N__22780\
        );

    \I__2016\ : InMux
    port map (
            O => \N__22786\,
            I => \N__22777\
        );

    \I__2015\ : LocalMux
    port map (
            O => \N__22783\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1\
        );

    \I__2014\ : LocalMux
    port map (
            O => \N__22780\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__22777\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1\
        );

    \I__2012\ : InMux
    port map (
            O => \N__22770\,
            I => \N__22767\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__22767\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.un2_count_bits_1_0_a2_2\
        );

    \I__2010\ : CascadeMux
    port map (
            O => \N__22764\,
            I => \N__22759\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__22763\,
            I => \N__22756\
        );

    \I__2008\ : CascadeMux
    port map (
            O => \N__22762\,
            I => \N__22752\
        );

    \I__2007\ : InMux
    port map (
            O => \N__22759\,
            I => \N__22746\
        );

    \I__2006\ : InMux
    port map (
            O => \N__22756\,
            I => \N__22746\
        );

    \I__2005\ : InMux
    port map (
            O => \N__22755\,
            I => \N__22740\
        );

    \I__2004\ : InMux
    port map (
            O => \N__22752\,
            I => \N__22737\
        );

    \I__2003\ : InMux
    port map (
            O => \N__22751\,
            I => \N__22734\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__22746\,
            I => \N__22731\
        );

    \I__2001\ : InMux
    port map (
            O => \N__22745\,
            I => \N__22724\
        );

    \I__2000\ : InMux
    port map (
            O => \N__22744\,
            I => \N__22724\
        );

    \I__1999\ : InMux
    port map (
            O => \N__22743\,
            I => \N__22724\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__22740\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__22737\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__22734\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__22731\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\
        );

    \I__1994\ : LocalMux
    port map (
            O => \N__22724\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\
        );

    \I__1993\ : InMux
    port map (
            O => \N__22713\,
            I => \N__22707\
        );

    \I__1992\ : InMux
    port map (
            O => \N__22712\,
            I => \N__22707\
        );

    \I__1991\ : LocalMux
    port map (
            O => \N__22707\,
            I => \N__22700\
        );

    \I__1990\ : InMux
    port map (
            O => \N__22706\,
            I => \N__22697\
        );

    \I__1989\ : InMux
    port map (
            O => \N__22705\,
            I => \N__22690\
        );

    \I__1988\ : InMux
    port map (
            O => \N__22704\,
            I => \N__22690\
        );

    \I__1987\ : InMux
    port map (
            O => \N__22703\,
            I => \N__22690\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__22700\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__22697\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__22690\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383\
        );

    \I__1983\ : InMux
    port map (
            O => \N__22683\,
            I => \N__22678\
        );

    \I__1982\ : InMux
    port map (
            O => \N__22682\,
            I => \N__22673\
        );

    \I__1981\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22673\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__22678\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__22673\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6\
        );

    \I__1978\ : CascadeMux
    port map (
            O => \N__22668\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0_cascade_\
        );

    \I__1977\ : InMux
    port map (
            O => \N__22665\,
            I => \N__22662\
        );

    \I__1976\ : LocalMux
    port map (
            O => \N__22662\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_4\
        );

    \I__1975\ : InMux
    port map (
            O => \N__22659\,
            I => \N__22653\
        );

    \I__1974\ : InMux
    port map (
            O => \N__22658\,
            I => \N__22653\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__22653\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_5\
        );

    \I__1972\ : InMux
    port map (
            O => \N__22650\,
            I => \N__22646\
        );

    \I__1971\ : InMux
    port map (
            O => \N__22649\,
            I => \N__22643\
        );

    \I__1970\ : LocalMux
    port map (
            O => \N__22646\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__22643\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7\
        );

    \I__1968\ : InMux
    port map (
            O => \N__22638\,
            I => \N__22632\
        );

    \I__1967\ : InMux
    port map (
            O => \N__22637\,
            I => \N__22632\
        );

    \I__1966\ : LocalMux
    port map (
            O => \N__22632\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_8\
        );

    \I__1965\ : InMux
    port map (
            O => \N__22629\,
            I => \N__22626\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__22626\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_4\
        );

    \I__1963\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22620\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__22620\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_5\
        );

    \I__1961\ : InMux
    port map (
            O => \N__22617\,
            I => \N__22614\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__22614\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_6\
        );

    \I__1959\ : InMux
    port map (
            O => \N__22611\,
            I => \N__22608\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__22608\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_0\
        );

    \I__1957\ : CEMux
    port map (
            O => \N__22605\,
            I => \N__22602\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__22602\,
            I => \N__22599\
        );

    \I__1955\ : Span4Mux_v
    port map (
            O => \N__22599\,
            I => \N__22596\
        );

    \I__1954\ : Odrv4
    port map (
            O => \N__22596\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_i\
        );

    \I__1953\ : IoInMux
    port map (
            O => \N__22593\,
            I => \N__22590\
        );

    \I__1952\ : LocalMux
    port map (
            O => \N__22590\,
            I => \N__22587\
        );

    \I__1951\ : Span4Mux_s2_v
    port map (
            O => \N__22587\,
            I => \N__22584\
        );

    \I__1950\ : Span4Mux_v
    port map (
            O => \N__22584\,
            I => \N__22581\
        );

    \I__1949\ : Span4Mux_v
    port map (
            O => \N__22581\,
            I => \N__22578\
        );

    \I__1948\ : Odrv4
    port map (
            O => \N__22578\,
            I => \N_1821_0\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__22575\,
            I => \N__22572\
        );

    \I__1946\ : InMux
    port map (
            O => \N__22572\,
            I => \N__22569\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__22569\,
            I => \N__22566\
        );

    \I__1944\ : Span12Mux_s8_h
    port map (
            O => \N__22566\,
            I => \N__22563\
        );

    \I__1943\ : Span12Mux_v
    port map (
            O => \N__22563\,
            I => \N__22560\
        );

    \I__1942\ : Span12Mux_h
    port map (
            O => \N__22560\,
            I => \N__22557\
        );

    \I__1941\ : Odrv12
    port map (
            O => \N__22557\,
            I => sdin1_c
        );

    \I__1940\ : InMux
    port map (
            O => \N__22554\,
            I => \N__22551\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__22551\,
            I => \N__22548\
        );

    \I__1938\ : Span12Mux_h
    port map (
            O => \N__22548\,
            I => \N__22545\
        );

    \I__1937\ : Span12Mux_v
    port map (
            O => \N__22545\,
            I => \N__22542\
        );

    \I__1936\ : Span12Mux_h
    port map (
            O => \N__22542\,
            I => \N__22539\
        );

    \I__1935\ : Odrv12
    port map (
            O => \N__22539\,
            I => sdin0_c
        );

    \I__1934\ : IoInMux
    port map (
            O => \N__22536\,
            I => \N__22533\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__22533\,
            I => \N__22530\
        );

    \I__1932\ : Span4Mux_s1_h
    port map (
            O => \N__22530\,
            I => \N__22527\
        );

    \I__1931\ : Sp12to4
    port map (
            O => \N__22527\,
            I => \N__22524\
        );

    \I__1930\ : Span12Mux_v
    port map (
            O => \N__22524\,
            I => \N__22521\
        );

    \I__1929\ : Odrv12
    port map (
            O => \N__22521\,
            I => mcu_data_c
        );

    \I__1928\ : InMux
    port map (
            O => \N__22518\,
            I => \N__22513\
        );

    \I__1927\ : InMux
    port map (
            O => \N__22517\,
            I => \N__22510\
        );

    \I__1926\ : InMux
    port map (
            O => \N__22516\,
            I => \N__22507\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__22513\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__22510\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__22507\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0\
        );

    \I__1922\ : InMux
    port map (
            O => \N__22500\,
            I => \N__22496\
        );

    \I__1921\ : InMux
    port map (
            O => \N__22499\,
            I => \N__22493\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__22496\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0\
        );

    \I__1919\ : LocalMux
    port map (
            O => \N__22493\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0\
        );

    \I__1918\ : InMux
    port map (
            O => \N__22488\,
            I => \N__22482\
        );

    \I__1917\ : InMux
    port map (
            O => \N__22487\,
            I => \N__22482\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__22482\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370\
        );

    \I__1915\ : CascadeMux
    port map (
            O => \N__22479\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_cascade_\
        );

    \I__1914\ : InMux
    port map (
            O => \N__22476\,
            I => \N__22471\
        );

    \I__1913\ : InMux
    port map (
            O => \N__22475\,
            I => \N__22466\
        );

    \I__1912\ : InMux
    port map (
            O => \N__22474\,
            I => \N__22466\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__22471\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__22466\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14\
        );

    \I__1909\ : InMux
    port map (
            O => \N__22461\,
            I => \N__22458\
        );

    \I__1908\ : LocalMux
    port map (
            O => \N__22458\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_1\
        );

    \I__1907\ : InMux
    port map (
            O => \N__22455\,
            I => \N__22452\
        );

    \I__1906\ : LocalMux
    port map (
            O => \N__22452\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_2\
        );

    \I__1905\ : InMux
    port map (
            O => \N__22449\,
            I => \N__22446\
        );

    \I__1904\ : LocalMux
    port map (
            O => \N__22446\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_3\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__22443\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_17_0_cascade_\
        );

    \I__1902\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22437\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__22437\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_12\
        );

    \I__1900\ : CascadeMux
    port map (
            O => \N__22434\,
            I => \N__22430\
        );

    \I__1899\ : CascadeMux
    port map (
            O => \N__22433\,
            I => \N__22427\
        );

    \I__1898\ : InMux
    port map (
            O => \N__22430\,
            I => \N__22424\
        );

    \I__1897\ : InMux
    port map (
            O => \N__22427\,
            I => \N__22421\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__22424\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13\
        );

    \I__1895\ : LocalMux
    port map (
            O => \N__22421\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13\
        );

    \I__1894\ : InMux
    port map (
            O => \N__22416\,
            I => \N__22405\
        );

    \I__1893\ : InMux
    port map (
            O => \N__22415\,
            I => \N__22405\
        );

    \I__1892\ : InMux
    port map (
            O => \N__22414\,
            I => \N__22405\
        );

    \I__1891\ : InMux
    port map (
            O => \N__22413\,
            I => \N__22400\
        );

    \I__1890\ : InMux
    port map (
            O => \N__22412\,
            I => \N__22400\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__22405\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__22400\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0\
        );

    \I__1887\ : CascadeMux
    port map (
            O => \N__22395\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0_cascade_\
        );

    \I__1886\ : InMux
    port map (
            O => \N__22392\,
            I => \N__22389\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__22389\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_375\
        );

    \I__1884\ : InMux
    port map (
            O => \N__22386\,
            I => \N__22383\
        );

    \I__1883\ : LocalMux
    port map (
            O => \N__22383\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_1\
        );

    \I__1882\ : InMux
    port map (
            O => \N__22380\,
            I => \N__22377\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__22377\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_0\
        );

    \I__1880\ : InMux
    port map (
            O => \N__22374\,
            I => \bfn_5_16_0_\
        );

    \I__1879\ : InMux
    port map (
            O => \N__22371\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0\
        );

    \I__1878\ : InMux
    port map (
            O => \N__22368\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1\
        );

    \I__1877\ : InMux
    port map (
            O => \N__22365\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2\
        );

    \I__1876\ : InMux
    port map (
            O => \N__22362\,
            I => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_3\
        );

    \I__1875\ : IoInMux
    port map (
            O => \N__22359\,
            I => \N__22356\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__22356\,
            I => \N__22353\
        );

    \I__1873\ : Span4Mux_s3_h
    port map (
            O => \N__22353\,
            I => \N__22350\
        );

    \I__1872\ : Span4Mux_v
    port map (
            O => \N__22350\,
            I => \N__22347\
        );

    \I__1871\ : Odrv4
    port map (
            O => \N__22347\,
            I => mcu_sclk_c
        );

    \I__1870\ : IoInMux
    port map (
            O => \N__22344\,
            I => \N__22341\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__22341\,
            I => \N__22338\
        );

    \I__1868\ : Span12Mux_s5_v
    port map (
            O => \N__22338\,
            I => \N__22335\
        );

    \I__1867\ : Span12Mux_h
    port map (
            O => \N__22335\,
            I => \N__22332\
        );

    \I__1866\ : Span12Mux_v
    port map (
            O => \N__22332\,
            I => \N__22329\
        );

    \I__1865\ : Span12Mux_v
    port map (
            O => \N__22329\,
            I => \N__22326\
        );

    \I__1864\ : Odrv12
    port map (
            O => \N__22326\,
            I => clock_ibuf_gb_io_gb_input
        );

    \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            I => \N__47994\
        );

    \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            I => \N__47993\
        );

    \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            I => \N__47991\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net\,
            I => \N__65638\
        );

    \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\,
            I => \N__47985\
        );

    \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net\,
            I => \N__47979\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net\,
            I => \N__65637\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net\,
            I => \N__65612\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net\,
            I => \N__65592\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net\,
            I => \N__65650\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net\,
            I => \N__65636\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net\,
            I => \N__65624\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net\,
            I => \N__65603\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net\,
            I => \N__65635\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net\,
            I => \N__65590\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net\,
            I => \N__65579\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net\,
            I => \N__65621\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net\,
            I => \N__65600\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net\,
            I => \N__65578\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net\,
            I => \N__65543\
        );

    \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C_net\,
            I => \N__47981\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net\,
            I => \N__65542\
        );

    \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            I => \N__47982\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net\,
            I => \N__65563\
        );

    \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net\,
            I => \N__47989\
        );

    \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net\,
            I => \N__47987\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net\,
            I => \N__65526\
        );

    \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net\,
            I => \N__47988\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net\,
            I => \N__65607\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net\,
            I => \N__65540\
        );

    \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\,
            I => \N__47995\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net\,
            I => \N__65647\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            I => \N__65630\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net\,
            I => \N__65620\
        );

    \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net\,
            I => \N__47986\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net\,
            I => \N__65574\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net\,
            I => \N__65561\
        );

    \INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC\ : INV
    port map (
            O => \INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC_net\,
            I => \N__32744\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net\,
            I => \N__65671\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C_net\,
            I => \N__65656\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            I => \N__65646\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\,
            I => \N__65629\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net\,
            I => \N__65619\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net\,
            I => \N__65596\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\,
            I => \N__65645\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net\,
            I => \N__65628\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net\,
            I => \N__65655\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            I => \N__65644\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net\,
            I => \N__65627\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            I => \N__65713\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\,
            I => \N__65693\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            I => \N__65654\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            I => \N__65643\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\,
            I => \N__65617\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net\,
            I => \N__65735\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net\,
            I => \N__65752\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            I => \N__65743\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net\,
            I => \N__65734\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net\,
            I => \N__65723\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net\,
            I => \N__65705\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C_net\,
            I => \N__65664\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\,
            I => \N__65753\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net\,
            I => \N__65751\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\,
            I => \N__65722\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            I => \N__65750\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net\,
            I => \N__65741\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net\,
            I => \N__65732\
        );

    \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C\ : INV
    port map (
            O => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net\,
            I => \N__65749\
        );

    \IN_MUX_bfv_18_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_18_0_\
        );

    \IN_MUX_bfv_6_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_18_0_\
        );

    \IN_MUX_bfv_9_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_19_0_\
        );

    \IN_MUX_bfv_20_17_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_20_17_0_\
        );

    \IN_MUX_bfv_20_18_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7\,
            carryinitout => \bfn_20_18_0_\
        );

    \IN_MUX_bfv_21_27_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_21_27_0_\
        );

    \IN_MUX_bfv_5_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_16_0_\
        );

    \IN_MUX_bfv_11_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_15_0_\
        );

    \IN_MUX_bfv_11_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_19_0_\
        );

    \IN_MUX_bfv_6_19_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_19_0_\
        );

    \IN_MUX_bfv_9_22_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_22_0_\
        );

    \IN_MUX_bfv_12_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_12_20_0_\
        );

    \IN_MUX_bfv_18_20_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_18_20_0_\
        );

    \IN_MUX_bfv_18_21_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_7\,
            carryinitout => \bfn_18_21_0_\
        );

    \IN_MUX_bfv_13_23_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_13_23_0_\
        );

    \clock_ibuf_gb_io_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__22344\,
            GLOBALBUFFEROUTPUT => clock_c_g
        );

    \scl_ibuf_RNI7T7F\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__51207\,
            GLOBALBUFFEROUTPUT => scl_c_g
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_0_14\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__43296\,
            GLOBALBUFFEROUTPUT => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_g\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__32250\,
            GLOBALBUFFEROUTPUT => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_g\
        );

    \rst_n_ibuf_RNIBNDC_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34806\,
            GLOBALBUFFEROUTPUT => rst_n_c_i_g
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__34818\,
            GLOBALBUFFEROUTPUT => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_g\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__25422\,
            GLOBALBUFFEROUTPUT => \I2C_top_level_inst1.c_state4_0_i_g\
        );

    \IO_PIN_INST_RNIR662\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__57699\,
            GLOBALBUFFEROUTPUT => s_sda_i_g
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIK8VR2_15_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__23022\,
            in1 => \N__65767\,
            in2 => \_gnd_net_\,
            in3 => \N__22890\,
            lcout => mcu_sclk_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1_LC_4_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22380\,
            in2 => \_gnd_net_\,
            in3 => \N__30475\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net\,
            ce => \N__23088\,
            sr => \N__62944\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_2_LC_4_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30476\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22386\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net\,
            ce => \N__23088\,
            sr => \N__62944\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_0_LC_4_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30477\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_1C_net\,
            ce => \N__23088\,
            sr => \N__62944\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_0_LC_5_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22414\,
            in1 => \N__22518\,
            in2 => \_gnd_net_\,
            in3 => \N__22374\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_16_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0\,
            clk => \N__65721\,
            ce => 'H',
            sr => \N__62950\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_1_LC_5_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22412\,
            in1 => \N__22788\,
            in2 => \_gnd_net_\,
            in3 => \N__22371\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1\,
            clk => \N__65721\,
            ce => 'H',
            sr => \N__62950\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_2_LC_5_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22415\,
            in1 => \N__22806\,
            in2 => \_gnd_net_\,
            in3 => \N__22368\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_2\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2\,
            clk => \N__65721\,
            ce => 'H',
            sr => \N__62950\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_3_LC_5_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22413\,
            in1 => \N__22826\,
            in2 => \_gnd_net_\,
            in3 => \N__22365\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bitsZ0Z_3\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_cry_3\,
            clk => \N__65721\,
            ce => 'H',
            sr => \N__62950\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_4_LC_5_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22416\,
            in1 => \N__22755\,
            in2 => \_gnd_net_\,
            in3 => \N__22362\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_bits_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65721\,
            ce => 'H',
            sr => \N__62950\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_3_LC_5_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000010100"
        )
    port map (
            in0 => \N__25530\,
            in1 => \N__22961\,
            in2 => \N__22941\,
            in3 => \N__25583\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65721\,
            ce => 'H',
            sr => \N__62950\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13_LC_5_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22440\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net\,
            ce => 'H',
            sr => \N__62945\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m16_LC_5_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__22859\,
            in1 => \N__22703\,
            in2 => \_gnd_net_\,
            in3 => \N__22744\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_17_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_12_LC_5_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100011111010"
        )
    port map (
            in0 => \N__23370\,
            in1 => \N__25629\,
            in2 => \N__22443\,
            in3 => \N__23349\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net\,
            ce => 'H',
            sr => \N__62945\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_14_LC_5_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111001011111010"
        )
    port map (
            in0 => \N__22475\,
            in1 => \N__22704\,
            in2 => \N__22434\,
            in3 => \N__22745\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net\,
            ce => 'H',
            sr => \N__62945\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI5JQ51_13_LC_5_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__22658\,
            in1 => \N__22858\,
            in2 => \N__22433\,
            in3 => \N__22499\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_377_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_6_LC_5_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100101010"
        )
    port map (
            in0 => \N__22682\,
            in1 => \N__22705\,
            in2 => \N__22762\,
            in3 => \N__22659\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_13C_net\,
            ce => 'H',
            sr => \N__62945\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI1LAH_14_LC_5_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22474\,
            in2 => \_gnd_net_\,
            in3 => \N__22681\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_344_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNITF8T1_0_LC_5_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__22517\,
            in1 => \N__22770\,
            in2 => \N__22395\,
            in3 => \N__22743\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_375\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNILFTV2_9_LC_5_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__25075\,
            in1 => \N__22487\,
            in2 => \N__25696\,
            in3 => \N__22392\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_datae_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10_LC_5_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25076\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net\,
            ce => 'H',
            sr => \N__62939\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_11_LC_5_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__22713\,
            in1 => \N__22857\,
            in2 => \N__22763\,
            in3 => \N__22488\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_55_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net\,
            ce => 'H',
            sr => \N__62939\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_en_count_data_i_LC_5_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__22856\,
            in1 => \N__25686\,
            in2 => \N__25751\,
            in3 => \N__25074\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.en_count_data_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_11_LC_5_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25736\,
            in2 => \_gnd_net_\,
            in3 => \N__22855\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNI9LA6_0_11_LC_5_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22479\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.N_370_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_15_LC_5_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22712\,
            in1 => \_gnd_net_\,
            in2 => \N__22764\,
            in3 => \N__22476\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_10C_net\,
            ce => 'H',
            sr => \N__62939\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1_LC_5_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25740\,
            in2 => \_gnd_net_\,
            in3 => \N__22611\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_2_LC_5_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25741\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22461\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_3_LC_5_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25742\,
            in2 => \_gnd_net_\,
            in3 => \N__22455\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_4_LC_5_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__25743\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22449\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_5_LC_5_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25744\,
            in2 => \_gnd_net_\,
            in3 => \N__22629\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_6_LC_5_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__25745\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22623\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_7_LC_5_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25746\,
            in2 => \_gnd_net_\,
            in3 => \N__22617\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_read\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_0_LC_5_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__25747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.ser_data_1C_net\,
            ce => \N__22605\,
            sr => \N__62929\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNI8PPB5_0_LC_5_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__65769\,
            in1 => \N__23211\,
            in2 => \N__23034\,
            in3 => \N__27210\,
            lcout => \N_1821_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIBD7Q2_15_LC_6_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110001001000000"
        )
    port map (
            in0 => \N__22883\,
            in1 => \N__23015\,
            in2 => \N__22575\,
            in3 => \N__22554\,
            lcout => mcu_data_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNIEJ431_0_LC_6_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__22804\,
            in1 => \N__22786\,
            in2 => \N__22827\,
            in3 => \N__22516\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m33_e_LC_6_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__23288\,
            in1 => \N__22650\,
            in2 => \_gnd_net_\,
            in3 => \N__22500\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.N_1458\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93_0_LC_6_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011111110110101"
        )
    port map (
            in0 => \N__27568\,
            in1 => \N__27678\,
            in2 => \N__29970\,
            in3 => \N__28863\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIKUT93Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIA8O66_0_LC_6_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100001001100"
        )
    port map (
            in0 => \N__25695\,
            in1 => \N__65768\,
            in2 => \N__22902\,
            in3 => \N__22833\,
            lcout => sclk1_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32_0_LC_6_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111111011111"
        )
    port map (
            in0 => \N__27567\,
            in1 => \N__22882\,
            in2 => \N__29969\,
            in3 => \N__22866\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIJEL32Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_bits_RNI4GBQ_1_LC_6_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__22825\,
            in1 => \N__22805\,
            in2 => \_gnd_net_\,
            in3 => \N__22787\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.un2_count_bits_1_0_a2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7_LC_6_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__22751\,
            in1 => \N__22706\,
            in2 => \_gnd_net_\,
            in3 => \N__22683\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\,
            ce => 'H',
            sr => \N__62940\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_4_LC_6_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__22637\,
            in1 => \N__25627\,
            in2 => \_gnd_net_\,
            in3 => \N__23347\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\,
            ce => 'H',
            sr => \N__62940\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_RNIICQD1_4_LC_6_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__22957\,
            in1 => \N__23621\,
            in2 => \N__25491\,
            in3 => \N__22922\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_347_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_9_LC_6_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__22638\,
            in1 => \_gnd_net_\,
            in2 => \N__22668\,
            in3 => \N__25628\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\,
            ce => 'H',
            sr => \N__62940\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_5_LC_6_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22665\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\,
            ce => 'H',
            sr => \N__62940\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_8_LC_6_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22649\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_7C_net\,
            ce => 'H',
            sr => \N__62940\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_c_0_LC_6_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25617\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_18_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_6_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25487\,
            in2 => \_gnd_net_\,
            in3 => \N__22968\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_6_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23625\,
            in2 => \_gnd_net_\,
            in3 => \N__22965\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_6_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22962\,
            in2 => \_gnd_net_\,
            in3 => \N__22929\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_4_LC_6_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100110001100"
        )
    port map (
            in0 => \N__25577\,
            in1 => \N__22923\,
            in2 => \N__25535\,
            in3 => \N__22926\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65733\,
            ce => 'H',
            sr => \N__62930\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_0_LC_6_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22987\,
            in1 => \N__23508\,
            in2 => \_gnd_net_\,
            in3 => \N__22911\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_6_19_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0\,
            clk => \N__65742\,
            ce => 'H',
            sr => \N__62920\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_1_LC_6_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22985\,
            in1 => \N__23547\,
            in2 => \_gnd_net_\,
            in3 => \N__22908\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1\,
            clk => \N__65742\,
            ce => 'H',
            sr => \N__62920\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_2_LC_6_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22988\,
            in1 => \N__23565\,
            in2 => \_gnd_net_\,
            in3 => \N__22905\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_2\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2\,
            clk => \N__65742\,
            ce => 'H',
            sr => \N__62920\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_3_LC_6_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22986\,
            in1 => \N__23528\,
            in2 => \_gnd_net_\,
            in3 => \N__23040\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_3\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_cry_3\,
            clk => \N__65742\,
            ce => 'H',
            sr => \N__62920\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_4_LC_6_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__22989\,
            in1 => \N__23450\,
            in2 => \_gnd_net_\,
            in3 => \N__23037\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bitsZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65742\,
            ce => 'H',
            sr => \N__62920\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIMOE52_15_LC_6_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23385\,
            in1 => \N__23591\,
            in2 => \N__23001\,
            in3 => \N__26994\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_333\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI02AE1_15_LC_6_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25804\,
            in1 => \N__23384\,
            in2 => \N__23592\,
            in3 => \N__25839\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_376\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_sck_m8_i_a2_1_LC_6_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__25838\,
            in1 => \N__26923\,
            in2 => \_gnd_net_\,
            in3 => \N__25802\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI0EFP1_13_LC_6_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23573\,
            in2 => \N__22992\,
            in3 => \N__23309\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_377_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6_LC_6_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011111110000"
        )
    port map (
            in0 => \N__23405\,
            in1 => \N__23449\,
            in2 => \N__23313\,
            in3 => \N__25803\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net\,
            ce => 'H',
            sr => \N__62912\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_14_LC_6_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101110000"
        )
    port map (
            in0 => \N__23448\,
            in1 => \N__23404\,
            in2 => \N__25845\,
            in3 => \N__23574\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net\,
            ce => 'H',
            sr => \N__62912\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_11_LC_6_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111001100"
        )
    port map (
            in0 => \N__23406\,
            in1 => \N__30472\,
            in2 => \N__23451\,
            in3 => \N__26924\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_6C_net\,
            ce => 'H',
            sr => \N__62912\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7_LC_6_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23124\,
            in2 => \_gnd_net_\,
            in3 => \N__30463\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.dout_read\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\,
            ce => \N__23087\,
            sr => \N__62901\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_RNINM921_23_LC_6_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__32633\,
            in1 => \N__26124\,
            in2 => \_gnd_net_\,
            in3 => \N__49560\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_237_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_RNIU7DV3_7_LC_6_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010000000000"
        )
    port map (
            in0 => \N__26982\,
            in1 => \N__23148\,
            in2 => \N__23142\,
            in3 => \N__23046\,
            lcout => \N_85_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_6_LC_6_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__30462\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23118\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\,
            ce => \N__23087\,
            sr => \N__62901\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_5_LC_6_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23112\,
            in2 => \_gnd_net_\,
            in3 => \N__30461\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\,
            ce => \N__23087\,
            sr => \N__62901\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_4_LC_6_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30460\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23094\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\,
            ce => \N__23087\,
            sr => \N__62901\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI7VAM_11_LC_6_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30458\,
            in2 => \_gnd_net_\,
            in3 => \N__26932\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_370_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_3_LC_6_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30459\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23106\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.ser_data_7C_net\,
            ce => \N__23087\,
            sr => \N__62901\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNISO0C4_0_LC_6_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__25869\,
            in1 => \N__32635\,
            in2 => \N__23754\,
            in3 => \N__26997\,
            lcout => \N_1820_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIS2262_0_LC_6_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010001000100"
        )
    port map (
            in0 => \N__27195\,
            in1 => \N__23220\,
            in2 => \N__32640\,
            in3 => \N__26999\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_u_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIPJA61_0_LC_6_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010110100001010"
        )
    port map (
            in0 => \N__26998\,
            in1 => \N__27194\,
            in2 => \N__27150\,
            in3 => \N__32636\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_RNIPJA61_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNID2OK2_0_LC_6_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32634\,
            in2 => \N__23214\,
            in3 => \N__31098\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.sclk_u_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_7_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__53314\,
            in1 => \N__40529\,
            in2 => \N__38319\,
            in3 => \N__41058\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_7_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__52781\,
            in2 => \N__23190\,
            in3 => \N__52522\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_7_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52236\,
            in2 => \N__23172\,
            in3 => \N__40551\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_7_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__23169\,
            in1 => \N__33456\,
            in2 => \N__23157\,
            in3 => \N__23154\,
            lcout => \I2C_top_level_inst1_s_data_oreg_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65639\,
            ce => \N__54525\,
            sr => \N__64964\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_7_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51927\,
            in1 => \N__25014\,
            in2 => \N__24855\,
            in3 => \N__48759\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28999\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_4C_net\,
            ce => 'H',
            sr => \N__62951\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_5_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41806\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65679\,
            ce => \N__44092\,
            sr => \N__64963\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_7_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41689\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65679\,
            ce => \N__44092\,
            sr => \N__64963\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16_LC_7_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23289\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62931\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_LC_7_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23226\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62931\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18_LC_7_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29049\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net\,
            ce => 'H',
            sr => \N__62921\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1_23_LC_7_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011000000"
        )
    port map (
            in0 => \N__36129\,
            in1 => \N__26802\,
            in2 => \N__29968\,
            in3 => \N__27579\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNI7VVC1Z0Z_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_RNIUP1S2_23_LC_7_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__23232\,
            in1 => \_gnd_net_\,
            in2 => \N__23268\,
            in3 => \N__25682\,
            lcout => \N_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01_0_LC_7_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__29958\,
            in1 => \N__27578\,
            in2 => \_gnd_net_\,
            in3 => \N__23244\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNI4QS01Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHF2R_0_LC_7_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29957\,
            in2 => \_gnd_net_\,
            in3 => \N__35860\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_reti_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_1_LC_7_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35861\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37173\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1867_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_0_LC_7_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101110011001100"
        )
    port map (
            in0 => \N__25626\,
            in1 => \N__25681\,
            in2 => \N__23366\,
            in3 => \N__23348\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_18C_net\,
            ce => 'H',
            sr => \N__62921\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIN9BU_0_LC_7_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23442\,
            in1 => \N__23546\,
            in2 => \N__23331\,
            in3 => \N__23507\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNINH4C_2_LC_7_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23527\,
            in2 => \_gnd_net_\,
            in3 => \N__23564\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.un2_count_bits_1_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_RNIEOU21_4_LC_7_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__25926\,
            in1 => \N__25962\,
            in2 => \N__25887\,
            in3 => \N__25995\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_347_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4_LC_7_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23297\,
            in2 => \N__23322\,
            in3 => \N__25458\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net\,
            ce => 'H',
            sr => \N__62913\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_9_LC_7_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__25459\,
            in1 => \_gnd_net_\,
            in2 => \N__23301\,
            in3 => \N__23485\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net\,
            ce => 'H',
            sr => \N__62913\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_5_LC_7_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__23319\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net\,
            ce => 'H',
            sr => \N__62913\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_8_LC_7_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23383\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_4C_net\,
            ce => 'H',
            sr => \N__62913\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16_LC_7_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23587\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62902\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_15_LC_7_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23446\,
            in1 => \N__23402\,
            in2 => \_gnd_net_\,
            in3 => \N__25840\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62902\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_13_LC_7_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23457\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62902\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_0_LC_7_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101000000"
        )
    port map (
            in0 => \N__25460\,
            in1 => \N__23486\,
            in2 => \N__23472\,
            in3 => \N__26976\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62902\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_bits_RNIAV8O_0_LC_7_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__23563\,
            in1 => \N__23545\,
            in2 => \N__23529\,
            in3 => \N__23506\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_383_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNO_0_12_LC_7_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23441\,
            in2 => \N__23490\,
            in3 => \N__26931\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.N_369_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_12_LC_7_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011110100"
        )
    port map (
            in0 => \N__23487\,
            in1 => \N__23471\,
            in2 => \N__23460\,
            in3 => \N__25461\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62902\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_7_LC_7_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__23447\,
            in1 => \N__23403\,
            in2 => \_gnd_net_\,
            in3 => \N__25808\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_16C_net\,
            ce => 'H',
            sr => \N__62902\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0_LC_7_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__26013\,
            in1 => \N__26061\,
            in2 => \_gnd_net_\,
            in3 => \N__23745\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net\,
            ce => 'H',
            sr => \N__62889\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_1_LC_7_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27193\,
            in2 => \_gnd_net_\,
            in3 => \N__27107\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_0C_net\,
            ce => 'H',
            sr => \N__62889\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNI9R351_9_LC_7_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30514\,
            in1 => \N__32632\,
            in2 => \_gnd_net_\,
            in3 => \N__26996\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.csb_u_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNINIFT1_0_LC_7_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__30473\,
            in1 => \N__27183\,
            in2 => \N__23760\,
            in3 => \N__27069\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_331_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIG6Q33_0_LC_7_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__27035\,
            in1 => \N__32631\,
            in2 => \N__23757\,
            in3 => \N__26995\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_LC_7_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27182\,
            in2 => \_gnd_net_\,
            in3 => \N__27068\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_391_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_ns_1_0__m7_0_a2_3_LC_7_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__26079\,
            in1 => \N__26097\,
            in2 => \N__27036\,
            in3 => \N__26115\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.m7_0_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec0_0_a2_i_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__38919\,
            in1 => \N__38823\,
            in2 => \_gnd_net_\,
            in3 => \N__26673\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1828_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_0_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__61964\,
            in1 => \N__26336\,
            in2 => \_gnd_net_\,
            in3 => \N__50387\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_469_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_1_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__61820\,
            in1 => \N__26337\,
            in2 => \_gnd_net_\,
            in3 => \N__50388\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_468_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_2_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000010100"
        )
    port map (
            in0 => \N__25536\,
            in1 => \N__23606\,
            in2 => \N__23646\,
            in3 => \N__25590\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65555\,
            ce => 'H',
            sr => \N__62961\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_12_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__58561\,
            in1 => \N__26288\,
            in2 => \_gnd_net_\,
            in3 => \N__50405\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_460_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_13_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__50403\,
            in1 => \_gnd_net_\,
            in2 => \N__26330\,
            in3 => \N__58332\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_459_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_14_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__58455\,
            in1 => \N__26292\,
            in2 => \_gnd_net_\,
            in3 => \N__50406\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_458_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_15_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__50404\,
            in1 => \_gnd_net_\,
            in2 => \N__26331\,
            in3 => \N__57509\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_457_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_16_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__57636\,
            in1 => \N__26296\,
            in2 => \_gnd_net_\,
            in3 => \N__50402\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_456_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_8_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__61963\,
            in1 => \N__23847\,
            in2 => \N__44665\,
            in3 => \N__38372\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_20_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__61545\,
            in1 => \N__26264\,
            in2 => \_gnd_net_\,
            in3 => \N__50390\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_452_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_o3_0_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59554\,
            in2 => \_gnd_net_\,
            in3 => \N__50456\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_393_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_3_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63909\,
            in2 => \N__23802\,
            in3 => \N__50391\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_466_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_4_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__50393\,
            in1 => \_gnd_net_\,
            in2 => \N__26325\,
            in3 => \N__63799\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_465_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_5_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__63661\,
            in1 => \N__26271\,
            in2 => \_gnd_net_\,
            in3 => \N__50394\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_464_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_22_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__50389\,
            in1 => \_gnd_net_\,
            in2 => \N__26324\,
            in3 => \N__61310\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_450_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_9_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__46501\,
            in1 => \N__26263\,
            in2 => \_gnd_net_\,
            in3 => \N__50392\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1562_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_25_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50348\,
            in2 => \N__26326\,
            in3 => \N__61014\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1563_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_23_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__61246\,
            in1 => \N__26277\,
            in2 => \_gnd_net_\,
            in3 => \N__50352\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_449_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_26_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50347\,
            in2 => \N__26327\,
            in3 => \N__60912\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_448_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_21_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__50351\,
            in1 => \N__26276\,
            in2 => \_gnd_net_\,
            in3 => \N__61449\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_451_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_29_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50350\,
            in2 => \N__26328\,
            in3 => \N__62265\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_446_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_10_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__58749\,
            in1 => \N__26272\,
            in2 => \_gnd_net_\,
            in3 => \N__50353\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_284_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_30_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50349\,
            in2 => \N__26329\,
            in3 => \N__62132\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_445_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_2_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__61730\,
            in1 => \N__26284\,
            in2 => \_gnd_net_\,
            in3 => \N__50354\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_467_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_24_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__61126\,
            in1 => \N__50407\,
            in2 => \_gnd_net_\,
            in3 => \N__26332\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_286_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__38912\,
            in1 => \N__38806\,
            in2 => \_gnd_net_\,
            in3 => \N__26665\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1826_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_0_a2_i_27_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__60805\,
            in1 => \N__50408\,
            in2 => \_gnd_net_\,
            in3 => \N__26333\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1564_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_11_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__58666\,
            in1 => \N__26334\,
            in2 => \_gnd_net_\,
            in3 => \N__50380\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_461_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_28_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__62337\,
            in1 => \N__26335\,
            in2 => \_gnd_net_\,
            in3 => \N__50379\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_447_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_5_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__24417\,
            in1 => \N__44616\,
            in2 => \N__24408\,
            in3 => \N__44372\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_6_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__25059\,
            in1 => \N__44614\,
            in2 => \N__25050\,
            in3 => \N__44370\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_6_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41757\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65616\,
            ce => \N__44106\,
            sr => \N__64966\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_7_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__25041\,
            in1 => \N__44615\,
            in2 => \N__25032\,
            in3 => \N__44371\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNI7VNRE_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__64259\,
            in1 => \N__38994\,
            in2 => \_gnd_net_\,
            in3 => \N__39015\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec3_0_a2_i_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__38905\,
            in1 => \N__38822\,
            in2 => \_gnd_net_\,
            in3 => \N__26672\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1827_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_7_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43570\,
            in1 => \N__37873\,
            in2 => \N__24873\,
            in3 => \N__64260\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_863\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.electr_config_test_1_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__24818\,
            in1 => \N__45486\,
            in2 => \N__35487\,
            in3 => \N__45087\,
            lcout => s1_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65652\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_c_RNIA3PRE_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000100010"
        )
    port map (
            in0 => \N__64261\,
            in1 => \N__38949\,
            in2 => \_gnd_net_\,
            in3 => \N__38973\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNO_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__35482\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50746\,
            lcout => \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_i_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__50747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35483\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state4_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_1_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__40602\,
            in1 => \N__33654\,
            in2 => \_gnd_net_\,
            in3 => \N__36235\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_597\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__36236\,
            in1 => \N__25395\,
            in2 => \_gnd_net_\,
            in3 => \N__30969\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_596_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010101000"
        )
    port map (
            in0 => \N__35973\,
            in1 => \N__29855\,
            in2 => \N__25404\,
            in3 => \N__25401\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_id_prdata_1_4_u_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_26_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60901\,
            in2 => \_gnd_net_\,
            in3 => \N__59381\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_oZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65667\,
            ce => \N__54119\,
            sr => \N__62922\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIRLAS1_2_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39621\,
            in1 => \N__46911\,
            in2 => \_gnd_net_\,
            in3 => \N__39141\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_1615\,
            ltout => \cemf_module_64ch_ctrl_inst1.N_1615_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_2_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__64229\,
            in1 => \_gnd_net_\,
            in2 => \N__25389\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1832_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_0_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64228\,
            in2 => \_gnd_net_\,
            in3 => \N__36237\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1830_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_3_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010011100000000"
        )
    port map (
            in0 => \N__39142\,
            in1 => \N__39576\,
            in2 => \N__54351\,
            in3 => \N__64230\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_memZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIP15Q1_9_LC_9_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__29951\,
            in1 => \N__27572\,
            in2 => \N__25701\,
            in3 => \N__25080\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.csb_u_i_a2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.c_state_RNIGVSD3_0_LC_9_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001110101111"
        )
    port map (
            in0 => \N__25755\,
            in1 => \N__25635\,
            in2 => \N__25704\,
            in3 => \N__25697\,
            lcout => \N_1822_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_RNI0JD21_LC_9_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000010"
        )
    port map (
            in0 => \N__30243\,
            in1 => \N__27831\,
            in2 => \N__27798\,
            in3 => \N__29950\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.csb_u_i_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_1_LC_9_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101100000100"
        )
    port map (
            in0 => \N__25778\,
            in1 => \N__25971\,
            in2 => \N__26895\,
            in3 => \N__25991\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65691\,
            ce => 'H',
            sr => \N__62903\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_2_LC_9_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000010100"
        )
    port map (
            in0 => \N__26893\,
            in1 => \N__25958\,
            in2 => \N__25938\,
            in3 => \N__25781\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65691\,
            ce => 'H',
            sr => \N__62903\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_3_LC_9_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000110110000"
        )
    port map (
            in0 => \N__25779\,
            in1 => \N__26894\,
            in2 => \N__25925\,
            in3 => \N__25899\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65691\,
            ce => 'H',
            sr => \N__62903\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_0_LC_9_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000010010"
        )
    port map (
            in0 => \N__25447\,
            in1 => \N__26889\,
            in2 => \N__39345\,
            in3 => \N__25780\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65691\,
            ce => 'H',
            sr => \N__62903\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_0_LC_9_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000010010"
        )
    port map (
            in0 => \N__25616\,
            in1 => \N__25523\,
            in2 => \N__39346\,
            in3 => \N__25582\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.count_data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65691\,
            ce => 'H',
            sr => \N__62903\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_data_1_LC_9_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101100000100"
        )
    port map (
            in0 => \N__25581\,
            in1 => \N__25545\,
            in2 => \N__25534\,
            in3 => \N__25483\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_read_inst1.count_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65691\,
            ce => 'H',
            sr => \N__62903\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_c_0_LC_9_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25440\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_19_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_LUT4_0_LC_9_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25990\,
            in2 => \_gnd_net_\,
            in3 => \N__25965\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_LUT4_0_LC_9_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25957\,
            in2 => \_gnd_net_\,
            in3 => \N__25929\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_LUT4_0_LC_9_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25918\,
            in2 => \_gnd_net_\,
            in3 => \N__25893\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_data_4_LC_9_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000111000100"
        )
    port map (
            in0 => \N__26888\,
            in1 => \N__25883\,
            in2 => \N__25782\,
            in3 => \N__25890\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65706\,
            ce => 'H',
            sr => \N__62890\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_RNIU62F_LC_9_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__27209\,
            in1 => \N__27149\,
            in2 => \_gnd_net_\,
            in3 => \N__31344\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.csb_u_i_a2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_m8_0_a2_LC_9_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__30515\,
            in1 => \N__26990\,
            in2 => \N__30474\,
            in3 => \N__26933\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_RNIAVP33_14_LC_9_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__25857\,
            in1 => \N__25844\,
            in2 => \N__25812\,
            in3 => \N__25809\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.count_datae_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_0_0_LC_9_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27208\,
            in2 => \_gnd_net_\,
            in3 => \N__27143\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.N_217_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22_LC_9_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__27141\,
            in1 => \N__26142\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net\,
            ce => \N__27236\,
            sr => \N__62872\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_21_LC_9_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27138\,
            in2 => \_gnd_net_\,
            in3 => \N__26136\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net\,
            ce => \N__27236\,
            sr => \N__62872\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_20_LC_9_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27140\,
            in1 => \N__27279\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net\,
            ce => \N__27236\,
            sr => \N__62872\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_23_LC_9_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27139\,
            in2 => \_gnd_net_\,
            in3 => \N__26130\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.dout_op\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_22C_net\,
            ce => \N__27236\,
            sr => \N__62872\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_0_LC_9_22_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26038\,
            in1 => \N__26114\,
            in2 => \_gnd_net_\,
            in3 => \N__26100\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_9_22_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0\,
            clk => \N__65744\,
            ce => 'H',
            sr => \N__62864\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_1_LC_9_22_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26036\,
            in1 => \N__26096\,
            in2 => \_gnd_net_\,
            in3 => \N__26082\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1\,
            clk => \N__65744\,
            ce => 'H',
            sr => \N__62864\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_2_LC_9_22_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26039\,
            in1 => \N__26078\,
            in2 => \_gnd_net_\,
            in3 => \N__26064\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_2\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2\,
            clk => \N__65744\,
            ce => 'H',
            sr => \N__62864\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_3_LC_9_22_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26037\,
            in1 => \N__26057\,
            in2 => \_gnd_net_\,
            in3 => \N__26043\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_3\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_cry_3\,
            clk => \N__65744\,
            ce => 'H',
            sr => \N__62864\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bits_4_LC_9_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__26040\,
            in1 => \N__26009\,
            in2 => \_gnd_net_\,
            in3 => \N__26016\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.count_bitsZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65744\,
            ce => 'H',
            sr => \N__62864\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_31_LC_10_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011001100"
        )
    port map (
            in0 => \N__59555\,
            in1 => \N__28174\,
            in2 => \N__62060\,
            in3 => \N__33951\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_31,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65537\,
            ce => \N__32516\,
            sr => \N__62960\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_31_LC_10_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50401\,
            in2 => \N__26339\,
            in3 => \N__62044\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_203_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_17_LC_10_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26312\,
            in2 => \N__50409\,
            in3 => \N__57393\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_455_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_18_LC_10_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50397\,
            in2 => \N__26338\,
            in3 => \N__59834\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_454_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_19_LC_10_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__50396\,
            in1 => \N__26316\,
            in2 => \_gnd_net_\,
            in3 => \N__61613\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_453_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec2_0_a2_i_o2_LC_10_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__38736\,
            in1 => \N__38675\,
            in2 => \N__64317\,
            in3 => \N__64268\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_221_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_6_LC_10_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001000"
        )
    port map (
            in0 => \N__63582\,
            in1 => \N__26320\,
            in2 => \N__50395\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_463_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_i_0_8_LC_10_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__63102\,
            in1 => \_gnd_net_\,
            in2 => \N__26340\,
            in3 => \N__50355\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_462_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_5_LC_10_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__63657\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59558\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65557\,
            ce => \N__48722\,
            sr => \N__62954\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_6_LC_10_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59557\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63583\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65557\,
            ce => \N__48722\,
            sr => \N__62954\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_8_LC_10_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59556\,
            in2 => \_gnd_net_\,
            in3 => \N__63103\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65557\,
            ce => \N__48722\,
            sr => \N__62954\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.we_elec1_0_a2_i_LC_10_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__38891\,
            in1 => \N__38802\,
            in2 => \_gnd_net_\,
            in3 => \N__26655\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1829_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_1_LC_10_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__26613\,
            in1 => \N__52737\,
            in2 => \N__26601\,
            in3 => \N__52524\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_1_LC_10_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52222\,
            in2 => \N__26586\,
            in3 => \N__54603\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_1_LC_10_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__26583\,
            in1 => \N__44617\,
            in2 => \N__44127\,
            in3 => \N__38382\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_1_LC_10_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__28422\,
            in1 => \N__53331\,
            in2 => \N__26571\,
            in3 => \N__57800\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_1_LC_10_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27384\,
            in1 => \N__33540\,
            in2 => \N__26568\,
            in3 => \N__26565\,
            lcout => \I2C_top_level_inst1_s_data_oreg_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65571\,
            ce => \N__54522\,
            sr => \N__64971\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_5_LC_10_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51924\,
            in1 => \N__26559\,
            in2 => \N__28392\,
            in3 => \N__32197\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_5_LC_10_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27495\,
            in1 => \N__26745\,
            in2 => \N__26748\,
            in3 => \N__26703\,
            lcout => \I2C_top_level_inst1_s_data_oreg_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65595\,
            ce => \N__54516\,
            sr => \N__64967\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_5_LC_10_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__53012\,
            in1 => \N__32171\,
            in2 => \N__53315\,
            in3 => \N__42216\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_5_LC_10_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__26739\,
            in1 => \N__52772\,
            in2 => \N__26724\,
            in3 => \N__52521\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_5_LC_10_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52227\,
            in2 => \N__26706\,
            in3 => \N__32127\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_6_LC_10_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51860\,
            in1 => \N__26697\,
            in2 => \N__28359\,
            in3 => \N__33779\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_LC_10_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29146\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\,
            ce => 'H',
            sr => \N__62923\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m12_LC_10_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26691\,
            in2 => \_gnd_net_\,
            in3 => \N__28874\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQK6I1_LC_10_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__26682\,
            in1 => \N__29145\,
            in2 => \N__26676\,
            in3 => \N__32992\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_271\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_7_LC_10_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__29235\,
            in1 => \N__26778\,
            in2 => \_gnd_net_\,
            in3 => \N__30137\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\,
            ce => 'H',
            sr => \N__62923\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_6_LC_10_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28995\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\,
            ce => 'H',
            sr => \N__62923\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_5_LC_10_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\,
            ce => 'H',
            sr => \N__62923\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_4_LC_10_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28917\,
            in2 => \_gnd_net_\,
            in3 => \N__29234\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6C_net\,
            ce => 'H',
            sr => \N__62923\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17_LC_10_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27778\,
            in1 => \N__26766\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_18_LC_10_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27774\,
            in2 => \_gnd_net_\,
            in3 => \N__26772\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_13_LC_10_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27776\,
            in1 => \N__27006\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_16_LC_10_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27773\,
            in2 => \_gnd_net_\,
            in3 => \N__26760\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_22_LC_10_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__27779\,
            in1 => \N__26838\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_15_LC_10_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27772\,
            in2 => \_gnd_net_\,
            in3 => \N__26844\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_14_LC_10_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27777\,
            in1 => \N__26754\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_21_LC_10_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27775\,
            in2 => \_gnd_net_\,
            in3 => \N__26832\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_17C_net\,
            ce => \N__27707\,
            sr => \N__62904\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10_LC_10_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27784\,
            in2 => \_gnd_net_\,
            in3 => \N__26826\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_20_LC_10_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27781\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26784\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_9_LC_10_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27787\,
            in2 => \_gnd_net_\,
            in3 => \N__26820\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_8_LC_10_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__27783\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_11_LC_10_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27785\,
            in2 => \_gnd_net_\,
            in3 => \N__26814\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_23_LC_10_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26808\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.dout_op\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_19_LC_10_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__26790\,
            in1 => \N__27786\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_12_LC_10_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27780\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27012\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_dataZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.ser_data_10C_net\,
            ce => \N__27708\,
            sr => \N__62891\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_LC_10_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__51190\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.s_stop\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32743\,
            ce => 'H',
            sr => \N__31005\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_en_count_data_i_LC_10_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__30513\,
            in1 => \N__27000\,
            in2 => \N__30471\,
            in3 => \N__26937\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.en_count_data_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12_LC_10_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27145\,
            in1 => \N__27261\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\,
            ce => \N__27235\,
            sr => \N__62866\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_15_LC_10_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__27147\,
            in1 => \N__26856\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\,
            ce => \N__27235\,
            sr => \N__62866\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_13_LC_10_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27144\,
            in2 => \_gnd_net_\,
            in3 => \N__26868\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\,
            ce => \N__27235\,
            sr => \N__62866\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_14_LC_10_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27146\,
            in1 => \N__26862\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\,
            ce => \N__27235\,
            sr => \N__62866\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_16_LC_10_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__27148\,
            in1 => \N__26850\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_12C_net\,
            ce => \N__27235\,
            sr => \N__62866\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18_LC_10_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27132\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27267\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_19_LC_10_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27285\,
            in2 => \_gnd_net_\,
            in3 => \N__27136\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_8_LC_10_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27137\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_17_LC_10_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__27131\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27273\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_11_LC_10_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27243\,
            in2 => \_gnd_net_\,
            in3 => \N__27135\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_9_LC_10_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__27133\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27255\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_10_LC_10_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27249\,
            in2 => \_gnd_net_\,
            in3 => \N__27134\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_dataZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.ser_data_18C_net\,
            ce => \N__27237\,
            sr => \N__62860\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_op_inst1.c_state_RNIB86D_1_0_LC_10_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27207\,
            in2 => \_gnd_net_\,
            in3 => \N__27142\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.N_391\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIT2U5_16_LC_10_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__28181\,
            in1 => \N__29367\,
            in2 => \_gnd_net_\,
            in3 => \N__27966\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_config\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_8_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__32382\,
            in1 => \N__27021\,
            in2 => \N__53329\,
            in3 => \N__40698\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_1_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38315\,
            in1 => \N__57834\,
            in2 => \N__51946\,
            in3 => \N__54639\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_10_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37881\,
            in1 => \N__43577\,
            in2 => \N__27372\,
            in3 => \N__64267\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_830\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_3_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__53016\,
            in1 => \N__49676\,
            in2 => \N__53330\,
            in3 => \N__49641\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_3_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35553\,
            in1 => \N__27357\,
            in2 => \N__27360\,
            in3 => \N__27318\,
            lcout => \I2C_top_level_inst1_s_data_oreg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65558\,
            ce => \N__54520\,
            sr => \N__64974\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_3_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51892\,
            in1 => \N__27519\,
            in2 => \N__28500\,
            in3 => \N__49719\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__27351\,
            in1 => \N__52736\,
            in2 => \N__27336\,
            in3 => \N__52523\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_3_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52221\,
            in2 => \N__27321\,
            in3 => \N__33741\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_31_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__28449\,
            in1 => \N__51936\,
            in2 => \N__38505\,
            in3 => \N__27390\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_31_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52439\,
            in1 => \N__27312\,
            in2 => \N__27300\,
            in3 => \N__52779\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_31_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46134\,
            in2 => \N__27468\,
            in3 => \N__52232\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_31_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_31_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__27465\,
            in1 => \N__27456\,
            in2 => \N__27459\,
            in3 => \N__28152\,
            lcout => \I2C_top_level_inst1_s_data_oreg_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65572\,
            ce => \N__54517\,
            sr => \N__64972\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_31_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__53445\,
            in1 => \N__53257\,
            in2 => \N__46227\,
            in3 => \N__52987\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_27_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__27450\,
            in1 => \N__44533\,
            in2 => \N__61632\,
            in3 => \N__44326\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_28_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__44327\,
            in1 => \N__61544\,
            in2 => \N__44591\,
            in3 => \N__27438\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_29_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__27426\,
            in1 => \N__44534\,
            in2 => \N__61448\,
            in3 => \N__44328\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_3_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48057\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65583\,
            ce => \N__44105\,
            sr => \N__64968\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_30_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__44329\,
            in1 => \N__61318\,
            in2 => \N__44592\,
            in3 => \N__27414\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_31_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__27402\,
            in1 => \N__44541\,
            in2 => \N__61252\,
            in3 => \N__44330\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_3_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__44508\,
            in1 => \N__27540\,
            in2 => \N__27534\,
            in3 => \N__44333\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_4_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__44334\,
            in1 => \N__27510\,
            in2 => \N__33081\,
            in3 => \N__44509\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_4_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__30174\,
            in1 => \N__51866\,
            in2 => \N__27498\,
            in3 => \N__42486\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_5_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38302\,
            in1 => \N__37705\,
            in2 => \N__32229\,
            in3 => \N__41127\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_4_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__53015\,
            in1 => \N__42252\,
            in2 => \N__53319\,
            in3 => \N__29697\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_4_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__28602\,
            in1 => \N__52234\,
            in2 => \_gnd_net_\,
            in3 => \N__33703\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_4_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__28137\,
            in1 => \N__27489\,
            in2 => \N__27483\,
            in3 => \N__27480\,
            lcout => \I2C_top_level_inst1_s_data_oreg_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65605\,
            ce => \N__54507\,
            sr => \N__64965\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_0_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27599\,
            in1 => \N__27612\,
            in2 => \_gnd_net_\,
            in3 => \N__27474\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_15_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0\,
            clk => \N__65618\,
            ce => 'H',
            sr => \N__62905\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_1_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27596\,
            in1 => \N__27639\,
            in2 => \_gnd_net_\,
            in3 => \N__27471\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1\,
            clk => \N__65618\,
            ce => 'H',
            sr => \N__62905\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_2_LC_11_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27600\,
            in1 => \N__27654\,
            in2 => \_gnd_net_\,
            in3 => \N__27687\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_2\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2\,
            clk => \N__65618\,
            ce => 'H',
            sr => \N__62905\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_3_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__27597\,
            in1 => \N__27627\,
            in2 => \_gnd_net_\,
            in3 => \N__27684\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_3\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_cry_3\,
            clk => \N__65618\,
            ce => 'H',
            sr => \N__62905\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bits_4_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__27666\,
            in1 => \N__27598\,
            in2 => \_gnd_net_\,
            in3 => \N__27681\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.count_bitsZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65618\,
            ce => 'H',
            sr => \N__62905\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1_LC_11_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27822\,
            in2 => \_gnd_net_\,
            in3 => \N__27771\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net\,
            ce => 'H',
            sr => \N__62892\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_0_LC_11_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__27770\,
            in1 => \_gnd_net_\,
            in2 => \N__27827\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ns_1_0__m7_3_LC_11_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__27665\,
            in1 => \N__27653\,
            in2 => \N__27642\,
            in3 => \N__27638\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m7_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_0_LC_11_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27626\,
            in2 => \N__27615\,
            in3 => \N__27611\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_1C_net\,
            ce => 'H',
            sr => \N__62892\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_LC_11_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27817\,
            in2 => \_gnd_net_\,
            in3 => \N__27768\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_d_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_1_0_LC_11_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__27823\,
            in1 => \N__27788\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_RNIDOFE_0_0_LC_11_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27821\,
            in2 => \_gnd_net_\,
            in3 => \N__27769\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_43_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIQO531_LC_11_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28956\,
            in1 => \N__29074\,
            in2 => \N__30122\,
            in3 => \N__30081\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_274_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9_LC_11_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__29075\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62882\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_LC_11_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__28957\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62882\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_8_LC_11_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29222\,
            in2 => \_gnd_net_\,
            in3 => \N__28887\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62882\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_16_LC_11_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30034\,
            in2 => \_gnd_net_\,
            in3 => \N__29221\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62882\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_17_LC_11_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29099\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62882\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_3_LC_11_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__29061\,
            in1 => \N__29037\,
            in2 => \N__29006\,
            in3 => \N__28958\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_ret_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62882\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIE8O3_0_LC_11_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__27869\,
            in1 => \N__27884\,
            in2 => \N__27855\,
            in3 => \N__29106\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_1996_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3_LC_11_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101011111111"
        )
    port map (
            in0 => \N__28909\,
            in1 => \_gnd_net_\,
            in2 => \N__27690\,
            in3 => \N__27912\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net\,
            ce => 'H',
            sr => \N__62874\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_1_LC_11_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__29942\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35853\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net\,
            ce => 'H',
            sr => \N__62874\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_LC_11_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29190\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_3C_net\,
            ce => 'H',
            sr => \N__62874\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_1_RNIFTTJ_LC_11_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27911\,
            in2 => \_gnd_net_\,
            in3 => \N__28908\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_287_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1OR71_LC_11_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27900\,
            in2 => \N__27888\,
            in3 => \N__29941\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_0_LC_11_19_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28861\,
            in1 => \N__27885\,
            in2 => \_gnd_net_\,
            in3 => \N__27873\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_19_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0\,
            clk => \N__65669\,
            ce => 'H',
            sr => \N__62867\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_1_LC_11_19_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28847\,
            in1 => \N__27870\,
            in2 => \_gnd_net_\,
            in3 => \N__27858\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1\,
            clk => \N__65669\,
            ce => 'H',
            sr => \N__62867\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_2_LC_11_19_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28862\,
            in1 => \N__27854\,
            in2 => \_gnd_net_\,
            in3 => \N__27840\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_2\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2\,
            clk => \N__65669\,
            ce => 'H',
            sr => \N__62867\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_3_LC_11_19_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__28848\,
            in1 => \N__29118\,
            in2 => \_gnd_net_\,
            in3 => \N__27837\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_3\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_cry_3\,
            clk => \N__65669\,
            ce => 'H',
            sr => \N__62867\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_4_LC_11_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__29130\,
            in1 => \N__28849\,
            in2 => \_gnd_net_\,
            in3 => \N__27834\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bitsZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65669\,
            ce => 'H',
            sr => \N__62867\
        );

    \cemf_module_64ch_ctrl_inst1.ch_cnt_0_LC_11_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__29256\,
            in1 => \N__36873\,
            in2 => \_gnd_net_\,
            in3 => \N__27978\,
            lcout => \cemf_module_64ch_ctrl_inst1.ch_cntZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65694\,
            ce => 'H',
            sr => \N__62854\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_0_LC_11_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27996\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65714\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNI07M9_LC_11_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__27977\,
            in1 => \N__29405\,
            in2 => \_gnd_net_\,
            in3 => \N__27965\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_410_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.N_410_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m56_i_LC_11_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111100010011"
        )
    port map (
            in0 => \N__30596\,
            in1 => \N__31456\,
            in2 => \N__27954\,
            in3 => \N__31479\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_68_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.N_68_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_i_i_0_o2_i_o2_0_4_LC_11_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__29389\,
            in1 => \N__35762\,
            in2 => \N__27951\,
            in3 => \N__29363\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_reti_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_8_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37707\,
            in1 => \N__53011\,
            in2 => \N__28803\,
            in3 => \N__40731\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_8_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38316\,
            in1 => \N__40759\,
            in2 => \N__51951\,
            in3 => \N__41025\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_8_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__27948\,
            in1 => \N__52744\,
            in2 => \N__27933\,
            in3 => \N__52527\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_8_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52203\,
            in2 => \N__27915\,
            in3 => \N__40833\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_8_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__28125\,
            in1 => \N__28119\,
            in2 => \N__28113\,
            in3 => \N__28110\,
            lcout => \I2C_top_level_inst1_s_data_oreg_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65527\,
            ce => \N__54523\,
            sr => \N__64985\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_14_LC_12_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28104\,
            in1 => \N__52761\,
            in2 => \N__28089\,
            in3 => \N__52520\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_14_LC_12_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__52206\,
            in1 => \_gnd_net_\,
            in2 => \N__28071\,
            in3 => \N__32097\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_14_LC_12_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__44368\,
            in1 => \N__63568\,
            in2 => \N__44662\,
            in3 => \N__28068\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_14_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__28698\,
            in1 => \N__51950\,
            in2 => \N__28053\,
            in3 => \N__38487\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_14_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__34968\,
            in1 => \N__30771\,
            in2 => \N__28050\,
            in3 => \N__28047\,
            lcout => \I2C_top_level_inst1_s_data_oreg_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65538\,
            ce => \N__54521\,
            sr => \N__64982\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_22_LC_12_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28041\,
            in1 => \N__44635\,
            in2 => \N__58440\,
            in3 => \N__44367\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_30_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__38550\,
            in1 => \N__53271\,
            in2 => \N__46293\,
            in3 => \N__53004\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_30_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28026\,
            in1 => \N__52780\,
            in2 => \N__28011\,
            in3 => \N__52445\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_30_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34026\,
            in2 => \N__28227\,
            in3 => \N__52233\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_30_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_30_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__28200\,
            in1 => \N__28224\,
            in2 => \N__28218\,
            in3 => \N__28206\,
            lcout => \I2C_top_level_inst1_s_data_oreg_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65547\,
            ce => \N__54518\,
            sr => \N__64978\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_30_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__51925\,
            in1 => \N__28470\,
            in2 => \N__38097\,
            in3 => \N__28215\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_30_LC_12_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28584\,
            in1 => \N__38276\,
            in2 => \N__28194\,
            in3 => \N__37689\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_30_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__62125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59441\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65559\,
            ce => \N__45572\,
            sr => \N__62932\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_31_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28182\,
            in1 => \N__38277\,
            in2 => \N__28146\,
            in3 => \N__37690\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_31_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__62024\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59442\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65559\,
            ce => \N__45572\,
            sr => \N__62932\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_4_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38268\,
            in1 => \N__37688\,
            in2 => \N__28566\,
            in3 => \N__28325\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_4_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63775\,
            in2 => \_gnd_net_\,
            in3 => \N__59443\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65559\,
            ce => \N__45572\,
            sr => \N__62932\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMAFN1_LC_12_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55198\,
            in1 => \N__55438\,
            in2 => \N__33714\,
            in3 => \N__28321\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9GQL2_LC_12_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__33710\,
            in1 => \N__54954\,
            in2 => \N__28326\,
            in3 => \N__54757\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_26_LC_12_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__28311\,
            in1 => \N__37844\,
            in2 => \_gnd_net_\,
            in3 => \N__66815\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_26_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__28299\,
            in1 => \N__32362\,
            in2 => \N__28281\,
            in3 => \N__34050\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_1_26_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_26_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__33432\,
            in1 => \N__28263\,
            in2 => \N__28257\,
            in3 => \N__28254\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_a3_1_3_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_26_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000101"
        )
    port map (
            in0 => \N__57249\,
            in1 => \_gnd_net_\,
            in2 => \N__66819\,
            in3 => \N__59851\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66814\,
            in2 => \_gnd_net_\,
            in3 => \N__57248\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1872_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_21_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64252\,
            in1 => \N__32363\,
            in2 => \N__43576\,
            in3 => \N__28242\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNITSQ5D_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__32361\,
            in1 => \N__43533\,
            in2 => \_gnd_net_\,
            in3 => \N__64251\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1318\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_9_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64208\,
            in1 => \N__28542\,
            in2 => \N__43562\,
            in3 => \N__37869\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_841\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_29_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37863\,
            in1 => \N__28527\,
            in2 => \N__43575\,
            in3 => \N__64202\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_632\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_3_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64204\,
            in1 => \N__28512\,
            in2 => \N__43560\,
            in3 => \N__37866\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_907\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_30_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37864\,
            in1 => \N__43491\,
            in2 => \N__28488\,
            in3 => \N__64205\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_621\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_31_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64201\,
            in1 => \N__28461\,
            in2 => \N__43559\,
            in3 => \N__37865\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_610\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_1_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32360\,
            in1 => \N__43492\,
            in2 => \N__28437\,
            in3 => \N__64207\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_5_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64206\,
            in1 => \N__28410\,
            in2 => \N__43561\,
            in3 => \N__37868\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_885\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_6_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37867\,
            in1 => \N__43487\,
            in2 => \N__28377\,
            in3 => \N__64203\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_874\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_9_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__52739\,
            in1 => \N__28347\,
            in2 => \N__28656\,
            in3 => \N__52370\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_4_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52371\,
            in1 => \N__28635\,
            in2 => \N__28620\,
            in3 => \N__52740\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_9_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__44590\,
            in1 => \N__28596\,
            in2 => \N__61862\,
            in3 => \N__44369\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_0_LC_12_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101010"
        )
    port map (
            in0 => \N__40060\,
            in1 => \N__61971\,
            in2 => \N__59445\,
            in3 => \N__33932\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_0_6_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__40000\,
            in1 => \N__40059\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_349\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_28_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__35651\,
            in1 => \N__59275\,
            in2 => \N__62376\,
            in3 => \N__33933\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_28,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_29_LC_12_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__33929\,
            in1 => \N__62259\,
            in2 => \N__59446\,
            in3 => \N__35603\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_29,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_3_LC_12_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__63914\,
            in1 => \N__59276\,
            in2 => \N__35573\,
            in3 => \N__33934\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_30_LC_12_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__33930\,
            in1 => \N__62147\,
            in2 => \N__59447\,
            in3 => \N__28583\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_30,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_4_LC_12_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__63822\,
            in1 => \N__59277\,
            in2 => \N__28562\,
            in3 => \N__33935\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_8_LC_12_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33931\,
            in1 => \N__28796\,
            in2 => \N__59448\,
            in3 => \N__63144\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65606\,
            ce => \N__32517\,
            sr => \N__62893\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_0_LC_12_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37805\,
            in1 => \N__43540\,
            in2 => \N__28782\,
            in3 => \N__64213\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_940\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_11_LC_12_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37806\,
            in1 => \N__43545\,
            in2 => \N__28764\,
            in3 => \N__64217\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_819\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_12_LC_12_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64215\,
            in1 => \N__28749\,
            in2 => \N__43579\,
            in3 => \N__37807\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_808\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_13_LC_12_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37808\,
            in1 => \N__43541\,
            in2 => \N__28731\,
            in3 => \N__64216\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_797\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_14_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64218\,
            in1 => \N__28713\,
            in2 => \N__43580\,
            in3 => \N__37809\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_786\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_15_LC_12_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37810\,
            in1 => \N__43549\,
            in2 => \N__28686\,
            in3 => \N__64219\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_775\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_20_LC_12_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64214\,
            in1 => \N__28665\,
            in2 => \N__43578\,
            in3 => \N__32364\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_283\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIT5I21_16_LC_12_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__29095\,
            in1 => \N__32973\,
            in2 => \N__29041\,
            in3 => \N__29999\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_549_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_LC_12_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29033\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_i_3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62875\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m10_LC_12_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28941\,
            in2 => \_gnd_net_\,
            in3 => \N__28819\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_286_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_19_LC_12_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28935\,
            in2 => \N__28920\,
            in3 => \N__29224\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62875\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_11_LC_12_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111111"
        )
    port map (
            in0 => \N__29223\,
            in1 => \_gnd_net_\,
            in2 => \N__30084\,
            in3 => \N__30121\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62875\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_0_LC_12_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__28820\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30077\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m15_LC_12_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__28910\,
            in1 => \N__30036\,
            in2 => \N__28890\,
            in3 => \N__28886\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_277_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_20_LC_12_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__28821\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29225\,
            lcout => \cemf_module_64ch_ctrl_inst1.end_conf_b\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62875\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_RNI63PT_LC_12_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__28809\,
            in1 => \N__30026\,
            in2 => \N__30054\,
            in3 => \N__29166\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5_LC_12_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29168\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\,
            ce => 'H',
            sr => \N__62868\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_12_LC_12_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29219\,
            in2 => \_gnd_net_\,
            in3 => \N__30083\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\,
            ce => 'H',
            sr => \N__62868\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_15_LC_12_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011111111"
        )
    port map (
            in0 => \N__29220\,
            in1 => \_gnd_net_\,
            in2 => \N__30035\,
            in3 => \N__30052\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\,
            ce => 'H',
            sr => \N__62868\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_13_LC_12_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29169\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\,
            ce => 'H',
            sr => \N__62868\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_LC_12_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__29178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_i_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_5C_net\,
            ce => 'H',
            sr => \N__62868\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_1_LC_12_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__29189\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29177\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIHNKP_12_LC_12_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__29167\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__29154\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.count_bits_RNIF6G1_4_LC_12_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29129\,
            in2 => \_gnd_net_\,
            in3 => \N__29117\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_i_a2_1_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIPVKP_16_LC_12_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29100\,
            in2 => \_gnd_net_\,
            in3 => \N__29079\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m45_0_LC_12_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__29060\,
            in1 => \N__29048\,
            in2 => \N__29007\,
            in3 => \N__28965\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_276i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_0_LC_12_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31090\,
            in1 => \N__30285\,
            in2 => \_gnd_net_\,
            in3 => \N__29271\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_12_20_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0\,
            clk => \N__65670\,
            ce => 'H',
            sr => \N__62855\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_1_LC_12_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31087\,
            in1 => \N__30300\,
            in2 => \_gnd_net_\,
            in3 => \N__29268\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1\,
            clk => \N__65670\,
            ce => 'H',
            sr => \N__62855\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_2_LC_12_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31091\,
            in1 => \N__30312\,
            in2 => \_gnd_net_\,
            in3 => \N__29265\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_2\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2\,
            clk => \N__65670\,
            ce => 'H',
            sr => \N__62855\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_3_LC_12_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__31088\,
            in1 => \N__30324\,
            in2 => \_gnd_net_\,
            in3 => \N__29262\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_3\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_cry_3\,
            clk => \N__65670\,
            ce => 'H',
            sr => \N__62855\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_4_LC_12_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__30336\,
            in1 => \N__31089\,
            in2 => \_gnd_net_\,
            in3 => \N__29259\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bitsZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65670\,
            ce => 'H',
            sr => \N__62855\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIFUVN_LC_12_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__29390\,
            in1 => \N__40037\,
            in2 => \_gnd_net_\,
            in3 => \N__32825\,
            lcout => \cemf_module_64ch_ctrl_inst1.en_ch_cnt_0_a2_0_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_RNO_0_LC_12_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__29250\,
            in1 => \N__29391\,
            in2 => \N__31455\,
            in3 => \N__36839\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un40_0_a2_4_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_m3_i_0_a2_LC_12_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101000101010"
        )
    port map (
            in0 => \N__32770\,
            in1 => \N__36869\,
            in2 => \N__36843\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1945\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_LC_12_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__30350\,
            in1 => \N__29366\,
            in2 => \N__35763\,
            in3 => \N__29394\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1851_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65695\,
            ce => 'H',
            sr => \N__62844\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_sync_LC_12_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__29412\,
            in1 => \N__31314\,
            in2 => \_gnd_net_\,
            in3 => \N__29406\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_syncZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65695\,
            ce => 'H',
            sr => \N__62844\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_LC_12_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__30349\,
            in1 => \N__29393\,
            in2 => \_gnd_net_\,
            in3 => \N__29365\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1844\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65695\,
            ce => 'H',
            sr => \N__62844\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_17_LC_12_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29392\,
            in2 => \_gnd_net_\,
            in3 => \N__29364\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65695\,
            ce => 'H',
            sr => \N__62844\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_16_LC_12_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35757\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65695\,
            ce => 'H',
            sr => \N__62844\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIANE51_11_LC_12_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101010101"
        )
    port map (
            in0 => \N__36552\,
            in1 => \N__63281\,
            in2 => \N__41529\,
            in3 => \N__50994\,
            lcout => sda_o,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_22_LC_13_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__52223\,
            in1 => \N__29277\,
            in2 => \_gnd_net_\,
            in3 => \N__38607\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_22_LC_13_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__30744\,
            in1 => \N__29316\,
            in2 => \N__29319\,
            in3 => \N__29532\,
            lcout => \I2C_top_level_inst1_s_data_oreg_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65518\,
            ce => \N__54524\,
            sr => \N__64996\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_22_LC_13_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__42279\,
            in1 => \N__53010\,
            in2 => \N__53328\,
            in3 => \N__38532\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_22_LC_13_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__29310\,
            in1 => \N__52743\,
            in2 => \N__29295\,
            in3 => \N__52438\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_22_LC_13_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51903\,
            in1 => \N__29538\,
            in2 => \N__33324\,
            in3 => \N__38436\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_28_LC_13_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__54177\,
            in1 => \N__53270\,
            in2 => \N__40623\,
            in3 => \N__52994\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_28_LC_13_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__29526\,
            in1 => \N__52768\,
            in2 => \N__29514\,
            in3 => \N__52486\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_28_LC_13_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49128\,
            in2 => \N__29496\,
            in3 => \N__52213\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_28_LC_13_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35631\,
            in1 => \N__29493\,
            in2 => \N__29487\,
            in3 => \N__29472\,
            lcout => \I2C_top_level_inst1_s_data_oreg_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65528\,
            ce => \N__54519\,
            sr => \N__64986\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_28_LC_13_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__29823\,
            in1 => \N__51904\,
            in2 => \N__48795\,
            in3 => \N__29484\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_15_LC_13_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__29466\,
            in1 => \N__52700\,
            in2 => \N__29448\,
            in3 => \N__52488\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_15_LC_13_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__52182\,
            in1 => \_gnd_net_\,
            in2 => \N__29430\,
            in3 => \N__46605\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_15_LC_13_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__44407\,
            in1 => \N__63481\,
            in2 => \N__44659\,
            in3 => \N__29427\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_15_LC_13_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__29661\,
            in1 => \N__51859\,
            in2 => \N__29649\,
            in3 => \N__48581\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_15_LC_13_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__34923\,
            in1 => \N__30759\,
            in2 => \N__29646\,
            in3 => \N__29643\,
            lcout => \I2C_top_level_inst1_s_data_oreg_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65539\,
            ce => \N__54513\,
            sr => \N__64983\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_23_LC_13_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__29637\,
            in1 => \N__44624\,
            in2 => \N__57475\,
            in3 => \N__44406\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_17_LC_13_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__52742\,
            in1 => \N__29622\,
            in2 => \N__29604\,
            in3 => \N__52487\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_17_LC_13_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52215\,
            in2 => \N__29586\,
            in3 => \N__46563\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_17_LC_13_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__44332\,
            in1 => \N__29583\,
            in2 => \N__46507\,
            in3 => \N__44548\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_17_LC_13_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__33135\,
            in1 => \N__51919\,
            in2 => \N__29568\,
            in3 => \N__51624\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_17_LC_13_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35316\,
            in1 => \N__30804\,
            in2 => \N__29565\,
            in3 => \N__29562\,
            lcout => \I2C_top_level_inst1_s_data_oreg_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65548\,
            ce => \N__54510\,
            sr => \N__64979\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_25_LC_13_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__44547\,
            in1 => \N__29556\,
            in2 => \N__57374\,
            in3 => \N__44331\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIUMB92_17_LC_13_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__57978\,
            in1 => \N__58156\,
            in2 => \N__42481\,
            in3 => \N__29689\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3Q5_LC_13_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60474\,
            in1 => \N__42247\,
            in2 => \N__29715\,
            in3 => \N__29712\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI7A3QZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_4_LC_13_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63785\,
            in2 => \_gnd_net_\,
            in3 => \N__59444\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65560\,
            ce => \N__54113\,
            sr => \N__62914\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0FK93_LC_13_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100110001"
        )
    port map (
            in0 => \N__42482\,
            in1 => \N__42248\,
            in2 => \N__46041\,
            in3 => \N__45867\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRL7_LC_13_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__53959\,
            in1 => \N__29706\,
            in2 => \N__29700\,
            in3 => \N__29690\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISHRLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7LCO7_LC_13_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53672\,
            in1 => \_gnd_net_\,
            in2 => \N__29676\,
            in3 => \N__30905\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0RV43_LC_13_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__45866\,
            in1 => \N__45992\,
            in2 => \N__38077\,
            in3 => \N__46270\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_6_LC_13_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__52220\,
            in1 => \N__29760\,
            in2 => \_gnd_net_\,
            in3 => \N__33678\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_6_LC_13_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__32049\,
            in1 => \N__29808\,
            in2 => \N__29673\,
            in3 => \N__29670\,
            lcout => \I2C_top_level_inst1_s_data_oreg_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65573\,
            ce => \N__54503\,
            sr => \N__64973\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_6_LC_13_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__31985\,
            in1 => \N__53281\,
            in2 => \N__53013\,
            in3 => \N__42175\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_6_LC_13_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__52741\,
            in1 => \N__29802\,
            in2 => \N__29781\,
            in3 => \N__52437\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_9_LC_13_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51906\,
            in1 => \N__29754\,
            in2 => \N__29748\,
            in3 => \N__49386\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_9_LC_13_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__30885\,
            in1 => \N__29724\,
            in2 => \N__29739\,
            in3 => \N__29730\,
            lcout => \I2C_top_level_inst1_s_data_oreg_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65584\,
            ce => \N__54502\,
            sr => \N__64969\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_9_LC_13_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__29736\,
            in1 => \N__52216\,
            in2 => \_gnd_net_\,
            in3 => \N__46641\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_9_LC_13_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52990\,
            in1 => \N__49842\,
            in2 => \N__53316\,
            in3 => \N__49423\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI0PB92_17_LC_13_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__58112\,
            in1 => \N__57941\,
            in2 => \N__32172\,
            in3 => \N__32207\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3Q5_LC_13_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60472\,
            in1 => \N__42208\,
            in2 => \N__29718\,
            in3 => \N__29814\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNICF3QZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6_LC_13_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__60149\,
            in1 => \N__29862\,
            in2 => \_gnd_net_\,
            in3 => \N__29888\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net\,
            ce => \N__59940\,
            sr => \N__62883\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI2RB92_17_LC_13_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100001011"
        )
    port map (
            in0 => \N__57942\,
            in1 => \N__31989\,
            in2 => \N__33786\,
            in3 => \N__58113\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3Q5_LC_13_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111110111111"
        )
    port map (
            in0 => \N__42177\,
            in1 => \N__32001\,
            in2 => \N__29895\,
            in3 => \N__60473\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIHK3QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNII2U76_LC_13_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60355\,
            in1 => \_gnd_net_\,
            in2 => \N__29892\,
            in3 => \N__29889\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIDTT76_LC_13_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__29877\,
            in1 => \N__60354\,
            in2 => \_gnd_net_\,
            in3 => \N__29871\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_5_LC_13_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__30822\,
            in1 => \_gnd_net_\,
            in2 => \N__29865\,
            in3 => \N__60148\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_6C_net\,
            ce => \N__59940\,
            sr => \N__62883\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIPJAS1_1_LC_13_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39653\,
            in1 => \N__46817\,
            in2 => \_gnd_net_\,
            in3 => \N__39140\,
            lcout => \N_1614\,
            ltout => \N_1614_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_a2_LC_13_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29856\,
            in2 => \N__29841\,
            in3 => \N__36201\,
            lcout => \N_979\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_28_LC_13_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43512\,
            in1 => \N__29838\,
            in2 => \N__37823\,
            in3 => \N__64153\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_643\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOCFN1_LC_13_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55351\,
            in1 => \N__55113\,
            in2 => \N__41125\,
            in3 => \N__32123\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_4_LC_13_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__43511\,
            in1 => \N__30186\,
            in2 => \N__37824\,
            in3 => \N__64152\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_896\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNIR6CE2_0_LC_13_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010100000"
        )
    port map (
            in0 => \N__30259\,
            in1 => \N__29920\,
            in2 => \N__29988\,
            in3 => \N__35854\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_291_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_LC_13_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30162\,
            in3 => \N__30159\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_retZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net\,
            ce => 'H',
            sr => \N__62869\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4_RNIB3H2_LC_13_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30150\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.N_272_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_RNO_0_0_LC_13_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30242\,
            in1 => \N__29986\,
            in2 => \N__30264\,
            in3 => \N__30989\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_0_LC_13_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1000100011111000"
        )
    port map (
            in0 => \N__30238\,
            in1 => \N__32982\,
            in2 => \N__30144\,
            in3 => \N__35856\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.c_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net\,
            ce => 'H',
            sr => \N__62869\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5EOM1_LC_13_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30141\,
            in1 => \N__30123\,
            in2 => \N__30099\,
            in3 => \N__30082\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ns_a2_0_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_LC_13_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__30053\,
            in1 => \N__30033\,
            in2 => \N__30003\,
            in3 => \N__30000\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_259_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_8_LC_13_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100110000000000"
        )
    port map (
            in0 => \N__35855\,
            in1 => \N__29987\,
            in2 => \N__29940\,
            in3 => \N__30260\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_291\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.c_state_ret_4C_net\,
            ce => 'H',
            sr => \N__62869\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_LC_13_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30555\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\,
            ce => 'H',
            sr => \N__62861\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3_RNIJA1F_LC_13_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30219\,
            in2 => \_gnd_net_\,
            in3 => \N__31123\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_o3_i_a2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI0RBC1_LC_13_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__30210\,
            in1 => \N__30554\,
            in2 => \N__30213\,
            in3 => \N__32884\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_340\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_LC_13_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__30203\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\,
            ce => 'H',
            sr => \N__62861\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_5_LC_13_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30556\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\,
            ce => 'H',
            sr => \N__62861\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_6_LC_13_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30204\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\,
            ce => 'H',
            sr => \N__62861\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI496Q_5_LC_13_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30380\,
            in2 => \_gnd_net_\,
            in3 => \N__30202\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m20_0_a2_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_10_LC_13_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__30381\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_3C_net\,
            ce => 'H',
            sr => \N__62861\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11_LC_13_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__30192\,
            in1 => \N__31029\,
            in2 => \_gnd_net_\,
            in3 => \N__31255\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            ce => 'H',
            sr => \N__62856\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_4_LC_13_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31256\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31385\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            ce => 'H',
            sr => \N__62856\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNIDC2S_4_LC_13_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30335\,
            in2 => \_gnd_net_\,
            in3 => \N__30323\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ns_i_a2_1_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.count_bits_RNI9N562_0_LC_13_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__30311\,
            in1 => \N__30299\,
            in2 => \N__30288\,
            in3 => \N__30284\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1987_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_3_LC_13_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101011001111"
        )
    port map (
            in0 => \N__31386\,
            in1 => \N__30270\,
            in2 => \N__30273\,
            in3 => \N__31364\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            ce => 'H',
            sr => \N__62856\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_8_LC_13_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31257\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31124\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            ce => 'H',
            sr => \N__62856\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_2_LC_13_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32568\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            ce => 'H',
            sr => \N__62856\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_10_LC_13_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__32567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_11C_net\,
            ce => 'H',
            sr => \N__62856\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIF2FF_12_LC_13_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__31283\,
            in1 => \N__30557\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_8_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_LC_13_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31086\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60127\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2FZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_RNION2F1_0_LC_13_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__30561\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1973_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_1_0_LC_13_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__30558\,
            in1 => \N__31336\,
            in2 => \_gnd_net_\,
            in3 => \N__32697\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNO_0_0_LC_13_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__31284\,
            in1 => \N__30537\,
            in2 => \N__30531\,
            in3 => \N__31161\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m52_0_a2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_LC_13_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31162\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5C_net\,
            ce => 'H',
            sr => \N__62849\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIO27J_LC_13_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__30363\,
            in1 => \N__31026\,
            in2 => \N__30528\,
            in3 => \N__31160\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_274\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9_LC_13_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31173\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62845\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_read_inst1.c_state_10_LC_13_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30519\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_state_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62845\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_7_LC_13_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30379\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_9C_net\,
            ce => 'H',
            sr => \N__62845\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_19_LC_13_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30354\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_state_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65681\,
            ce => 'H',
            sr => \N__62838\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_LC_13_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000101110111011"
        )
    port map (
            in0 => \N__30609\,
            in1 => \N__30595\,
            in2 => \N__31458\,
            in3 => \N__31478\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65681\,
            ce => 'H',
            sr => \N__62838\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.m59_i_LC_13_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000111"
        )
    port map (
            in0 => \N__31451\,
            in1 => \N__31477\,
            in2 => \N__30597\,
            in3 => \N__30608\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_1816_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_7_LC_13_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40111\,
            in2 => \_gnd_net_\,
            in3 => \N__40001\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_state_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65681\,
            ce => 'H',
            sr => \N__62838\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_0_LC_13_23_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34272\,
            in2 => \N__31590\,
            in3 => \N__31589\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_0\,
            ltout => OPEN,
            carryin => \bfn_13_23_0_\,
            carryout => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_1_LC_13_23_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34190\,
            in2 => \_gnd_net_\,
            in3 => \N__30576\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_1\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_0\,
            carryout => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_2_LC_13_23_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34244\,
            in2 => \_gnd_net_\,
            in3 => \N__30573\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_2\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_1\,
            carryout => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_bit_counter_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0_3_LC_13_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34217\,
            in2 => \_gnd_net_\,
            in3 => \N__30570\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNO_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetter_LC_13_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50820\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_resetterZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47997\,
            ce => 'H',
            sr => \N__62829\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_RNO_LC_13_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__30567\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35457\,
            lcout => \I2C_top_level_inst1.I2C_Control_StartUp_inst.rst_neg_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.start_detect_LC_13_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51186\,
            lcout => \I2C_top_level_inst1.s_start\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_Control_StartUp_inst.start_detectC_net\,
            ce => 'H',
            sr => \N__30753\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_22_LC_14_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__37701\,
            in1 => \N__42681\,
            in2 => \N__38304\,
            in3 => \N__30867\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_2_LC_14_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__30738\,
            in1 => \N__44675\,
            in2 => \N__32925\,
            in3 => \N__44418\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_13_LC_14_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__30720\,
            in1 => \N__52760\,
            in2 => \N__30708\,
            in3 => \N__52471\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_13_LC_14_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52205\,
            in2 => \N__30690\,
            in3 => \N__46173\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_13_LC_14_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__30687\,
            in1 => \N__44663\,
            in2 => \N__63670\,
            in3 => \N__44413\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_13_LC_14_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__30672\,
            in1 => \N__51902\,
            in2 => \N__30657\,
            in3 => \N__38079\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_13_LC_14_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35004\,
            in1 => \N__30654\,
            in2 => \N__30648\,
            in3 => \N__30780\,
            lcout => \I2C_top_level_inst1_s_data_oreg_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65522\,
            ce => \N__54514\,
            sr => \N__64992\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_18_LC_14_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__30645\,
            in1 => \N__38373\,
            in2 => \N__30630\,
            in3 => \N__52701\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_18_LC_14_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52186\,
            in2 => \N__30798\,
            in3 => \N__49173\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_18_LC_14_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__33498\,
            in1 => \N__30786\,
            in2 => \N__30795\,
            in3 => \N__30792\,
            lcout => \I2C_top_level_inst1_s_data_oreg_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65529\,
            ce => \N__54511\,
            sr => \N__64987\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_18_LC_14_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__32412\,
            in1 => \N__38303\,
            in2 => \N__31626\,
            in3 => \N__48862\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_18_LC_14_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__53258\,
            in1 => \N__51438\,
            in2 => \N__51905\,
            in3 => \N__51402\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_10_LC_14_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__49340\,
            in1 => \N__52923\,
            in2 => \N__53256\,
            in3 => \N__49269\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_11_LC_14_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52925\,
            in1 => \N__46380\,
            in2 => \N__53262\,
            in3 => \N__42527\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_13_LC_14_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__53179\,
            in1 => \N__46272\,
            in2 => \N__40896\,
            in3 => \N__52924\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_14_LC_14_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52922\,
            in1 => \N__33564\,
            in2 => \N__53430\,
            in3 => \N__53175\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_15_LC_14_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__53180\,
            in1 => \N__52926\,
            in2 => \N__53382\,
            in3 => \N__46212\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_17_LC_14_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__53181\,
            in1 => \N__52927\,
            in2 => \N__54165\,
            in3 => \N__51586\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_1_LC_14_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61861\,
            in2 => \_gnd_net_\,
            in3 => \N__59142\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_2_LC_14_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59145\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61729\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_3_LC_14_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__63910\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59149\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_5_LC_14_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63645\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_6_LC_14_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63526\,
            in2 => \_gnd_net_\,
            in3 => \N__59143\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_7_LC_14_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59147\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63467\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_8_LC_14_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59144\,
            in2 => \_gnd_net_\,
            in3 => \N__63119\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_9_LC_14_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59148\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46525\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65549\,
            ce => \N__54112\,
            sr => \N__62906\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMMQI1_LC_14_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55221\,
            in1 => \N__55399\,
            in2 => \N__46172\,
            in3 => \N__42812\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GH5_LC_14_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__46271\,
            in1 => \N__60540\,
            in2 => \N__30852\,
            in3 => \N__30813\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIN5GHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOJAV5_LC_14_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60329\,
            in2 => \N__30849\,
            in3 => \N__30846\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13_LC_14_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41256\,
            in2 => \N__30840\,
            in3 => \N__60150\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net\,
            ce => \N__60005\,
            sr => \N__62894\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI8OT76_LC_14_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30831\,
            in1 => \N__60328\,
            in2 => \_gnd_net_\,
            in3 => \N__30837\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_4_LC_14_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__49983\,
            in1 => \_gnd_net_\,
            in2 => \N__30825\,
            in3 => \N__60151\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_13C_net\,
            ce => \N__60005\,
            sr => \N__62894\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU1492_17_LC_14_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__57935\,
            in1 => \N__58157\,
            in2 => \N__38078\,
            in3 => \N__40888\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIK8FN1_LC_14_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55183\,
            in1 => \N__55387\,
            in2 => \N__35538\,
            in3 => \N__33730\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7EQL2_LC_14_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__35537\,
            in1 => \N__54953\,
            in2 => \N__33737\,
            in3 => \N__54756\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRL7_LC_14_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53976\,
            in1 => \N__49669\,
            in2 => \N__30807\,
            in3 => \N__40791\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINCRLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI2GCO7_LC_14_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53670\,
            in2 => \N__30939\,
            in3 => \N__30936\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3_LC_14_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55584\,
            in2 => \N__30930\,
            in3 => \N__55650\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net\,
            ce => \N__55521\,
            sr => \N__62884\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICQCO7_LC_14_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__30927\,
            in1 => \N__53669\,
            in2 => \_gnd_net_\,
            in3 => \N__32139\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_5_LC_14_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30891\,
            in2 => \N__30918\,
            in3 => \N__55652\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net\,
            ce => \N__55521\,
            sr => \N__62884\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_4_LC_14_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55651\,
            in1 => \N__30915\,
            in2 => \_gnd_net_\,
            in3 => \N__30909\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_3C_net\,
            ce => \N__55521\,
            sr => \N__62884\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_9_LC_14_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38301\,
            in1 => \N__37706\,
            in2 => \N__30879\,
            in3 => \N__46671\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_9_LC_14_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33939\,
            in1 => \N__30878\,
            in2 => \N__59163\,
            in3 => \N__46461\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_21_LC_14_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__61436\,
            in1 => \N__59023\,
            in2 => \N__33365\,
            in3 => \N__33940\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_22_LC_14_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33936\,
            in1 => \N__30866\,
            in2 => \N__59160\,
            in3 => \N__61319\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_23_LC_14_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__61253\,
            in1 => \N__59024\,
            in2 => \N__37934\,
            in3 => \N__33941\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_24_LC_14_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__33937\,
            in1 => \N__61131\,
            in2 => \N__59161\,
            in3 => \N__35264\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_24,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_25_LC_14_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__35198\,
            in1 => \N__59025\,
            in2 => \N__61020\,
            in3 => \N__33942\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_25,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_26_LC_14_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__33938\,
            in1 => \N__60913\,
            in2 => \N__59162\,
            in3 => \N__30962\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.s_data_system_oZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65585\,
            ce => \N__32489\,
            sr => \N__62876\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_0_LC_14_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__62479\,
            in1 => \N__36540\,
            in2 => \_gnd_net_\,
            in3 => \N__38674\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_a2_3_LC_14_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38726\,
            in2 => \N__30948\,
            in3 => \N__64157\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.N_1959_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_0_0_tz_LC_14_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111001111"
        )
    port map (
            in0 => \N__36753\,
            in1 => \N__38699\,
            in2 => \N__30945\,
            in3 => \N__36807\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.re_elec0_tz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst2.rdata_tri_enable_LC_14_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__38821\,
            in1 => \_gnd_net_\,
            in2 => \N__30942\,
            in3 => \N__38904\,
            lcout => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst2_rdata_tri_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst0.rdata_tri_enable_LC_14_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__38903\,
            in1 => \N__38820\,
            in2 => \_gnd_net_\,
            in3 => \N__32311\,
            lcout => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst0_rdata_tri_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65597\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_2_LC_14_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__31605\,
            in1 => \N__34280\,
            in2 => \_gnd_net_\,
            in3 => \N__34148\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net\,
            ce => 'H',
            sr => \N__64970\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_8_LC_14_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__41424\,
            in1 => \N__36651\,
            in2 => \_gnd_net_\,
            in3 => \N__34421\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_2C_net\,
            ce => 'H',
            sr => \N__64970\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_o2_7_LC_14_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56246\,
            in2 => \_gnd_net_\,
            in3 => \N__38673\,
            lcout => \N_1592_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_detect_RNO_LC_14_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__39186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Control_StartUp_inst.N_8_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1EQD_LC_14_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_272_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_2_RNIUMRG2_0_LC_14_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30990\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.N_278_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_14_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19_LC_14_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000110011"
        )
    port map (
            in0 => \N__31041\,
            in1 => \N__30978\,
            in2 => \_gnd_net_\,
            in3 => \N__31263\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net\,
            ce => 'H',
            sr => \N__62857\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_RNIBV54_LC_14_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32646\,
            in2 => \_gnd_net_\,
            in3 => \N__31051\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_10_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIFSQ8_17_LC_14_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__32666\,
            in1 => \N__32696\,
            in2 => \N__30972\,
            in3 => \N__32883\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_547_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_7_LC_14_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__31262\,
            in1 => \_gnd_net_\,
            in2 => \N__31125\,
            in3 => \N__31131\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net\,
            ce => 'H',
            sr => \N__62857\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIPCFF_19_LC_14_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__31052\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31119\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.en_count_bits_0_i_a2_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIO9811_11_LC_14_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31027\,
            in1 => \N__31384\,
            in2 => \N__31101\,
            in3 => \N__31225\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_277_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_20_LC_14_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__31053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31261\,
            lcout => \cemf_module_64ch_ctrl_inst1.end_conf_a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net\,
            ce => 'H',
            sr => \N__62857\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_18_LC_14_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32667\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_19C_net\,
            ce => 'H',
            sr => \N__62857\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_RNILJCF_LC_14_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__31035\,
            in1 => \N__31218\,
            in2 => \N__31302\,
            in3 => \N__31280\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_270\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_LC_14_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_12_LC_14_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31028\,
            in2 => \_gnd_net_\,
            in3 => \N__31258\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_15_LC_14_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011101"
        )
    port map (
            in0 => \N__31259\,
            in1 => \N__31290\,
            in2 => \N__31227\,
            in3 => \N__31301\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_9_LC_14_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32271\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_14_LC_14_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__32272\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_13_LC_14_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31282\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_16_LC_14_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__31260\,
            in1 => \_gnd_net_\,
            in2 => \N__31226\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retC_net\,
            ce => 'H',
            sr => \N__62850\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIK0RN1_16_LC_14_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__31171\,
            in1 => \N__32698\,
            in2 => \N__31185\,
            in3 => \N__31139\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_LC_14_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31203\,
            in3 => \N__31191\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_retZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net\,
            ce => 'H',
            sr => \N__62846\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIIF971_13_LC_14_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__32673\,
            in1 => \N__32566\,
            in2 => \N__32276\,
            in3 => \N__32297\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_276_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_6_LC_14_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__31140\,
            in1 => \N__31184\,
            in2 => \N__32703\,
            in3 => \N__31172\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_1967\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net\,
            ce => 'H',
            sr => \N__62846\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNIEJSO_0_LC_14_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32592\,
            in2 => \_gnd_net_\,
            in3 => \N__36956\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_reti_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_LC_14_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31395\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net\,
            ce => 'H',
            sr => \N__62846\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_1_RNI7P0A1_LC_14_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__31392\,
            in1 => \N__31383\,
            in2 => \N__31365\,
            in3 => \N__32591\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.N_273\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_LC_14_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111010001000100"
        )
    port map (
            in0 => \N__36957\,
            in1 => \N__31350\,
            in2 => \N__31343\,
            in3 => \N__32904\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.c_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13C_net\,
            ce => 'H',
            sr => \N__62846\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIMH2I_LC_14_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__32950\,
            in1 => \N__37168\,
            in2 => \N__34551\,
            in3 => \N__35755\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNI6VG51_LC_14_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32782\,
            in2 => \N__31320\,
            in3 => \N__32818\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addrlde_i_0_a2_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43_0_LC_14_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__36696\,
            in1 => \N__36868\,
            in2 => \N__31317\,
            in3 => \N__39743\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIFIK43Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIS0GS_LC_14_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__39742\,
            in1 => \N__32949\,
            in2 => \_gnd_net_\,
            in3 => \N__32817\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1852_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_10_LC_14_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35796\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65657\,
            ce => 'H',
            sr => \N__62839\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_RNIIDR41_LC_14_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__35756\,
            in1 => \N__34543\,
            in2 => \N__32718\,
            in3 => \N__36695\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2\,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1946_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.next_sequence_1_c_state_ret_6_RNICL4J4_LC_14_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__36836\,
            in1 => \N__31551\,
            in2 => \N__31539\,
            in3 => \N__31536\,
            lcout => \N_528_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_2_LC_14_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31413\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_1_LC_14_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31503\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_2_LC_14_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__31488\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.sync_50hz_q_RNI5H26_2_LC_14_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31494\,
            in2 => \_gnd_net_\,
            in3 => \N__31487\,
            lcout => \cemf_module_64ch_ctrl_inst1.n_state41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__un35_li_0_i_i_a2_0_a2_1_LC_14_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__36904\,
            in1 => \N__32951\,
            in2 => \N__31457\,
            in3 => \N__34512\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_li_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_1_LC_14_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50790\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65672\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0_LC_14_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__34331\,
            in1 => \N__32540\,
            in2 => \N__63301\,
            in3 => \N__31407\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\,
            ce => 'H',
            sr => \N__64991\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_1_LC_14_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__32538\,
            in1 => \N__34332\,
            in2 => \N__63273\,
            in3 => \N__31401\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\,
            ce => 'H',
            sr => \N__64991\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_3_LC_14_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__34334\,
            in1 => \N__32541\,
            in2 => \N__63302\,
            in3 => \N__31617\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\,
            ce => 'H',
            sr => \N__64991\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_2_LC_14_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__32539\,
            in1 => \N__34333\,
            in2 => \N__63274\,
            in3 => \N__31611\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\,
            ce => 'H',
            sr => \N__64991\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIH7DQ_3_LC_14_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__34216\,
            in1 => \N__34240\,
            in2 => \_gnd_net_\,
            in3 => \N__34189\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_275_0\,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_275_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNI7FJ71_0_LC_14_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010100000"
        )
    port map (
            in0 => \N__34116\,
            in1 => \_gnd_net_\,
            in2 => \N__31596\,
            in3 => \N__34276\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_1_LC_14_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__34335\,
            in1 => \N__63231\,
            in2 => \N__31593\,
            in3 => \N__36573\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_0C_net\,
            ce => 'H',
            sr => \N__64991\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI344J1_1_LC_14_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__63230\,
            in1 => \N__34330\,
            in2 => \N__34125\,
            in3 => \N__34299\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_13_LC_14_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37116\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65696\,
            ce => 'H',
            sr => \N__62823\
        );

    \serializer_mod_inst.current_state_1_LC_14_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45174\,
            in2 => \_gnd_net_\,
            in3 => \N__45064\,
            lcout => \serializer_mod_inst.current_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65724\,
            ce => 'H',
            sr => \N__62813\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_2_LC_15_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__33087\,
            in1 => \N__31575\,
            in2 => \N__51926\,
            in3 => \N__49752\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_2_LC_15_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31569\,
            in1 => \N__52769\,
            in2 => \N__31764\,
            in3 => \N__52513\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_2_LC_15_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52204\,
            in2 => \N__31746\,
            in3 => \N__43005\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_2_LC_15_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35280\,
            in1 => \N__33297\,
            in2 => \N__31743\,
            in3 => \N__31740\,
            lcout => \I2C_top_level_inst1_s_data_oreg_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65514\,
            ce => \N__54515\,
            sr => \N__65002\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_10_LC_15_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31734\,
            in1 => \N__52674\,
            in2 => \N__31716\,
            in3 => \N__52494\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_10_LC_15_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__42738\,
            in1 => \_gnd_net_\,
            in2 => \N__31698\,
            in3 => \N__52123\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_10_LC_15_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__44640\,
            in1 => \N__31695\,
            in2 => \N__61712\,
            in3 => \N__44414\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_10_LC_15_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__31677\,
            in1 => \N__51791\,
            in2 => \N__31668\,
            in3 => \N__49307\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_10_LC_15_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__31665\,
            in1 => \N__37890\,
            in2 => \N__31653\,
            in3 => \N__31650\,
            lcout => \I2C_top_level_inst1_s_data_oreg_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65519\,
            ce => \N__54512\,
            sr => \N__64998\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_18_LC_15_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52495\,
            in1 => \N__31644\,
            in2 => \N__58766\,
            in3 => \N__44639\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_11_LC_15_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31935\,
            in1 => \N__52673\,
            in2 => \N__31914\,
            in3 => \N__52493\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_11_LC_15_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52122\,
            in2 => \N__31893\,
            in3 => \N__42915\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_11_LC_15_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__44409\,
            in1 => \N__63905\,
            in2 => \N__44660\,
            in3 => \N__31890\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_11_LC_15_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__51790\,
            in1 => \N__31872\,
            in2 => \N__31857\,
            in3 => \N__42558\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_11_LC_15_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__31854\,
            in1 => \N__31848\,
            in2 => \N__31842\,
            in3 => \N__35079\,
            lcout => \I2C_top_level_inst1_s_data_oreg_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65523\,
            ce => \N__54508\,
            sr => \N__64993\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_19_LC_15_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31839\,
            in1 => \N__44628\,
            in2 => \N__58634\,
            in3 => \N__44408\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_20_LC_15_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__31821\,
            in1 => \N__52676\,
            in2 => \N__31803\,
            in3 => \N__52381\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_20_LC_15_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52124\,
            in2 => \N__31785\,
            in3 => \N__35691\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_20_LC_15_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__31782\,
            in1 => \N__38374\,
            in2 => \N__58593\,
            in3 => \N__44664\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_20_LC_15_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__32028\,
            in1 => \N__38278\,
            in2 => \N__32013\,
            in3 => \N__42423\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_20_LC_15_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38034\,
            in1 => \N__33465\,
            in2 => \N__32010\,
            in3 => \N__32007\,
            lcout => \I2C_top_level_inst1_s_data_oreg_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65530\,
            ce => \N__54504\,
            sr => \N__64988\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQEFN1_LC_15_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__33673\,
            in1 => \N__55217\,
            in2 => \N__41088\,
            in3 => \N__55431\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIDKQL2_LC_15_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__55001\,
            in1 => \N__33674\,
            in2 => \N__54836\,
            in3 => \N__41087\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRL7_LC_15_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53949\,
            in1 => \N__31981\,
            in2 => \N__31965\,
            in3 => \N__33747\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI6SRLZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SL7_LC_15_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011101111111111"
        )
    port map (
            in0 => \N__40510\,
            in1 => \N__45513\,
            in2 => \N__53994\,
            in3 => \N__40560\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB1SLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIM4DO7_LC_15_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32058\,
            in1 => \_gnd_net_\,
            in2 => \N__31962\,
            in3 => \N__53695\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHVCO7_LC_15_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__53694\,
            in1 => \N__31953\,
            in2 => \_gnd_net_\,
            in3 => \N__31959\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6_LC_15_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__31947\,
            in1 => \_gnd_net_\,
            in2 => \N__31938\,
            in3 => \N__55693\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net\,
            ce => \N__55522\,
            sr => \N__62895\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_7_LC_15_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55694\,
            in1 => \N__32064\,
            in2 => \_gnd_net_\,
            in3 => \N__32057\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_6C_net\,
            ce => \N__55522\,
            sr => \N__62895\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_6_LC_15_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38269\,
            in1 => \N__37694\,
            in2 => \N__32040\,
            in3 => \N__41083\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_6_LC_15_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33946\,
            in1 => \N__32039\,
            in2 => \N__59544\,
            in3 => \N__63543\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_16_LC_15_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__57632\,
            in1 => \N__59333\,
            in2 => \N__34910\,
            in3 => \N__33947\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_17_LC_15_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33943\,
            in1 => \N__35330\,
            in2 => \N__59541\,
            in3 => \N__57423\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_18_LC_15_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__59850\,
            in1 => \N__59334\,
            in2 => \N__33521\,
            in3 => \N__33948\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_19_LC_15_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33944\,
            in1 => \N__35234\,
            in2 => \N__59542\,
            in3 => \N__61639\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_2_LC_15_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__61711\,
            in1 => \N__59335\,
            in2 => \N__35303\,
            in3 => \N__33949\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_20_LC_15_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111001000100"
        )
    port map (
            in0 => \N__33945\,
            in1 => \N__33479\,
            in2 => \N__59543\,
            in3 => \N__61526\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65550\,
            ce => \N__32512\,
            sr => \N__62885\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2HK93_LC_15_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__45842\,
            in1 => \N__46013\,
            in2 => \N__32208\,
            in3 => \N__42212\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRL7_LC_15_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53969\,
            in1 => \N__32170\,
            in2 => \N__32142\,
            in3 => \N__32133\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1NRLZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBIQL2_LC_15_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__54928\,
            in1 => \N__54736\,
            in2 => \N__41126\,
            in3 => \N__32110\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_5_LC_15_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63677\,
            in2 => \_gnd_net_\,
            in3 => \N__59141\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65562\,
            ce => \N__49059\,
            sr => \N__62877\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOOQI1_LC_15_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55154\,
            in1 => \N__55386\,
            in2 => \N__42644\,
            in3 => \N__32080\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_14_LC_15_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58496\,
            in2 => \_gnd_net_\,
            in3 => \N__59140\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65562\,
            ce => \N__49059\,
            sr => \N__62877\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIBU5H2_LC_15_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__54929\,
            in1 => \N__54735\,
            in2 => \N__42645\,
            in3 => \N__32081\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_7_LC_15_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000000011111111"
        )
    port map (
            in0 => \N__34092\,
            in1 => \N__50449\,
            in2 => \N__63472\,
            in3 => \N__33798\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65575\,
            ce => \N__32488\,
            sr => \N__62870\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_m2_0_LC_15_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000011111000"
        )
    port map (
            in0 => \N__36306\,
            in1 => \N__34844\,
            in2 => \N__34671\,
            in3 => \N__38665\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_i_0_LC_15_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__38706\,
            in1 => \N__34670\,
            in2 => \N__32067\,
            in3 => \N__62481\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_iZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_1_LC_15_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61863\,
            in2 => \_gnd_net_\,
            in3 => \N__34091\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65575\,
            ce => \N__32488\,
            sr => \N__62870\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa_0_a2_0_LC_15_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36272\,
            in1 => \N__34843\,
            in2 => \_gnd_net_\,
            in3 => \N__38664\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.n_data_system_o_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_15_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__38666\,
            in1 => \N__34851\,
            in2 => \_gnd_net_\,
            in3 => \N__36324\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.N_1825_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_27_LC_15_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__35177\,
            in1 => \N__59139\,
            in2 => \N__60816\,
            in3 => \N__33922\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_27,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65575\,
            ce => \N__32488\,
            sr => \N__62870\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_5_LC_15_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__33919\,
            in1 => \N__32222\,
            in2 => \N__63697\,
            in3 => \N__59016\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_10_LC_15_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__58783\,
            in1 => \N__37904\,
            in2 => \N__33950\,
            in3 => \N__59012\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_11_LC_15_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__33916\,
            in1 => \N__58660\,
            in2 => \N__35099\,
            in3 => \N__59013\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_12_LC_15_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__58596\,
            in1 => \N__59010\,
            in2 => \N__35060\,
            in3 => \N__33920\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_13_LC_15_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010011100100"
        )
    port map (
            in0 => \N__33917\,
            in1 => \N__35018\,
            in2 => \N__58357\,
            in3 => \N__59014\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_14_LC_15_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__58500\,
            in1 => \N__59011\,
            in2 => \N__34988\,
            in3 => \N__33921\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_15_LC_15_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000011011000"
        )
    port map (
            in0 => \N__33918\,
            in1 => \N__57520\,
            in2 => \N__34943\,
            in3 => \N__59015\,
            lcout => cemf_module_64ch_ctrl_inst1_s_data_system_o_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65586\,
            ce => \N__32490\,
            sr => \N__62862\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_16_LC_15_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64071\,
            in1 => \N__32451\,
            in2 => \N__43431\,
            in3 => \N__37803\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_764\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_18_LC_15_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32336\,
            in1 => \N__43370\,
            in2 => \N__32433\,
            in3 => \N__64072\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1911\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISS83_0_0_LC_15_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66799\,
            in2 => \_gnd_net_\,
            in3 => \N__57238\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1843_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_8_LC_15_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32337\,
            in1 => \N__32400\,
            in2 => \N__32385\,
            in3 => \N__64070\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1920\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst3.rdata_tri_enable_LC_15_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__38893\,
            in1 => \N__38808\,
            in2 => \_gnd_net_\,
            in3 => \N__32313\,
            lcout => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst3_rdata_tri_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.ram_module_top_inst.ram_module_inst1.rdata_tri_enable_LC_15_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__38892\,
            in1 => \N__38807\,
            in2 => \_gnd_net_\,
            in3 => \N__32312\,
            lcout => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_ram_module_top_inst_ram_module_inst1_rdata_tri_enable,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65598\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_LC_15_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__32557\,
            in1 => \N__32298\,
            in2 => \N__32277\,
            in3 => \N__32671\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net\,
            ce => 'H',
            sr => \N__62851\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_17_LC_15_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32702\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_stateZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net\,
            ce => 'H',
            sr => \N__62851\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_8_LC_15_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32672\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_i_3_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net\,
            ce => 'H',
            sr => \N__62851\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_1_LC_15_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__32602\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36967\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_12C_net\,
            ce => 'H',
            sr => \N__62851\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_RNIETUR_1_LC_15_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36477\,
            in1 => \N__36435\,
            in2 => \_gnd_net_\,
            in3 => \N__66274\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1372_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI216D_2_LC_15_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__43813\,
            in1 => \N__36595\,
            in2 => \_gnd_net_\,
            in3 => \N__34420\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1379_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI2QEM_0_LC_15_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__50881\,
            in1 => \N__43671\,
            in2 => \_gnd_net_\,
            in3 => \N__34170\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_113_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI35U51_14_LC_15_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__34147\,
            in1 => \N__34359\,
            in2 => \_gnd_net_\,
            in3 => \N__34295\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_11_0_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_14_LC_15_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010111001111"
        )
    port map (
            in0 => \N__32751\,
            in1 => \N__50865\,
            in2 => \N__34358\,
            in3 => \N__43931\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_12_LC_15_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__43902\,
            in1 => \N__48256\,
            in2 => \_gnd_net_\,
            in3 => \N__36676\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_12_LC_15_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__36638\,
            in1 => \N__63197\,
            in2 => \N__32520\,
            in3 => \N__32727\,
            lcout => \I2C_top_level_inst1.s_enable_desp_tx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net\,
            ce => 'H',
            sr => \N__64980\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_12_LC_15_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__43932\,
            in1 => \N__32750\,
            in2 => \_gnd_net_\,
            in3 => \N__34375\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_13_LC_15_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36639\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63198\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net\,
            ce => 'H',
            sr => \N__64980\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_LC_15_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110010001100"
        )
    port map (
            in0 => \N__50864\,
            in1 => \N__34354\,
            in2 => \N__43686\,
            in3 => \N__36677\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_new_addressZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net\,
            ce => 'H',
            sr => \N__64980\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_4_LC_15_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__36675\,
            in1 => \N__43903\,
            in2 => \_gnd_net_\,
            in3 => \N__48257\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1381_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_4_LC_15_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110110000"
        )
    port map (
            in0 => \N__43904\,
            in1 => \N__36640\,
            in2 => \N__32721\,
            in3 => \N__36599\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_12C_net\,
            ce => 'H',
            sr => \N__64980\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO59R_2_LC_15_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100011"
        )
    port map (
            in0 => \N__32899\,
            in1 => \N__36958\,
            in2 => \N__32862\,
            in3 => \N__35725\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_5_LC_15_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000001100000001"
        )
    port map (
            in0 => \N__32857\,
            in1 => \N__35748\,
            in2 => \N__36968\,
            in3 => \N__32903\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_392\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65631\,
            ce => 'H',
            sr => \N__62840\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_4_LC_15_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__32902\,
            in1 => \N__36960\,
            in2 => \_gnd_net_\,
            in3 => \N__32858\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_state_i_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65631\,
            ce => 'H',
            sr => \N__62840\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_3_LC_15_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32709\,
            in2 => \_gnd_net_\,
            in3 => \N__32901\,
            lcout => \cemf_module_64ch_ctrl_inst1.start_conf_b\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65631\,
            ce => 'H',
            sr => \N__62840\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_RNI2QTM_20_LC_15_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000110011"
        )
    port map (
            in0 => \N__32900\,
            in1 => \N__36959\,
            in2 => \_gnd_net_\,
            in3 => \N__32856\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.N_1817_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_2_LC_15_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__32865\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65631\,
            ce => 'H',
            sr => \N__62840\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIM2JK_2_LC_15_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35818\,
            in2 => \_gnd_net_\,
            in3 => \N__32855\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1846_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_4_LC_15_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__35819\,
            in1 => \N__35881\,
            in2 => \_gnd_net_\,
            in3 => \N__32993\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65631\,
            ce => 'H',
            sr => \N__62840\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_RNI3S391_LC_15_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100000111"
        )
    port map (
            in0 => \N__32838\,
            in1 => \N__36955\,
            in2 => \N__32826\,
            in3 => \N__37083\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1874_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNISDQ71_10_LC_15_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001110000"
        )
    port map (
            in0 => \N__36954\,
            in1 => \N__37161\,
            in2 => \N__36909\,
            in3 => \N__36717\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1873_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIP3H21_LC_15_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36837\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__32783\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_RNIAUPM2_LC_15_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__37082\,
            in1 => \N__34521\,
            in2 => \N__32799\,
            in3 => \N__32796\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1950\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_1_RNIVHBV1_LC_15_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__32790\,
            in1 => \N__32784\,
            in2 => \_gnd_net_\,
            in3 => \N__34511\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.stop_fpga2_0_0_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNIUA133_LC_15_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__39757\,
            in1 => \N__32952\,
            in2 => \N__33027\,
            in3 => \N__36900\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1949_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_RNII03U6_LC_15_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__34599\,
            in1 => \N__33024\,
            in2 => \N__33018\,
            in3 => \N__35400\,
            lcout => stop_fpga2_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_5_LC_15_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__35888\,
            in2 => \_gnd_net_\,
            in3 => \N__32997\,
            lcout => \cemf_module_64ch_ctrl_inst1.clr_sys_reg\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_1_LC_15_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34629\,
            in2 => \_gnd_net_\,
            in3 => \N__35396\,
            lcout => \cemf_module_64ch_ctrl_inst1.start_conf_a\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_7_LC_15_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__35367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35922\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1847\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \serializer_mod_inst.shift_reg_55_LC_15_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47883\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40122\,
            lcout => \serializer_mod_inst.shift_regZ0Z_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \serializer_mod_inst.shift_reg_113_LC_15_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__32931\,
            in1 => \N__45389\,
            in2 => \_gnd_net_\,
            in3 => \N__44901\,
            lcout => \serializer_mod_inst.shift_regZ0Z_113\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_0_LC_15_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34494\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \serializer_mod_inst.shift_reg_112_LC_15_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__33060\,
            in1 => \N__45388\,
            in2 => \_gnd_net_\,
            in3 => \N__44900\,
            lcout => \serializer_mod_inst.shift_regZ0Z_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65658\,
            ce => 'H',
            sr => \N__62830\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_2_LC_15_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48105\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65673\,
            ce => \N__44088\,
            sr => \N__64997\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_4_LC_15_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41376\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65673\,
            ce => \N__44088\,
            sr => \N__64997\
        );

    \serializer_mod_inst.shift_reg_111_LC_15_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47879\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34740\,
            lcout => \serializer_mod_inst.shift_regZ0Z_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65682\,
            ce => 'H',
            sr => \N__62818\
        );

    \serializer_mod_inst.shift_reg_119_LC_15_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33033\,
            in2 => \_gnd_net_\,
            in3 => \N__47880\,
            lcout => \serializer_mod_inst.shift_regZ0Z_119\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65682\,
            ce => 'H',
            sr => \N__62818\
        );

    \serializer_mod_inst.shift_reg_39_LC_15_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47882\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33183\,
            lcout => \serializer_mod_inst.shift_regZ0Z_39\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65682\,
            ce => 'H',
            sr => \N__62818\
        );

    \serializer_mod_inst.shift_reg_121_LC_15_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33045\,
            in2 => \_gnd_net_\,
            in3 => \N__47881\,
            lcout => \serializer_mod_inst.shift_regZ0Z_121\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65682\,
            ce => 'H',
            sr => \N__62818\
        );

    \serializer_mod_inst.shift_reg_120_LC_15_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__44964\,
            in1 => \N__33051\,
            in2 => \_gnd_net_\,
            in3 => \N__45247\,
            lcout => \serializer_mod_inst.shift_regZ0Z_120\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65682\,
            ce => 'H',
            sr => \N__62818\
        );

    \serializer_mod_inst.shift_reg_36_LC_15_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33165\,
            lcout => \serializer_mod_inst.shift_regZ0Z_36\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65697\,
            ce => 'H',
            sr => \N__62814\
        );

    \serializer_mod_inst.shift_reg_37_LC_15_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45031\,
            in1 => \N__33039\,
            in2 => \_gnd_net_\,
            in3 => \N__45177\,
            lcout => \serializer_mod_inst.shift_regZ0Z_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65697\,
            ce => 'H',
            sr => \N__62814\
        );

    \serializer_mod_inst.shift_reg_118_LC_15_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34863\,
            in2 => \_gnd_net_\,
            in3 => \N__47877\,
            lcout => \serializer_mod_inst.shift_regZ0Z_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65697\,
            ce => 'H',
            sr => \N__62814\
        );

    \serializer_mod_inst.shift_reg_33_LC_15_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45030\,
            in1 => \N__34563\,
            in2 => \_gnd_net_\,
            in3 => \N__45176\,
            lcout => \serializer_mod_inst.shift_regZ0Z_33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65697\,
            ce => 'H',
            sr => \N__62814\
        );

    \serializer_mod_inst.shift_reg_38_LC_15_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45178\,
            in1 => \N__33189\,
            in2 => \_gnd_net_\,
            in3 => \N__45032\,
            lcout => \serializer_mod_inst.shift_regZ0Z_38\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65697\,
            ce => 'H',
            sr => \N__62814\
        );

    \serializer_mod_inst.shift_reg_76_LC_15_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40245\,
            lcout => \serializer_mod_inst.shift_regZ0Z_76\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65715\,
            ce => 'H',
            sr => \N__62810\
        );

    \serializer_mod_inst.shift_reg_34_LC_15_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__33177\,
            in1 => \N__45175\,
            in2 => \_gnd_net_\,
            in3 => \N__45057\,
            lcout => \serializer_mod_inst.shift_regZ0Z_34\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65715\,
            ce => 'H',
            sr => \N__62810\
        );

    \serializer_mod_inst.shift_reg_35_LC_15_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33171\,
            in2 => \_gnd_net_\,
            in3 => \N__47869\,
            lcout => \serializer_mod_inst.shift_regZ0Z_35\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65715\,
            ce => 'H',
            sr => \N__62810\
        );

    \serializer_mod_inst.shift_reg_77_LC_15_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33159\,
            in2 => \_gnd_net_\,
            in3 => \N__47871\,
            lcout => \serializer_mod_inst.shift_regZ0Z_77\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65715\,
            ce => 'H',
            sr => \N__62810\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_17_LC_16_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64246\,
            in1 => \N__33153\,
            in2 => \N__43572\,
            in3 => \N__37878\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_753\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_19_LC_16_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37879\,
            in1 => \N__43529\,
            in2 => \N__33123\,
            in3 => \N__64249\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_731\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_2_LC_16_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64248\,
            in1 => \N__33102\,
            in2 => \N__43574\,
            in3 => \N__37877\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_918\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_22_LC_16_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37874\,
            in1 => \N__43519\,
            in2 => \N__33345\,
            in3 => \N__64245\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_698\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_23_LC_16_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64247\,
            in1 => \N__33312\,
            in2 => \N__43573\,
            in3 => \N__37880\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_687\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_2_LC_16_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__52983\,
            in1 => \N__53792\,
            in2 => \N__53318\,
            in3 => \N__49965\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_25_LC_16_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64243\,
            in1 => \N__33291\,
            in2 => \N__43571\,
            in3 => \N__37875\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_665\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_27_LC_16_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37876\,
            in1 => \N__43518\,
            in2 => \N__33273\,
            in3 => \N__64244\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_654\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_19_LC_16_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__33255\,
            in1 => \N__52672\,
            in2 => \N__33237\,
            in3 => \N__52440\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_19_LC_16_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__33216\,
            in1 => \N__33210\,
            in2 => \N__51867\,
            in3 => \N__51510\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_19_LC_16_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35217\,
            in1 => \N__33438\,
            in2 => \N__33204\,
            in3 => \N__33195\,
            lcout => \I2C_top_level_inst1_s_data_oreg_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65513\,
            ce => \N__54509\,
            sr => \N__65003\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_19_LC_16_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__52145\,
            in1 => \N__33201\,
            in2 => \_gnd_net_\,
            in3 => \N__48681\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_19_LC_16_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52982\,
            in1 => \N__57330\,
            in2 => \N__53324\,
            in3 => \N__51477\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_1_LC_16_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__56606\,
            in1 => \N__47415\,
            in2 => \N__47307\,
            in3 => \N__42888\,
            lcout => \s_paddr_I2C_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65517\,
            ce => \N__50091\,
            sr => \N__64999\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_2_LC_16_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47414\,
            in1 => \N__56607\,
            in2 => \N__47271\,
            in3 => \N__42870\,
            lcout => \s_paddr_I2C_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65517\,
            ce => \N__50091\,
            sr => \N__64999\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_1_0_LC_16_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__35989\,
            in1 => \N__36268\,
            in2 => \N__43514\,
            in3 => \N__64172\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_214_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_0_LC_16_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__64174\,
            in1 => \N__43436\,
            in2 => \N__36273\,
            in3 => \N__35988\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_213_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIRQ9DD_0_LC_16_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__43435\,
            in1 => \N__33431\,
            in2 => \_gnd_net_\,
            in3 => \N__64173\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1319_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_0_LC_16_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__33408\,
            in1 => \N__33393\,
            in2 => \N__33375\,
            in3 => \N__52441\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_0_LC_16_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52054\,
            in2 => \N__33372\,
            in3 => \N__48921\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_21_LC_16_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__52903\,
            in1 => \N__37642\,
            in2 => \N__33369\,
            in3 => \N__46317\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_1_LC_16_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37641\,
            in1 => \N__52901\,
            in2 => \N__34641\,
            in3 => \N__60710\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIH49MI_2_LC_16_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__64235\,
            in1 => \N__35987\,
            in2 => \N__43581\,
            in3 => \N__36305\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_216_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_18_LC_16_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__33525\,
            in1 => \N__52902\,
            in2 => \N__33501\,
            in3 => \N__51368\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_20_LC_16_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__52904\,
            in1 => \N__37643\,
            in2 => \N__33486\,
            in3 => \N__40986\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_4_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_0_LC_16_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__35986\,
            in1 => \N__36362\,
            in2 => \N__43582\,
            in3 => \N__64236\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1876_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_7_LC_16_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__45534\,
            in1 => \N__33825\,
            in2 => \N__33459\,
            in3 => \N__37640\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15_LC_16_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60158\,
            in1 => \_gnd_net_\,
            in2 => \N__33600\,
            in3 => \N__33635\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net\,
            ce => \N__60004\,
            sr => \N__62881\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI26492_17_LC_16_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__53375\,
            in1 => \N__58190\,
            in2 => \N__48585\,
            in3 => \N__58005\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGH5_LC_16_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__60565\,
            in1 => \N__42396\,
            in2 => \N__33441\,
            in3 => \N__46211\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI1GGHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI2UAV5_LC_16_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__33636\,
            in1 => \_gnd_net_\,
            in2 => \N__33639\,
            in3 => \N__60381\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITOAV5_LC_16_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__33627\,
            in1 => \N__60380\,
            in2 => \_gnd_net_\,
            in3 => \N__33579\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_14_LC_16_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33621\,
            in2 => \N__33603\,
            in3 => \N__60157\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_15C_net\,
            ce => \N__60004\,
            sr => \N__62881\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI04492_17_LC_16_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__58004\,
            in1 => \N__38479\,
            in2 => \N__58198\,
            in3 => \N__53420\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGH5_LC_16_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60558\,
            in1 => \N__33557\,
            in2 => \N__33591\,
            in3 => \N__33588\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISAGHZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2TV43_LC_16_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__45990\,
            in1 => \N__45832\,
            in2 => \N__38480\,
            in3 => \N__33556\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8D7_LC_16_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__53419\,
            in1 => \N__53978\,
            in2 => \N__33573\,
            in3 => \N__33570\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHI8DZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_14_LC_16_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58497\,
            in2 => \_gnd_net_\,
            in3 => \N__59382\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65536\,
            ce => \N__58869\,
            sr => \N__62873\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI2V153_LC_16_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__45991\,
            in1 => \N__48964\,
            in2 => \N__45868\,
            in3 => \N__49003\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDD7_LC_16_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__53979\,
            in1 => \N__42777\,
            in2 => \N__33792\,
            in3 => \N__51251\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIHNDDZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISQUF7_LC_16_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__36141\,
            in1 => \_gnd_net_\,
            in2 => \N__33789\,
            in3 => \N__53691\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_23_LC_16_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61247\,
            in2 => \_gnd_net_\,
            in3 => \N__59383\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65536\,
            ce => \N__58869\,
            sr => \N__62873\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4JK93_LC_16_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__45831\,
            in1 => \N__45989\,
            in2 => \N__42176\,
            in3 => \N__33775\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_1_LC_16_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61867\,
            in2 => \_gnd_net_\,
            in3 => \N__59188\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_3_LC_16_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59185\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63939\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_4_LC_16_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63809\,
            in2 => \_gnd_net_\,
            in3 => \N__59190\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_6_LC_16_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59186\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63580\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_26_LC_16_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60921\,
            in2 => \_gnd_net_\,
            in3 => \N__59189\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_0Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_20_LC_16_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59183\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61525\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_12_LC_16_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58589\,
            in2 => \_gnd_net_\,
            in3 => \N__59187\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_30_LC_16_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59184\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62184\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65546\,
            ce => \N__49033\,
            sr => \N__62865\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_15_LC_16_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011000000"
        )
    port map (
            in0 => \N__64312\,
            in1 => \N__55927\,
            in2 => \N__50625\,
            in3 => \N__64081\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1654_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_15_LC_16_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50592\,
            in2 => \N__34011\,
            in3 => \N__49875\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65556\,
            ce => 'H',
            sr => \N__64975\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNI6TP01_7_LC_16_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__63448\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59164\,
            lcout => \N_12_0\,
            ltout => \N_12_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_mem_7_LC_16_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__34008\,
            in3 => \N__64073\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pwdata_memZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_o2_LC_16_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__36294\,
            in1 => \N__36785\,
            in2 => \_gnd_net_\,
            in3 => \N__34852\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_539_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.c_data_system_o_RNO_0_7_LC_16_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101001111110011"
        )
    port map (
            in0 => \N__36396\,
            in1 => \N__33821\,
            in2 => \N__33807\,
            in3 => \N__33804\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_5_LC_16_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__50558\,
            in1 => \N__56308\,
            in2 => \_gnd_net_\,
            in3 => \N__38657\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.n_data_system_o_0_a3_2_7_LC_16_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__59165\,
            in1 => \N__34856\,
            in2 => \N__36789\,
            in3 => \N__36295\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_1786_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_26_LC_16_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001011"
        )
    port map (
            in0 => \N__34083\,
            in1 => \N__34074\,
            in2 => \N__66813\,
            in3 => \N__64074\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_4093_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.N_536_i_i_o2_LC_16_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100010"
        )
    port map (
            in0 => \N__46807\,
            in1 => \N__64117\,
            in2 => \N__39660\,
            in3 => \N__39145\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1868_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISBI9D_0_LC_16_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010000000"
        )
    port map (
            in0 => \N__43366\,
            in1 => \N__37804\,
            in2 => \N__64209\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_LC_16_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__47111\,
            in1 => \N__34062\,
            in2 => \_gnd_net_\,
            in3 => \N__39144\,
            lcout => \N_409\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_o2_0_a2_2_LC_16_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__47172\,
            in1 => \N__54334\,
            in2 => \N__56151\,
            in3 => \N__41609\,
            lcout => cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2,
            ltout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_pready_i_o2_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIAC0UC_7_LC_16_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__47110\,
            in1 => \N__50244\,
            in2 => \N__34056\,
            in3 => \N__39143\,
            lcout => \N_1838_0\,
            ltout => \N_1838_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ91HD_0_LC_16_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__43365\,
            in1 => \_gnd_net_\,
            in2 => \N__34053\,
            in3 => \N__34049\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE6LS1_15_LC_16_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43235\,
            in1 => \N__43268\,
            in2 => \N__43205\,
            in3 => \N__43034\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_2043_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_12_LC_16_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__64574\,
            in1 => \N__47411\,
            in2 => \N__41487\,
            in3 => \N__43023\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65582\,
            ce => \N__50087\,
            sr => \N__64976\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_13_LC_16_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47409\,
            in1 => \N__64576\,
            in2 => \N__41469\,
            in3 => \N__43257\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65582\,
            ce => \N__50087\,
            sr => \N__64976\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_14_LC_16_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__64575\,
            in1 => \N__47412\,
            in2 => \N__41454\,
            in3 => \N__43224\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65582\,
            ce => \N__50087\,
            sr => \N__64976\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_15_LC_16_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47410\,
            in1 => \N__64577\,
            in2 => \N__41439\,
            in3 => \N__43185\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65582\,
            ce => \N__50087\,
            sr => \N__64976\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_0_LC_16_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__57685\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.s_data_ireg_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => \N__36503\,
            sr => \N__62843\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_1_LC_16_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48262\,
            lcout => \I2C_top_level_inst1.s_data_ireg_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => \N__36503\,
            sr => \N__62843\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_7_LC_16_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41733\,
            lcout => \I2C_top_level_inst1.s_data_ireg_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => \N__36503\,
            sr => \N__62843\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_5_LC_16_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41375\,
            lcout => \I2C_top_level_inst1.s_data_ireg_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => \N__36503\,
            sr => \N__62843\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_2_LC_16_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48140\,
            lcout => \I2C_top_level_inst1.s_data_ireg_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => \N__36503\,
            sr => \N__62843\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_4_LC_16_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48032\,
            lcout => \I2C_top_level_inst1.s_data_ireg_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47983\,
            ce => \N__36503\,
            sr => \N__62843\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIEDSM_1_LC_16_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111111"
        )
    port map (
            in0 => \N__34167\,
            in1 => \N__34449\,
            in2 => \N__34149\,
            in3 => \N__34313\,
            lcout => \I2C_top_level_inst1.N_327_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_6_LC_16_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__50874\,
            in1 => \N__36634\,
            in2 => \_gnd_net_\,
            in3 => \N__34168\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1400_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_6_LC_16_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__36657\,
            in1 => \N__34404\,
            in2 => \N__34302\,
            in3 => \N__34381\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net\,
            ce => 'H',
            sr => \N__64984\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNILBK01_6_LC_16_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101110101011"
        )
    port map (
            in0 => \N__50873\,
            in1 => \N__34166\,
            in2 => \N__34458\,
            in3 => \N__41574\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1374_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_bit_counter_RNIAT631_3_LC_16_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__34281\,
            in1 => \N__34248\,
            in2 => \N__34224\,
            in3 => \N__34197\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0\,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1354_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_7_LC_16_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__50872\,
            in1 => \_gnd_net_\,
            in2 => \N__34173\,
            in3 => \N__34169\,
            lcout => \I2C_top_level_inst1.s_load_addr1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net\,
            ce => 'H',
            sr => \N__64984\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_11_LC_16_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011000000000000"
        )
    port map (
            in0 => \N__41576\,
            in1 => \N__50871\,
            in2 => \N__36647\,
            in3 => \N__34454\,
            lcout => \I2C_top_level_inst1.s_load_wdata\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_6C_net\,
            ce => 'H',
            sr => \N__64984\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_1_LC_16_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010011111100"
        )
    port map (
            in0 => \N__34453\,
            in1 => \N__34146\,
            in2 => \N__50885\,
            in3 => \N__41575\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_2_10_LC_16_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__34455\,
            in1 => \N__41521\,
            in2 => \N__43733\,
            in3 => \N__66275\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1399_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_10_LC_16_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001011"
        )
    port map (
            in0 => \N__43720\,
            in1 => \N__50884\,
            in2 => \N__34473\,
            in3 => \N__41577\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIIMIE_11_LC_16_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__50883\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50979\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0\,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1373_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_10_LC_16_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000001"
        )
    port map (
            in0 => \N__43721\,
            in1 => \N__34456\,
            in2 => \N__34470\,
            in3 => \N__34382\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1395_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_10_LC_16_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__34457\,
            in1 => \N__36643\,
            in2 => \N__34467\,
            in3 => \N__34464\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net\,
            ce => 'H',
            sr => \N__64989\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_9_LC_16_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__36642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34428\,
            lcout => \I2C_top_level_inst1.s_load_addr0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net\,
            ce => 'H',
            sr => \N__64989\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_14_LC_16_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__34403\,
            in1 => \N__41522\,
            in2 => \_gnd_net_\,
            in3 => \N__66276\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1409_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_14_LC_16_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110111110101"
        )
    port map (
            in0 => \N__34392\,
            in1 => \N__43938\,
            in2 => \N__34386\,
            in3 => \N__34383\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_state_10C_net\,
            ce => 'H',
            sr => \N__64989\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_2_LC_16_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37149\,
            in1 => \N__37108\,
            in2 => \N__34557\,
            in3 => \N__36735\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_14_LC_16_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34556\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_381_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65626\,
            ce => 'H',
            sr => \N__62828\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_8_LC_16_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__34555\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36736\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1880\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65626\,
            ce => 'H',
            sr => \N__62828\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_10_LC_16_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37032\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_71_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65626\,
            ce => 'H',
            sr => \N__62828\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI6HM8_10_LC_16_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36734\,
            in2 => \_gnd_net_\,
            in3 => \N__36714\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_1848_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.N_1848_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIVI6G_15_LC_16_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37148\,
            in2 => \N__34515\,
            in3 => \N__35724\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1884_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_15_LC_16_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36737\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65626\,
            ce => 'H',
            sr => \N__62828\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_11_LC_16_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__36715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65626\,
            ce => 'H',
            sr => \N__62828\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI2MBM1_5_LC_16_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__34654\,
            in1 => \N__35394\,
            in2 => \N__34639\,
            in3 => \N__34597\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_520_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_0_LC_16_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37031\,
            in2 => \N__34488\,
            in3 => \N__37064\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_0_a2_6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_LC_16_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1101010111111111"
        )
    port map (
            in0 => \N__35795\,
            in1 => \N__34485\,
            in2 => \N__34476\,
            in3 => \N__34701\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65642\,
            ce => 'H',
            sr => \N__62822\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNO_1_LC_16_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__35360\,
            in1 => \N__35915\,
            in2 => \N__34710\,
            in3 => \N__37019\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un41_i_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_12_RNIDMPS1_LC_16_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34695\,
            in1 => \N__34680\,
            in2 => \_gnd_net_\,
            in3 => \N__34689\,
            lcout => \c_state_ret_12_RNIDMPS1_0\,
            ltout => \c_state_ret_12_RNIDMPS1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.current_state_0_LC_16_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001000010000"
        )
    port map (
            in0 => \N__45469\,
            in1 => \N__44899\,
            in2 => \N__34674\,
            in3 => \N__45498\,
            lcout => \serializer_mod_inst.current_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65642\,
            ce => 'H',
            sr => \N__62822\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_LC_16_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000001010001"
        )
    port map (
            in0 => \N__34655\,
            in1 => \N__35395\,
            in2 => \N__34640\,
            in3 => \N__34598\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_i_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65642\,
            ce => 'H',
            sr => \N__62822\
        );

    \serializer_mod_inst.shift_reg_7_LC_16_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101101000001010"
        )
    port map (
            in0 => \N__44894\,
            in1 => \_gnd_net_\,
            in2 => \N__45464\,
            in3 => \N__41847\,
            lcout => \serializer_mod_inst.shift_regZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65653\,
            ce => 'H',
            sr => \N__62817\
        );

    \serializer_mod_inst.shift_reg_11_LC_16_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37239\,
            in1 => \N__45422\,
            in2 => \_gnd_net_\,
            in3 => \N__44895\,
            lcout => \serializer_mod_inst.shift_regZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65653\,
            ce => 'H',
            sr => \N__62817\
        );

    \serializer_mod_inst.shift_reg_8_LC_16_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__34575\,
            in1 => \N__45426\,
            in2 => \_gnd_net_\,
            in3 => \N__44896\,
            lcout => \serializer_mod_inst.shift_regZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65653\,
            ce => 'H',
            sr => \N__62817\
        );

    \serializer_mod_inst.shift_reg_31_LC_16_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__44214\,
            in1 => \N__45411\,
            in2 => \_gnd_net_\,
            in3 => \N__45033\,
            lcout => \serializer_mod_inst.shift_regZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65668\,
            ce => 'H',
            sr => \N__62812\
        );

    \serializer_mod_inst.shift_reg_32_LC_16_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44949\,
            in2 => \N__45462\,
            in3 => \N__34569\,
            lcout => \serializer_mod_inst.shift_regZ0Z_32\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65668\,
            ce => 'H',
            sr => \N__62812\
        );

    \serializer_mod_inst.shift_reg_48_LC_16_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37347\,
            in1 => \N__45415\,
            in2 => \_gnd_net_\,
            in3 => \N__45034\,
            lcout => \serializer_mod_inst.shift_regZ0Z_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65668\,
            ce => 'H',
            sr => \N__62812\
        );

    \serializer_mod_inst.shift_reg_115_LC_16_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34746\,
            in2 => \_gnd_net_\,
            in3 => \N__47876\,
            lcout => \serializer_mod_inst.shift_regZ0Z_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65668\,
            ce => 'H',
            sr => \N__62812\
        );

    \serializer_mod_inst.shift_reg_114_LC_16_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34755\,
            in2 => \_gnd_net_\,
            in3 => \N__47875\,
            lcout => \serializer_mod_inst.shift_regZ0Z_114\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65668\,
            ce => 'H',
            sr => \N__62812\
        );

    \serializer_mod_inst.shift_reg_79_LC_16_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45027\,
            in1 => \N__34722\,
            in2 => \_gnd_net_\,
            in3 => \N__45406\,
            lcout => \serializer_mod_inst.shift_regZ0Z_79\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65680\,
            ce => 'H',
            sr => \N__62809\
        );

    \serializer_mod_inst.shift_reg_110_LC_16_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45403\,
            in1 => \N__41922\,
            in2 => \_gnd_net_\,
            in3 => \N__45028\,
            lcout => \serializer_mod_inst.shift_regZ0Z_110\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65680\,
            ce => 'H',
            sr => \N__62809\
        );

    \serializer_mod_inst.shift_reg_40_LC_16_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45026\,
            in1 => \N__34734\,
            in2 => \_gnd_net_\,
            in3 => \N__45404\,
            lcout => \serializer_mod_inst.shift_regZ0Z_40\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65680\,
            ce => 'H',
            sr => \N__62809\
        );

    \serializer_mod_inst.shift_reg_78_LC_16_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45405\,
            in1 => \N__34728\,
            in2 => \_gnd_net_\,
            in3 => \N__45029\,
            lcout => \serializer_mod_inst.shift_regZ0Z_78\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65680\,
            ce => 'H',
            sr => \N__62809\
        );

    \serializer_mod_inst.shift_reg_41_LC_16_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34716\,
            in2 => \_gnd_net_\,
            in3 => \N__47874\,
            lcout => \serializer_mod_inst.shift_regZ0Z_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65680\,
            ce => 'H',
            sr => \N__62809\
        );

    \serializer_mod_inst.shift_reg_67_LC_16_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45058\,
            in2 => \N__45357\,
            in3 => \N__40176\,
            lcout => \serializer_mod_inst.shift_regZ0Z_67\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65692\,
            ce => 'H',
            sr => \N__62806\
        );

    \serializer_mod_inst.shift_reg_69_LC_16_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45059\,
            in2 => \N__45358\,
            in3 => \N__34884\,
            lcout => \serializer_mod_inst.shift_regZ0Z_69\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65692\,
            ce => 'H',
            sr => \N__62806\
        );

    \serializer_mod_inst.shift_reg_68_LC_16_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47812\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__34890\,
            lcout => \serializer_mod_inst.shift_regZ0Z_68\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65692\,
            ce => 'H',
            sr => \N__62806\
        );

    \serializer_mod_inst.shift_reg_116_LC_16_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__34878\,
            in1 => \N__47811\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \serializer_mod_inst.shift_regZ0Z_116\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65692\,
            ce => 'H',
            sr => \N__62806\
        );

    \serializer_mod_inst.shift_reg_117_LC_16_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__34869\,
            in1 => \N__45232\,
            in2 => \_gnd_net_\,
            in3 => \N__45060\,
            lcout => \serializer_mod_inst.shift_regZ0Z_117\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65692\,
            ce => 'H',
            sr => \N__62806\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa_0_a2_0_LC_16_27_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__38679\,
            in1 => \N__36366\,
            in2 => \_gnd_net_\,
            in3 => \N__34857\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.n_data_system_o_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \rst_n_ibuf_RNIBNDC_LC_16_32_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35464\,
            lcout => rst_n_c_i,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_12_LC_17_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__52146\,
            in1 => \N__41234\,
            in2 => \N__53317\,
            in3 => \N__40961\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_12_LC_17_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__34800\,
            in1 => \N__52675\,
            in2 => \N__34779\,
            in3 => \N__52484\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_12_LC_17_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53000\,
            in2 => \N__34758\,
            in3 => \N__46350\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_12_LC_17_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__35154\,
            in1 => \N__44661\,
            in2 => \N__63831\,
            in3 => \N__44427\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_12_LC_17_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__35136\,
            in1 => \N__51824\,
            in2 => \N__35124\,
            in3 => \N__41202\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_12_LC_17_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__35037\,
            in1 => \N__35121\,
            in2 => \N__35115\,
            in3 => \N__35112\,
            lcout => \I2C_top_level_inst1_s_data_oreg_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65520\,
            ce => \N__54505\,
            sr => \N__65005\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_11_LC_17_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38220\,
            in1 => \N__37649\,
            in2 => \N__35106\,
            in3 => \N__42951\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_12_LC_17_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37650\,
            in1 => \N__38221\,
            in2 => \N__35070\,
            in3 => \N__42705\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_13_LC_17_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38216\,
            in1 => \N__37645\,
            in2 => \N__35031\,
            in3 => \N__42813\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_14_LC_17_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37644\,
            in1 => \N__38215\,
            in2 => \N__34992\,
            in3 => \N__42643\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_15_LC_17_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38218\,
            in1 => \N__37648\,
            in2 => \N__34953\,
            in3 => \N__42612\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_16_LC_17_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37647\,
            in1 => \N__38219\,
            in2 => \N__34914\,
            in3 => \N__42582\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_17_LC_17_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38217\,
            in1 => \N__37646\,
            in2 => \N__35340\,
            in3 => \N__45617\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_3_0_LC_17_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__36355\,
            in1 => \N__35996\,
            in2 => \N__43583\,
            in3 => \N__64234\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_215_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_2_LC_17_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__37656\,
            in1 => \N__35304\,
            in2 => \N__35283\,
            in3 => \N__42975\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_24_LC_17_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__38238\,
            in1 => \N__35268\,
            in2 => \N__35250\,
            in3 => \N__37657\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_24_LC_17_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__61103\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59388\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65531\,
            ce => \N__45570\,
            sr => \N__62907\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_19_LC_17_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38237\,
            in1 => \N__37655\,
            in2 => \N__35241\,
            in3 => \N__48705\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_25_LC_17_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__37658\,
            in1 => \N__38239\,
            in2 => \N__44238\,
            in3 => \N__35205\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_27_LC_17_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__35184\,
            in1 => \N__38214\,
            in2 => \N__35163\,
            in3 => \N__37654\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_27_LC_17_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60797\,
            in2 => \_gnd_net_\,
            in3 => \N__59384\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65541\,
            ce => \N__45568\,
            sr => \N__62896\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_28_LC_17_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__35655\,
            in1 => \N__38213\,
            in2 => \N__35619\,
            in3 => \N__37653\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_28_LC_17_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62336\,
            in2 => \_gnd_net_\,
            in3 => \N__59385\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65541\,
            ce => \N__45568\,
            sr => \N__62896\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_29_LC_17_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__35610\,
            in1 => \N__38211\,
            in2 => \N__35589\,
            in3 => \N__37652\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_29_LC_17_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__62264\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59386\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65541\,
            ce => \N__45568\,
            sr => \N__62896\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_3_LC_17_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__35580\,
            in1 => \N__37651\,
            in2 => \N__35533\,
            in3 => \N__38212\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_3_LC_17_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63923\,
            in2 => \_gnd_net_\,
            in3 => \N__59387\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65541\,
            ce => \N__45568\,
            sr => \N__62896\
        );

    \serializer_mod_inst.serial_out_test_e_0_LC_17_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__44007\,
            in1 => \N__45485\,
            in2 => \_gnd_net_\,
            in3 => \N__45090\,
            lcout => serial_out_testing_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65551\,
            ce => \N__35481\,
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIIO3I_0_LC_17_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40096\,
            in2 => \_gnd_net_\,
            in3 => \N__39791\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1965\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIOU3I_6_LC_17_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__40097\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40002\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_522_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_2_RNIMEFF_LC_17_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40041\,
            in2 => \_gnd_net_\,
            in3 => \N__40098\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_525_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIO4JK_4_LC_17_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__35892\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35862\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1845_reti_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNIP1G7_15_LC_17_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37169\,
            in2 => \_gnd_net_\,
            in3 => \N__35761\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_1854_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIGUF7_LC_17_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__36183\,
            in1 => \N__53692\,
            in2 => \_gnd_net_\,
            in3 => \N__45708\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINLUF7_LC_17_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__53693\,
            in1 => \N__38403\,
            in2 => \_gnd_net_\,
            in3 => \N__36159\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIKSI1_LC_17_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__55155\,
            in1 => \N__42412\,
            in2 => \N__55451\,
            in3 => \N__35680\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5Q7H2_LC_17_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__35681\,
            in1 => \N__55010\,
            in2 => \N__42419\,
            in3 => \N__54802\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DD7_LC_17_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53977\,
            in1 => \N__38566\,
            in2 => \N__35667\,
            in3 => \N__40800\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI28DDZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIDBUF7_LC_17_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53671\,
            in1 => \_gnd_net_\,
            in2 => \N__35664\,
            in3 => \N__35661\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20_LC_17_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49191\,
            in2 => \N__36192\,
            in3 => \N__55686\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net\,
            ce => \N__55563\,
            sr => \N__62878\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_21_LC_17_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55687\,
            in1 => \N__36189\,
            in2 => \_gnd_net_\,
            in3 => \N__36182\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net\,
            ce => \N__55563\,
            sr => \N__62878\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_22_LC_17_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__36171\,
            in1 => \N__55688\,
            in2 => \_gnd_net_\,
            in3 => \N__36158\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net\,
            ce => \N__55563\,
            sr => \N__62878\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_23_LC_17_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__55689\,
            in1 => \N__36147\,
            in2 => \_gnd_net_\,
            in3 => \N__36140\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.dout_conf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_20C_net\,
            ce => \N__55563\,
            sr => \N__62878\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIH49MI_2_0_LC_17_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__35990\,
            in1 => \N__36317\,
            in2 => \N__43569\,
            in3 => \N__64066\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1875_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.addr_mem_0_a2_i_1_LC_17_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__64067\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__35991\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1831_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__36259\,
            in1 => \N__38656\,
            in2 => \N__35997\,
            in3 => \N__64068\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.N_1824_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPOSB_11_LC_17_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56868\,
            in2 => \_gnd_net_\,
            in3 => \N__57718\,
            lcout => \N_1841_0\,
            ltout => \N_1841_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_LC_17_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__35992\,
            in1 => \N__36354\,
            in2 => \N__35925\,
            in3 => \N__64069\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.N_112_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_12_LC_17_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66184\,
            in2 => \_gnd_net_\,
            in3 => \N__57719\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65576\,
            ce => 'H',
            sr => \N__64981\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_11_LC_17_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111000001000000"
        )
    port map (
            in0 => \N__50943\,
            in1 => \N__50559\,
            in2 => \N__50490\,
            in3 => \N__47517\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65576\,
            ce => 'H',
            sr => \N__64981\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_13_LC_17_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011101100"
        )
    port map (
            in0 => \N__43173\,
            in1 => \N__56869\,
            in2 => \N__56245\,
            in3 => \N__66185\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65576\,
            ce => 'H',
            sr => \N__64981\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNINHAS1_0_LC_17_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39036\,
            in1 => \N__46764\,
            in2 => \_gnd_net_\,
            in3 => \N__39113\,
            lcout => \N_1613\,
            ltout => \N_1613_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001100"
        )
    port map (
            in0 => \N__39612\,
            in1 => \N__46900\,
            in2 => \N__36369\,
            in3 => \N__39132\,
            lcout => \N_1860_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000001010"
        )
    port map (
            in0 => \N__36219\,
            in1 => \N__39611\,
            in2 => \N__46910\,
            in3 => \N__39116\,
            lcout => \N_202_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII7LO3_2_LC_17_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__39114\,
            in1 => \N__46896\,
            in2 => \N__39617\,
            in3 => \N__36218\,
            lcout => \N_1859_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.n_data_system_o_1_sqmuxa_0_a2_0_i_o2_LC_17_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010100000"
        )
    port map (
            in0 => \N__36220\,
            in1 => \N__39613\,
            in2 => \N__46909\,
            in3 => \N__39115\,
            lcout => \N_1861_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.prdata_1_4_u_i_m2_0_LC_17_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__48519\,
            in1 => \N__45588\,
            in2 => \_gnd_net_\,
            in3 => \N__36221\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_id.N_604\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI7T453_9_LC_17_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__47043\,
            in1 => \N__47013\,
            in2 => \N__46950\,
            in3 => \N__47456\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_404_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIE7FP3_4_LC_17_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47243\,
            in2 => \N__36417\,
            in3 => \N__47206\,
            lcout => \N_396\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_6_0_a3_0_o2_LC_17_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__36402\,
            in1 => \N__36408\,
            in2 => \N__36384\,
            in3 => \N__36414\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_399_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_4_LC_17_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41377\,
            lcout => \I2C_top_level_inst1.s_command_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__47921\,
            sr => \N__62858\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_5_LC_17_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41796\,
            lcout => \I2C_top_level_inst1.s_command_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__47921\,
            sr => \N__62858\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_6_LC_17_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41734\,
            lcout => \I2C_top_level_inst1.s_command_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__47921\,
            sr => \N__62858\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIFO5I1_7_LC_17_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39455\,
            in2 => \_gnd_net_\,
            in3 => \N__39109\,
            lcout => \N_1803\,
            ltout => \N_1803_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_26_LC_17_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37182\,
            in1 => \N__36519\,
            in2 => \N__36387\,
            in3 => \N__36375\,
            lcout => \N_410\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_7_LC_17_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41688\,
            lcout => \I2C_top_level_inst1.s_command_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47978\,
            ce => \N__47921\,
            sr => \N__62858\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6_26_LC_17_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39512\,
            in1 => \N__39536\,
            in2 => \N__39486\,
            in3 => \N__39566\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_6Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_a2_6_0_LC_17_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__41729\,
            in1 => \N__41786\,
            in2 => \N__41658\,
            in3 => \N__41348\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_300_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_6_LC_17_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41787\,
            lcout => \I2C_top_level_inst1.s_data_ireg_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47980\,
            ce => \N__36510\,
            sr => \N__62852\
        );

    \I2C_top_level_inst1.RX_Shift_Register_inst.data_o_3_LC_17_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.s_data_ireg_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47980\,
            ce => \N__36510\,
            sr => \N__62852\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_a2_1_0_LC_17_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__48020\,
            in1 => \N__48132\,
            in2 => \_gnd_net_\,
            in3 => \N__48080\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1425_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0_LC_17_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100001000100"
        )
    port map (
            in0 => \N__36486\,
            in1 => \N__36449\,
            in2 => \_gnd_net_\,
            in3 => \N__36472\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            ce => 'H',
            sr => \N__64990\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNIUAQ1_11_LC_17_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50983\,
            in2 => \_gnd_net_\,
            in3 => \N__43954\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0\,
            ltout => \I2C_top_level_inst1.I2C_FSM_inst.N_1367_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_1_LC_17_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100011000000000"
        )
    port map (
            in0 => \N__36473\,
            in1 => \N__36431\,
            in2 => \N__36453\,
            in3 => \N__36450\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_byte_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            ce => 'H',
            sr => \N__64990\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_r_w_LC_17_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010000000100"
        )
    port map (
            in0 => \N__43664\,
            in1 => \N__51299\,
            in2 => \N__43901\,
            in3 => \N__48258\,
            lcout => \I2C_top_level_inst1.s_r_w\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            ce => 'H',
            sr => \N__64990\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_0_LC_17_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000110100001111"
        )
    port map (
            in0 => \N__43790\,
            in1 => \N__43665\,
            in2 => \N__43638\,
            in3 => \N__43852\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            ce => 'H',
            sr => \N__64990\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_3_LC_17_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__43853\,
            in1 => \N__43828\,
            in2 => \_gnd_net_\,
            in3 => \N__43789\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            ce => 'H',
            sr => \N__64990\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_6_LC_17_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__36678\,
            in1 => \N__47914\,
            in2 => \_gnd_net_\,
            in3 => \N__43887\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_5_LC_17_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36641\,
            in2 => \_gnd_net_\,
            in3 => \N__36600\,
            lcout => \I2C_top_level_inst1.s_load_command\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.I2C_FSM_inst.c_byte_counter_0C_net\,
            ce => 'H',
            sr => \N__64990\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_1_LC_17_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__36579\,
            in1 => \N__36561\,
            in2 => \N__43748\,
            in3 => \N__43956\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_1_1_LC_17_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__47912\,
            in1 => \N__41406\,
            in2 => \_gnd_net_\,
            in3 => \N__43885\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.c_state_ns_i_i_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNI8SIH_3_LC_17_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__43886\,
            in1 => \N__47913\,
            in2 => \N__43749\,
            in3 => \N__41413\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.N_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.s_sda_o_tx_RNITO2M_LC_17_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__63292\,
            in1 => \N__36981\,
            in2 => \N__36555\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.N_259\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_552_i_0_a2_LC_17_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__36530\,
            in1 => \N__62456\,
            in2 => \_gnd_net_\,
            in3 => \N__56878\,
            lcout => \N_552_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7_26_LC_17_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39878\,
            in1 => \N__39893\,
            in2 => \N__39711\,
            in3 => \N__39908\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_7Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.s_sda_o_q_1_LC_17_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36975\,
            lcout => \I2C_top_level_inst1.s_sda_o_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.s_sda_o_tx_LC_17_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__36987\,
            lcout => \I2C_top_level_inst1.s_sda_o_txZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65632\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.s_sda_o_q_0_LC_17_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61989\,
            lcout => \I2C_top_level_inst1.s_sda_o_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_RNI8HA01_1_LC_17_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36969\,
            in2 => \_gnd_net_\,
            in3 => \N__36908\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_1855_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.N_1855_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_RNI6LR22_LC_17_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37005\,
            in2 => \N__36846\,
            in3 => \N__36838\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_1857_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.N_1857_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.prdata15_0_o3_0_a2_LC_17_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111100000000"
        )
    port map (
            in0 => \N__36770\,
            in1 => \N__36689\,
            in2 => \N__36792\,
            in3 => \N__39146\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.N_384\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.n_data_system_o_1_sqmuxa_0_a2_2_o2_0_LC_17_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__36771\,
            in1 => \N__37048\,
            in2 => \_gnd_net_\,
            in3 => \N__37107\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.N_1840_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_RNI1ITL_8_LC_17_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__37106\,
            in1 => \N__36738\,
            in2 => \N__37050\,
            in3 => \N__36716\,
            lcout => \cemf_module_64ch_ctrl_inst1.N_383\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8_26_LC_17_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__39848\,
            in1 => \N__39863\,
            in2 => \N__39834\,
            in3 => \N__39421\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_0_i_o2_0_a3_8Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_12_LC_17_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__37160\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_state_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65659\,
            ce => 'H',
            sr => \N__62831\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_ret_9_LC_17_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37159\,
            in2 => \_gnd_net_\,
            in3 => \N__37109\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.N_1862\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65659\,
            ce => 'H',
            sr => \N__62831\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_8_LC_17_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37068\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_state_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65659\,
            ce => 'H',
            sr => \N__62831\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_9_LC_17_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37049\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65659\,
            ce => 'H',
            sr => \N__62831\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.un35_4_0__c_state_ret_6_LC_17_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37020\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_retZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65659\,
            ce => 'H',
            sr => \N__62831\
        );

    \serializer_mod_inst.shift_reg_1_LC_17_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__44898\,
            in1 => \N__45427\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \serializer_mod_inst.shift_regZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65674\,
            ce => 'H',
            sr => \N__62824\
        );

    \serializer_mod_inst.shift_reg_12_LC_17_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__36999\,
            in2 => \_gnd_net_\,
            in3 => \N__47857\,
            lcout => \serializer_mod_inst.shift_regZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65674\,
            ce => 'H',
            sr => \N__62824\
        );

    \serializer_mod_inst.shift_reg_49_LC_17_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__36993\,
            in1 => \N__45428\,
            in2 => \_gnd_net_\,
            in3 => \N__44902\,
            lcout => \serializer_mod_inst.shift_regZ0Z_49\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65674\,
            ce => 'H',
            sr => \N__62824\
        );

    \serializer_mod_inst.shift_reg_91_LC_17_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44897\,
            in2 => \N__45465\,
            in3 => \N__39915\,
            lcout => \serializer_mod_inst.shift_regZ0Z_91\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65674\,
            ce => 'H',
            sr => \N__62824\
        );

    \serializer_mod_inst.shift_reg_51_LC_17_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__47858\,
            in1 => \_gnd_net_\,
            in2 => \N__39930\,
            in3 => \_gnd_net_\,
            lcout => \serializer_mod_inst.shift_regZ0Z_51\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65674\,
            ce => 'H',
            sr => \N__62824\
        );

    \serializer_mod_inst.shift_reg_52_LC_17_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47859\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37245\,
            lcout => \serializer_mod_inst.shift_regZ0Z_52\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65674\,
            ce => 'H',
            sr => \N__62824\
        );

    \serializer_mod_inst.shift_reg_10_LC_17_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37188\,
            in1 => \N__45416\,
            in2 => \_gnd_net_\,
            in3 => \N__45083\,
            lcout => \serializer_mod_inst.shift_regZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_56_LC_17_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44948\,
            in2 => \N__45463\,
            in3 => \N__37233\,
            lcout => \serializer_mod_inst.shift_regZ0Z_56\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_15_LC_17_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37212\,
            in1 => \N__45418\,
            in2 => \_gnd_net_\,
            in3 => \N__45085\,
            lcout => \serializer_mod_inst.shift_regZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_122_LC_17_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37221\,
            in2 => \_gnd_net_\,
            in3 => \N__47851\,
            lcout => \serializer_mod_inst.shift_regZ0Z_122\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_14_LC_17_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37200\,
            in1 => \N__45417\,
            in2 => \_gnd_net_\,
            in3 => \N__45084\,
            lcout => \serializer_mod_inst.shift_regZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_13_LC_17_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__37206\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__47852\,
            lcout => \serializer_mod_inst.shift_regZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_9_LC_17_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37194\,
            in2 => \_gnd_net_\,
            in3 => \N__47853\,
            lcout => \serializer_mod_inst.shift_regZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65683\,
            ce => 'H',
            sr => \N__62819\
        );

    \serializer_mod_inst.shift_reg_18_LC_17_25_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47850\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37269\,
            lcout => \serializer_mod_inst.shift_regZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65698\,
            ce => 'H',
            sr => \N__62815\
        );

    \serializer_mod_inst.shift_reg_16_LC_17_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45066\,
            in1 => \N__37287\,
            in2 => \_gnd_net_\,
            in3 => \N__45407\,
            lcout => \serializer_mod_inst.shift_regZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65698\,
            ce => 'H',
            sr => \N__62815\
        );

    \serializer_mod_inst.shift_reg_80_LC_17_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45410\,
            in1 => \N__37281\,
            in2 => \_gnd_net_\,
            in3 => \N__45069\,
            lcout => \serializer_mod_inst.shift_regZ0Z_80\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65698\,
            ce => 'H',
            sr => \N__62815\
        );

    \serializer_mod_inst.shift_reg_108_LC_17_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37257\,
            in2 => \_gnd_net_\,
            in3 => \N__47849\,
            lcout => \serializer_mod_inst.shift_regZ0Z_108\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65698\,
            ce => 'H',
            sr => \N__62815\
        );

    \serializer_mod_inst.shift_reg_17_LC_17_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45408\,
            in1 => \N__37275\,
            in2 => \_gnd_net_\,
            in3 => \N__45068\,
            lcout => \serializer_mod_inst.shift_regZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65698\,
            ce => 'H',
            sr => \N__62815\
        );

    \serializer_mod_inst.shift_reg_19_LC_17_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45067\,
            in1 => \N__37263\,
            in2 => \_gnd_net_\,
            in3 => \N__45409\,
            lcout => \serializer_mod_inst.shift_regZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65698\,
            ce => 'H',
            sr => \N__62815\
        );

    \serializer_mod_inst.shift_reg_107_LC_17_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37353\,
            in2 => \_gnd_net_\,
            in3 => \N__47810\,
            lcout => \serializer_mod_inst.shift_regZ0Z_107\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65716\,
            ce => 'H',
            sr => \N__62811\
        );

    \serializer_mod_inst.shift_reg_70_LC_17_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45076\,
            in1 => \N__37251\,
            in2 => \_gnd_net_\,
            in3 => \N__45241\,
            lcout => \serializer_mod_inst.shift_regZ0Z_70\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65716\,
            ce => 'H',
            sr => \N__62811\
        );

    \serializer_mod_inst.shift_reg_104_LC_17_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000010101010"
        )
    port map (
            in0 => \N__45074\,
            in1 => \_gnd_net_\,
            in2 => \N__40158\,
            in3 => \N__45239\,
            lcout => \serializer_mod_inst.shift_regZ0Z_104\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65716\,
            ce => 'H',
            sr => \N__62811\
        );

    \serializer_mod_inst.shift_reg_106_LC_17_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000010101010"
        )
    port map (
            in0 => \N__45075\,
            in1 => \_gnd_net_\,
            in2 => \N__37323\,
            in3 => \N__45240\,
            lcout => \serializer_mod_inst.shift_regZ0Z_106\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65716\,
            ce => 'H',
            sr => \N__62811\
        );

    \serializer_mod_inst.shift_reg_47_LC_17_27_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47864\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37314\,
            lcout => \serializer_mod_inst.shift_regZ0Z_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65725\,
            ce => 'H',
            sr => \N__62807\
        );

    \serializer_mod_inst.shift_reg_95_LC_17_27_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45047\,
            in1 => \N__37335\,
            in2 => \_gnd_net_\,
            in3 => \N__45360\,
            lcout => \serializer_mod_inst.shift_regZ0Z_95\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65725\,
            ce => 'H',
            sr => \N__62807\
        );

    \serializer_mod_inst.shift_reg_94_LC_17_27_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47865\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37293\,
            lcout => \serializer_mod_inst.shift_regZ0Z_94\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65725\,
            ce => 'H',
            sr => \N__62807\
        );

    \serializer_mod_inst.shift_reg_105_LC_17_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37329\,
            in2 => \_gnd_net_\,
            in3 => \N__47863\,
            lcout => \serializer_mod_inst.shift_regZ0Z_105\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65725\,
            ce => 'H',
            sr => \N__62807\
        );

    \serializer_mod_inst.shift_reg_46_LC_17_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40272\,
            in1 => \N__45359\,
            in2 => \_gnd_net_\,
            in3 => \N__45048\,
            lcout => \serializer_mod_inst.shift_regZ0Z_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65725\,
            ce => 'H',
            sr => \N__62807\
        );

    \serializer_mod_inst.shift_reg_97_LC_17_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37461\,
            in1 => \N__45442\,
            in2 => \_gnd_net_\,
            in3 => \N__45053\,
            lcout => \serializer_mod_inst.shift_regZ0Z_97\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65736\,
            ce => 'H',
            sr => \N__62805\
        );

    \serializer_mod_inst.shift_reg_92_LC_17_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37308\,
            in2 => \_gnd_net_\,
            in3 => \N__47867\,
            lcout => \serializer_mod_inst.shift_regZ0Z_92\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65736\,
            ce => 'H',
            sr => \N__62805\
        );

    \serializer_mod_inst.shift_reg_93_LC_17_28_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47868\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__37299\,
            lcout => \serializer_mod_inst.shift_regZ0Z_93\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65736\,
            ce => 'H',
            sr => \N__62805\
        );

    \serializer_mod_inst.shift_reg_96_LC_17_28_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__37467\,
            in1 => \N__45441\,
            in2 => \_gnd_net_\,
            in3 => \N__45052\,
            lcout => \serializer_mod_inst.shift_regZ0Z_96\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65736\,
            ce => 'H',
            sr => \N__62805\
        );

    \serializer_mod_inst.shift_reg_98_LC_17_29_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45049\,
            in1 => \N__37455\,
            in2 => \_gnd_net_\,
            in3 => \N__45445\,
            lcout => \serializer_mod_inst.shift_regZ0Z_98\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65745\,
            ce => 'H',
            sr => \N__62804\
        );

    \serializer_mod_inst.enable_config_LC_17_29_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45443\,
            in2 => \_gnd_net_\,
            in3 => \N__45051\,
            lcout => enable_config_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65745\,
            ce => 'H',
            sr => \N__62804\
        );

    \serializer_mod_inst.serial_out_LC_17_29_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__45050\,
            in1 => \N__44003\,
            in2 => \_gnd_net_\,
            in3 => \N__45444\,
            lcout => elec_config_out_c,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65745\,
            ce => 'H',
            sr => \N__62804\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_24_LC_18_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__37713\,
            in1 => \N__51891\,
            in2 => \N__48537\,
            in3 => \N__42291\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_24_LC_18_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__37422\,
            in1 => \N__37407\,
            in2 => \N__37410\,
            in3 => \N__37359\,
            lcout => \I2C_top_level_inst1_s_data_oreg_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65521\,
            ce => \N__54506\,
            sr => \N__65016\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_24_LC_18_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__54222\,
            in1 => \N__53286\,
            in2 => \N__40437\,
            in3 => \N__52989\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_24_LC_18_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__37401\,
            in1 => \N__52756\,
            in2 => \N__37383\,
            in3 => \N__52512\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_24_LC_18_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__46578\,
            in1 => \_gnd_net_\,
            in2 => \N__37362\,
            in3 => \N__52199\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_23_LC_18_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__37700\,
            in1 => \N__38311\,
            in2 => \N__37938\,
            in3 => \N__49497\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_10_LC_18_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__37914\,
            in1 => \N__37699\,
            in2 => \N__38318\,
            in3 => \N__42765\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_6_24_LC_18_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__37843\,
            in1 => \N__43584\,
            in2 => \N__37731\,
            in3 => \N__64250\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_676\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_0_LC_18_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__40113\,
            in1 => \N__37698\,
            in2 => \N__38317\,
            in3 => \N__48942\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_23_LC_18_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__51846\,
            in1 => \N__37557\,
            in2 => \N__37548\,
            in3 => \N__49004\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_23_LC_18_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__37524\,
            in1 => \N__37533\,
            in2 => \N__37527\,
            in3 => \N__37473\,
            lcout => \I2C_top_level_inst1_s_data_oreg_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65532\,
            ce => \N__54498\,
            sr => \N__65006\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_23_LC_18_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52988\,
            in1 => \N__48974\,
            in2 => \N__53306\,
            in3 => \N__51252\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_23_LC_18_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__37518\,
            in1 => \N__52738\,
            in2 => \N__37497\,
            in3 => \N__52496\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_23_LC_18_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001110000"
        )
    port map (
            in0 => \N__49464\,
            in1 => \N__52191\,
            in2 => \N__37476\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_20_LC_18_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__53194\,
            in1 => \N__42447\,
            in2 => \N__51915\,
            in3 => \N__38576\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_2_21_LC_18_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__45744\,
            in1 => \N__53195\,
            in2 => \N__45768\,
            in3 => \N__51871\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_5_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQV592_17_LC_18_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__58165\,
            in1 => \N__58015\,
            in2 => \N__38577\,
            in3 => \N__42446\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJJFV5_LC_18_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60353\,
            in1 => \N__38025\,
            in2 => \_gnd_net_\,
            in3 => \N__46086\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21_LC_18_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__37986\,
            in2 => \N__38019\,
            in3 => \N__60187\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net\,
            ce => \N__60009\,
            sr => \N__62915\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LH5_LC_18_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60604\,
            in1 => \N__40985\,
            in2 => \N__38016\,
            in3 => \N__38007\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNID0LHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIEEFV5_LC_18_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60358\,
            in1 => \_gnd_net_\,
            in2 => \N__37998\,
            in3 => \N__37995\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_20_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_20_LC_18_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60186\,
            in1 => \_gnd_net_\,
            in2 => \N__37989\,
            in3 => \N__51525\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_21C_net\,
            ce => \N__60009\,
            sr => \N__62915\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_21_LC_18_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__37980\,
            in1 => \N__52755\,
            in2 => \N__37959\,
            in3 => \N__52446\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_1_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_21_LC_18_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52198\,
            in2 => \N__38397\,
            in3 => \N__45678\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_3_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_21_LC_18_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__38394\,
            in1 => \N__58350\,
            in2 => \N__44647\,
            in3 => \N__38375\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_21_LC_18_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__38328\,
            in1 => \N__38222\,
            in2 => \N__38127\,
            in3 => \N__45699\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_6_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_21_LC_18_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__38124\,
            in1 => \N__38118\,
            in2 => \N__38106\,
            in3 => \N__38103\,
            lcout => \I2C_top_level_inst1_s_data_oreg_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65552\,
            ce => \N__54496\,
            sr => \N__65000\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_12_LC_18_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58595\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_21_LC_18_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59633\,
            in2 => \_gnd_net_\,
            in3 => \N__61406\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_30_LC_18_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59638\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62165\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_13_LC_18_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59632\,
            in2 => \_gnd_net_\,
            in3 => \N__58351\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_22_LC_18_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59639\,
            in1 => \N__61352\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_31_LC_18_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59635\,
            in2 => \_gnd_net_\,
            in3 => \N__62070\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_14_LC_18_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59637\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58498\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_23_LC_18_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59634\,
            in2 => \_gnd_net_\,
            in3 => \N__61193\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65564\,
            ce => \N__48723\,
            sr => \N__62897\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIMOSI1_LC_18_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55163\,
            in1 => \N__55423\,
            in2 => \N__42674\,
            in3 => \N__38596\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALH5_LC_18_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60557\,
            in1 => \N__42277\,
            in2 => \N__38445\,
            in3 => \N__38442\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNINALHZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIU3692_17_LC_18_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__57914\,
            in1 => \N__58120\,
            in2 => \N__38429\,
            in3 => \N__38518\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_22_LC_18_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61353\,
            in2 => \_gnd_net_\,
            in3 => \N__59553\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65577\,
            ce => \N__49034\,
            sr => \N__62886\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI0T153_LC_18_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__42278\,
            in1 => \N__46050\,
            in2 => \N__45915\,
            in3 => \N__38425\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDD7_LC_18_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__38519\,
            in1 => \N__54005\,
            in2 => \N__38406\,
            in3 => \N__38583\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICIDDZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9U7H2_LC_18_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__54798\,
            in1 => \N__42670\,
            in2 => \N__55035\,
            in3 => \N__38597\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_10_LC_18_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59647\,
            in2 => \_gnd_net_\,
            in3 => \N__58787\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_11_LC_18_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59643\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58692\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_20_LC_18_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__61530\,
            in1 => \N__59650\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_12_LC_18_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59644\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58594\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_21_LC_18_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59649\,
            in2 => \_gnd_net_\,
            in3 => \N__61421\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_30_LC_18_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59646\,
            in1 => \N__62179\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_13_LC_18_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59648\,
            in2 => \_gnd_net_\,
            in3 => \N__58349\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_22_LC_18_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59645\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61354\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65587\,
            ce => \N__54114\,
            sr => \N__62879\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_26_LC_18_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__56407\,
            in1 => \N__47546\,
            in2 => \N__66192\,
            in3 => \N__56593\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65599\,
            ce => 'H',
            sr => \N__64977\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBDJD_23_LC_18_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__57242\,
            in1 => \N__56406\,
            in2 => \_gnd_net_\,
            in3 => \N__56733\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_8_0_m2_ns_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI3S672_1_LC_18_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101000111"
        )
    port map (
            in0 => \N__48329\,
            in1 => \N__56592\,
            in2 => \N__38709\,
            in3 => \N__50145\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_5_LC_18_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011011100"
        )
    port map (
            in0 => \N__47547\,
            in1 => \N__56949\,
            in2 => \N__43142\,
            in3 => \N__66191\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65599\,
            ce => 'H',
            sr => \N__64977\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_6_LC_18_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__66187\,
            in1 => \N__47545\,
            in2 => \_gnd_net_\,
            in3 => \N__43135\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65599\,
            ce => 'H',
            sr => \N__64977\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_21_LC_18_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66186\,
            in2 => \_gnd_net_\,
            in3 => \N__56916\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65599\,
            ce => 'H',
            sr => \N__64977\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf_cmf.un1_n_data_system_o17_i_0_0_o2_0_LC_18_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__56915\,
            in1 => \N__43134\,
            in2 => \N__43612\,
            in3 => \N__56948\,
            lcout => \N_1842_0\,
            ltout => \N_1842_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.psel_1_N_680_i_i_a2_LC_18_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__65945\,
            in1 => \N__56828\,
            in2 => \N__38682\,
            in3 => \N__38637\,
            lcout => \N_1975\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9_LC_18_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__63045\,
            in1 => \N__63246\,
            in2 => \_gnd_net_\,
            in3 => \N__46524\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_9C_net\,
            ce => \N__63029\,
            sr => \N__62863\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI1SAS1_5_LC_18_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39513\,
            in1 => \N__47246\,
            in2 => \_gnd_net_\,
            in3 => \N__39106\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_addr_RNI1SAS1_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI3UAS1_6_LC_18_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39485\,
            in1 => \N__47164\,
            in2 => \_gnd_net_\,
            in3 => \N__39107\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_addr_RNI3UAS1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNI50BS1_7_LC_18_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__39108\,
            in1 => \N__47093\,
            in2 => \_gnd_net_\,
            in3 => \N__39456\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_addr_RNI50BS1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_RNIVPAS1_4_LC_18_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__47196\,
            in1 => \N__39537\,
            in2 => \_gnd_net_\,
            in3 => \N__39105\,
            lcout => \cemf_module_64ch_ctrl_inst1.c_addr_RNIVPAS1_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_LC_18_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39042\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_18_18_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_LUT4_0_LC_18_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39282\,
            in2 => \N__39011\,
            in3 => \N__38976\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_LUT4_0_LC_18_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__38960\,
            in2 => \N__39315\,
            in3 => \N__38931\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPT1_LC_18_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39286\,
            in2 => \N__38928\,
            in3 => \N__38835\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2_c_RNI3RPTZ0Z1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQT1_LC_18_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39253\,
            in2 => \N__38832\,
            in3 => \N__38742\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3_c_RNI6VQTZ0Z1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_3\,
            carryout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93ST1_LC_18_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101000110101"
        )
    port map (
            in0 => \N__56147\,
            in1 => \N__39426\,
            in2 => \N__39147\,
            in3 => \N__38739\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_4_c_RNI93STZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rst_LC_18_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__39281\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Control_StartUp_inst.stop_resetter_rstZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47984\,
            ce => 'H',
            sr => \N__39174\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNIJHC9_1_LC_18_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55968\,
            in2 => \_gnd_net_\,
            in3 => \N__56352\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_1_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_3_LC_18_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110011"
        )
    port map (
            in0 => \N__41385\,
            in1 => \N__47433\,
            in2 => \N__39153\,
            in3 => \N__64570\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_3_LC_18_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__54289\,
            in1 => \N__47384\,
            in2 => \N__39150\,
            in3 => \N__42852\,
            lcout => \s_paddr_I2C_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65633\,
            ce => \N__50080\,
            sr => \N__64994\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNO_LC_18_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__39564\,
            in1 => \N__54288\,
            in2 => \_gnd_net_\,
            in3 => \N__39133\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.un3_addr_mem_cry_0_c_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_5_LC_18_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__64571\,
            in1 => \N__47382\,
            in2 => \N__41766\,
            in3 => \N__43116\,
            lcout => \s_paddr_I2C_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65633\,
            ce => \N__50080\,
            sr => \N__64994\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_6_LC_18_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47381\,
            in1 => \N__64573\,
            in2 => \N__41703\,
            in3 => \N__43101\,
            lcout => \s_paddr_I2C_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65633\,
            ce => \N__50080\,
            sr => \N__64994\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_7_LC_18_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011001110000000"
        )
    port map (
            in0 => \N__64572\,
            in1 => \N__47383\,
            in2 => \N__41628\,
            in3 => \N__43086\,
            lcout => \s_paddr_I2C_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65633\,
            ce => \N__50080\,
            sr => \N__64994\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_0_LC_18_20_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39813\,
            in1 => \N__39032\,
            in2 => \_gnd_net_\,
            in3 => \N__39018\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsm_0\,
            ltout => OPEN,
            carryin => \bfn_18_20_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_1_LC_18_20_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39809\,
            in1 => \N__39646\,
            in2 => \_gnd_net_\,
            in3 => \N__39624\,
            lcout => \cemf_module_64ch_ctrl_inst1.paddr_fsm_1\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_0\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_2_LC_18_20_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39814\,
            in1 => \N__39595\,
            in2 => \_gnd_net_\,
            in3 => \N__39579\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_2,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_1\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_3_LC_18_20_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101111101110"
        )
    port map (
            in0 => \N__39810\,
            in1 => \N__39565\,
            in2 => \_gnd_net_\,
            in3 => \N__39540\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_3,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_2\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_4_LC_18_20_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39815\,
            in1 => \N__39535\,
            in2 => \_gnd_net_\,
            in3 => \N__39516\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_4,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_3\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_5_LC_18_20_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39811\,
            in1 => \N__39505\,
            in2 => \_gnd_net_\,
            in3 => \N__39489\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_5,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_4\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_6_LC_18_20_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39816\,
            in1 => \N__39475\,
            in2 => \_gnd_net_\,
            in3 => \N__39459\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_6,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_5\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_7_LC_18_20_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39812\,
            in1 => \N__39448\,
            in2 => \_gnd_net_\,
            in3 => \N__39429\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.paddr_fsmZ0Z_7\,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_6\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_7\,
            clk => \N__65649\,
            ce => \N__39696\,
            sr => \N__62847\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_8_LC_18_21_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39799\,
            in1 => \N__39425\,
            in2 => \_gnd_net_\,
            in3 => \N__39405\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_8,
            ltout => OPEN,
            carryin => \bfn_18_21_0_\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_9_LC_18_21_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39794\,
            in1 => \N__39909\,
            in2 => \_gnd_net_\,
            in3 => \N__39897\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_9,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_8\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_10_LC_18_21_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39796\,
            in1 => \N__39894\,
            in2 => \_gnd_net_\,
            in3 => \N__39882\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_10,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_9\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_11_LC_18_21_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39792\,
            in1 => \N__39879\,
            in2 => \_gnd_net_\,
            in3 => \N__39867\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_11,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_10\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_12_LC_18_21_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39797\,
            in1 => \N__39864\,
            in2 => \_gnd_net_\,
            in3 => \N__39852\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_12,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_11\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_13_LC_18_21_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39793\,
            in1 => \N__39849\,
            in2 => \_gnd_net_\,
            in3 => \N__39837\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_13,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_12\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_14_LC_18_21_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39798\,
            in1 => \N__39833\,
            in2 => \_gnd_net_\,
            in3 => \N__39819\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_14,
            ltout => OPEN,
            carryin => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_13\,
            carryout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_cry_14\,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_addr_15_LC_18_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__39795\,
            in1 => \N__39710\,
            in2 => \_gnd_net_\,
            in3 => \N__39714\,
            lcout => cemf_module_64ch_ctrl_inst1_paddr_fsm_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65660\,
            ce => \N__39695\,
            sr => \N__62841\
        );

    \serializer_mod_inst.shift_reg_86_LC_18_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__47873\,
            in1 => \N__40197\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \serializer_mod_inst.shift_regZ0Z_86\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65675\,
            ce => 'H',
            sr => \N__62835\
        );

    \serializer_mod_inst.shift_reg_87_LC_18_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__44929\,
            in1 => \N__39666\,
            in2 => \_gnd_net_\,
            in3 => \N__45459\,
            lcout => \serializer_mod_inst.shift_regZ0Z_87\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65675\,
            ce => 'H',
            sr => \N__62835\
        );

    \serializer_mod_inst.shift_reg_54_LC_18_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39957\,
            in2 => \_gnd_net_\,
            in3 => \N__47872\,
            lcout => \serializer_mod_inst.shift_regZ0Z_54\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65675\,
            ce => 'H',
            sr => \N__62835\
        );

    \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_state_0_6_LC_18_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__40112\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40033\,
            lcout => \cemf_module_64ch_ctrl_inst1.cemf_module_64ch_fsm_int1.c_stateZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65675\,
            ce => 'H',
            sr => \N__62835\
        );

    \serializer_mod_inst.shift_reg_53_LC_18_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110100000"
        )
    port map (
            in0 => \N__45458\,
            in1 => \_gnd_net_\,
            in2 => \N__39966\,
            in3 => \N__44930\,
            lcout => \serializer_mod_inst.shift_regZ0Z_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65675\,
            ce => 'H',
            sr => \N__62835\
        );

    \serializer_mod_inst.shift_reg_88_LC_18_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45065\,
            in2 => \N__39951\,
            in3 => \N__45391\,
            lcout => \serializer_mod_inst.shift_regZ0Z_88\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65684\,
            ce => 'H',
            sr => \N__62832\
        );

    \serializer_mod_inst.shift_reg_101_LC_18_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40131\,
            in1 => \N__45390\,
            in2 => \_gnd_net_\,
            in3 => \N__45082\,
            lcout => \serializer_mod_inst.shift_regZ0Z_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65684\,
            ce => 'H',
            sr => \N__62832\
        );

    \serializer_mod_inst.shift_reg_89_LC_18_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39942\,
            in2 => \_gnd_net_\,
            in3 => \N__47855\,
            lcout => \serializer_mod_inst.shift_regZ0Z_89\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65684\,
            ce => 'H',
            sr => \N__62832\
        );

    \serializer_mod_inst.shift_reg_50_LC_18_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__39936\,
            in2 => \_gnd_net_\,
            in3 => \N__47854\,
            lcout => \serializer_mod_inst.shift_regZ0Z_50\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65684\,
            ce => 'H',
            sr => \N__62832\
        );

    \serializer_mod_inst.shift_reg_90_LC_18_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47856\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__39921\,
            lcout => \serializer_mod_inst.shift_regZ0Z_90\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65684\,
            ce => 'H',
            sr => \N__62832\
        );

    \serializer_mod_inst.shift_reg_85_LC_18_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45071\,
            in1 => \N__40146\,
            in2 => \_gnd_net_\,
            in3 => \N__45451\,
            lcout => \serializer_mod_inst.shift_regZ0Z_85\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65699\,
            ce => 'H',
            sr => \N__62825\
        );

    \serializer_mod_inst.shift_reg_2_LC_18_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45070\,
            in1 => \N__40188\,
            in2 => \_gnd_net_\,
            in3 => \N__45449\,
            lcout => \serializer_mod_inst.shift_regZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65699\,
            ce => 'H',
            sr => \N__62825\
        );

    \serializer_mod_inst.shift_reg_102_LC_18_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45448\,
            in1 => \N__40182\,
            in2 => \_gnd_net_\,
            in3 => \N__45072\,
            lcout => \serializer_mod_inst.shift_regZ0Z_102\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65699\,
            ce => 'H',
            sr => \N__62825\
        );

    \serializer_mod_inst.shift_reg_66_LC_18_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45450\,
            in1 => \N__44019\,
            in2 => \_gnd_net_\,
            in3 => \N__45073\,
            lcout => \serializer_mod_inst.shift_regZ0Z_66\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65699\,
            ce => 'H',
            sr => \N__62825\
        );

    \serializer_mod_inst.shift_reg_103_LC_18_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40164\,
            in2 => \_gnd_net_\,
            in3 => \N__47848\,
            lcout => \serializer_mod_inst.shift_regZ0Z_103\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65699\,
            ce => 'H',
            sr => \N__62825\
        );

    \serializer_mod_inst.shift_reg_44_LC_18_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40284\,
            in2 => \_gnd_net_\,
            in3 => \N__47845\,
            lcout => \serializer_mod_inst.shift_regZ0Z_44\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_84_LC_18_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__47847\,
            in1 => \_gnd_net_\,
            in2 => \N__40206\,
            in3 => \_gnd_net_\,
            lcout => \serializer_mod_inst.shift_regZ0Z_84\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_22_LC_18_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41814\,
            in2 => \_gnd_net_\,
            in3 => \N__47843\,
            lcout => \serializer_mod_inst.shift_regZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_42_LC_18_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40140\,
            in1 => \N__45447\,
            in2 => \_gnd_net_\,
            in3 => \N__45086\,
            lcout => \serializer_mod_inst.shift_regZ0Z_42\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_100_LC_18_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40227\,
            in2 => \_gnd_net_\,
            in3 => \N__47842\,
            lcout => \serializer_mod_inst.shift_regZ0Z_100\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_43_LC_18_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47844\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40290\,
            lcout => \serializer_mod_inst.shift_regZ0Z_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_45_LC_18_25_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40278\,
            in2 => \_gnd_net_\,
            in3 => \N__47846\,
            lcout => \serializer_mod_inst.shift_regZ0Z_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65717\,
            ce => 'H',
            sr => \N__62820\
        );

    \serializer_mod_inst.shift_reg_72_LC_18_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45077\,
            in1 => \N__40257\,
            in2 => \_gnd_net_\,
            in3 => \N__45245\,
            lcout => \serializer_mod_inst.shift_regZ0Z_72\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_71_LC_18_26_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40263\,
            in1 => \N__45242\,
            in2 => \_gnd_net_\,
            in3 => \N__45079\,
            lcout => \serializer_mod_inst.shift_regZ0Z_71\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_74_LC_18_26_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45078\,
            in1 => \N__40212\,
            in2 => \_gnd_net_\,
            in3 => \N__45246\,
            lcout => \serializer_mod_inst.shift_regZ0Z_74\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_75_LC_18_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40251\,
            in1 => \N__45243\,
            in2 => \_gnd_net_\,
            in3 => \N__45080\,
            lcout => \serializer_mod_inst.shift_regZ0Z_75\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_99_LC_18_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__40236\,
            lcout => \serializer_mod_inst.shift_regZ0Z_99\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_73_LC_18_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47741\,
            in2 => \_gnd_net_\,
            in3 => \N__40218\,
            lcout => \serializer_mod_inst.shift_regZ0Z_73\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_83_LC_18_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40422\,
            in1 => \N__45244\,
            in2 => \_gnd_net_\,
            in3 => \N__45081\,
            lcout => \serializer_mod_inst.shift_regZ0Z_83\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65726\,
            ce => 'H',
            sr => \N__62816\
        );

    \serializer_mod_inst.shift_reg_82_LC_18_28_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40401\,
            in2 => \_gnd_net_\,
            in3 => \N__47866\,
            lcout => \serializer_mod_inst.shift_regZ0Z_82\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65746\,
            ce => 'H',
            sr => \N__62808\
        );

    \serializer_mod_inst.shift_reg_81_LC_18_28_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__40413\,
            in1 => \N__45457\,
            in2 => \_gnd_net_\,
            in3 => \N__45089\,
            lcout => \serializer_mod_inst.shift_regZ0Z_81\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65746\,
            ce => 'H',
            sr => \N__62808\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_27_LC_19_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__53008\,
            in1 => \N__51279\,
            in2 => \N__40584\,
            in3 => \N__53282\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_29_LC_19_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__51264\,
            in1 => \N__53296\,
            in2 => \N__59748\,
            in3 => \N__52999\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_29_LC_19_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__40395\,
            in1 => \N__52770\,
            in2 => \N__40374\,
            in3 => \N__52485\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_29_LC_19_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49110\,
            in2 => \N__40353\,
            in3 => \N__52214\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_29_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_29_LC_19_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__40350\,
            in1 => \N__40335\,
            in2 => \N__40329\,
            in3 => \N__40296\,
            lcout => \I2C_top_level_inst1_s_data_oreg_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65533\,
            ce => \N__54499\,
            sr => \N__65017\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_29_LC_19_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__40326\,
            in1 => \N__51890\,
            in2 => \N__48774\,
            in3 => \N__40311\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI4TB92_17_LC_19_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58016\,
            in1 => \N__58185\,
            in2 => \N__40530\,
            in3 => \N__48749\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6VB92_17_LC_19_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58186\,
            in1 => \N__58017\,
            in2 => \N__40773\,
            in3 => \N__40696\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3Q5_LC_19_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60591\,
            in1 => \N__40717\,
            in2 => \N__40491\,
            in3 => \N__40782\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIRU3QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNISCU76_LC_19_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60357\,
            in2 => \N__40488\,
            in3 => \N__40485\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8_LC_19_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60203\,
            in1 => \_gnd_net_\,
            in2 => \N__40479\,
            in3 => \N__40443\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net\,
            ce => \N__59994\,
            sr => \N__62933\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3Q5_LC_19_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60517\,
            in1 => \N__45529\,
            in2 => \N__40476\,
            in3 => \N__40569\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIMP3QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIN7U76_LC_19_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60356\,
            in1 => \_gnd_net_\,
            in2 => \N__40467\,
            in3 => \N__40464\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_7_LC_19_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__40458\,
            in1 => \_gnd_net_\,
            in2 => \N__40446\,
            in3 => \N__60202\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_8C_net\,
            ce => \N__59994\,
            sr => \N__62933\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_24_LC_19_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__61125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59702\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_16_LC_19_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59696\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57601\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_28_LC_19_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__62369\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59704\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_8_LC_19_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__63149\,
            in1 => \_gnd_net_\,
            in2 => \N__59728\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_26_LC_19_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59695\,
            in2 => \_gnd_net_\,
            in3 => \N__60914\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_1Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_18_LC_19_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59697\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59852\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_27_LC_19_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__60776\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59703\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_1_LC_19_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59698\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61859\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65553\,
            ce => \N__58879\,
            sr => \N__62924\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISGFN1_LC_19_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55256\,
            in1 => \N__55447\,
            in2 => \N__41053\,
            in3 => \N__40543\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIFMQL2_LC_19_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__40544\,
            in1 => \N__55031\,
            in2 => \N__41054\,
            in3 => \N__54820\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_7_LC_19_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59706\,
            in1 => \N__63476\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65565\,
            ce => \N__49083\,
            sr => \N__62916\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNISSQI1_LC_19_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55446\,
            in1 => \N__55257\,
            in2 => \N__42010\,
            in3 => \N__42577\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_16_LC_19_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59705\,
            in1 => \N__57619\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65565\,
            ce => \N__49083\,
            sr => \N__62916\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIF26H2_LC_19_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__54963\,
            in1 => \N__54819\,
            in2 => \N__42011\,
            in3 => \N__42578\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUIFN1_LC_19_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55258\,
            in1 => \N__55448\,
            in2 => \N__41021\,
            in3 => \N__40822\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_8_LC_19_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59707\,
            in2 => \_gnd_net_\,
            in3 => \N__63150\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65565\,
            ce => \N__49083\,
            sr => \N__62916\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI8NK93_LC_19_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__45869\,
            in1 => \N__40766\,
            in2 => \N__46068\,
            in3 => \N__40721\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SL7_LC_19_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__54004\,
            in1 => \N__40697\,
            in2 => \N__40653\,
            in3 => \N__40806\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIG6SLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIR9DO7_LC_19_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53690\,
            in2 => \N__40650\,
            in3 => \N__40647\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8_LC_19_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__40641\,
            in2 => \N__40626\,
            in3 => \N__55723\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net\,
            ce => \N__55539\,
            sr => \N__62908\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNISLPF7_LC_19_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__40842\,
            in1 => \N__53689\,
            in2 => \_gnd_net_\,
            in3 => \N__40851\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_14_LC_19_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41139\,
            in2 => \N__40836\,
            in3 => \N__55722\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_8C_net\,
            ce => \N__55539\,
            sr => \N__62908\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIHOQL2_LC_19_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55030\,
            in1 => \N__54821\,
            in2 => \N__41020\,
            in3 => \N__40823\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQKV43_LC_19_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__45871\,
            in1 => \N__46042\,
            in2 => \N__49255\,
            in3 => \N__49285\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISAK93_LC_19_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__46043\,
            in1 => \N__45872\,
            in2 => \N__49747\,
            in3 => \N__49948\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISO153_LC_19_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__45873\,
            in1 => \N__46045\,
            in2 => \N__42445\,
            in3 => \N__40973\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUCK93_LC_19_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__46044\,
            in1 => \N__45874\,
            in2 => \N__49636\,
            in3 => \N__49693\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUOV43_LC_19_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__45875\,
            in1 => \N__46046\,
            in2 => \N__41197\,
            in3 => \N__46339\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_10_LC_19_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59640\,
            in2 => \_gnd_net_\,
            in3 => \N__58788\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65588\,
            ce => \N__58867\,
            sr => \N__62898\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_2_LC_19_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59642\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61737\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65588\,
            ce => \N__58867\,
            sr => \N__62898\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_20_LC_19_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59641\,
            in2 => \_gnd_net_\,
            in3 => \N__61531\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65588\,
            ce => \N__58867\,
            sr => \N__62898\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKKQI1_LC_19_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55250\,
            in1 => \N__55409\,
            in2 => \N__42701\,
            in3 => \N__40957\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7Q5H2_LC_19_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55029\,
            in1 => \N__54783\,
            in2 => \N__40962\,
            in3 => \N__42697\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_0_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI788D7_LC_19_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__54001\,
            in1 => \N__41221\,
            in2 => \N__40935\,
            in3 => \N__40932\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_0_i_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIIBPF7_LC_19_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53712\,
            in2 => \N__40926\,
            in3 => \N__40923\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12_LC_19_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46101\,
            in2 => \N__40917\,
            in3 => \N__55695\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net\,
            ce => \N__55538\,
            sr => \N__62887\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8D7_LC_19_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111111111"
        )
    port map (
            in0 => \N__40914\,
            in1 => \N__54002\,
            in2 => \N__40892\,
            in3 => \N__42819\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNICD8DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNINGPF7_LC_19_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53713\,
            in1 => \_gnd_net_\,
            in2 => \N__40860\,
            in3 => \N__40857\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_13_LC_19_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55696\,
            in1 => \_gnd_net_\,
            in2 => \N__41148\,
            in3 => \N__41145\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_12C_net\,
            ce => \N__55538\,
            sr => \N__62887\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_1_LC_19_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59546\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61871\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_2_LC_19_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__61738\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59550\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_5_LC_19_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59547\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63702\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_6_LC_19_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__63584\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59551\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_7_LC_19_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59548\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63471\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_8_LC_19_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59552\,
            in2 => \_gnd_net_\,
            in3 => \N__63145\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_8,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_9_LC_19_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59549\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46523\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_10_LC_19_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58779\,
            in2 => \_gnd_net_\,
            in3 => \N__59545\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65608\,
            ce => \N__45567\,
            sr => \N__62880\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIE9AV5_LC_19_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__60345\,
            in1 => \N__41292\,
            in2 => \_gnd_net_\,
            in3 => \N__41154\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11_LC_19_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49857\,
            in2 => \N__41286\,
            in3 => \N__60164\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net\,
            ce => \N__59984\,
            sr => \N__62871\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GH5_LC_19_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101011111"
        )
    port map (
            in0 => \N__41283\,
            in1 => \N__60516\,
            in2 => \N__41169\,
            in3 => \N__46346\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII0GHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIJEAV5_LC_19_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60346\,
            in2 => \N__41274\,
            in3 => \N__41271\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_12_LC_19_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101100011011000"
        )
    port map (
            in0 => \N__60165\,
            in1 => \N__41265\,
            in2 => \N__41259\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_11C_net\,
            ce => \N__59984\,
            sr => \N__62871\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISV392_17_LC_19_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__58158\,
            in1 => \N__57980\,
            in2 => \N__41238\,
            in3 => \N__41201\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQT392_17_LC_19_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__57979\,
            in1 => \N__58159\,
            in2 => \N__42528\,
            in3 => \N__42554\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFH5_LC_19_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60515\,
            in1 => \N__46376\,
            in2 => \N__41157\,
            in3 => \N__42921\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIDRFHZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIR9FE1_9_LC_19_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__46938\,
            in1 => \N__47042\,
            in2 => \N__56440\,
            in3 => \N__47007\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_7_3_i_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_10_LC_19_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__43059\,
            in1 => \N__41304\,
            in2 => \N__64584\,
            in3 => \N__47380\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65634\,
            ce => \N__50076\,
            sr => \N__64995\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_4_LC_19_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47378\,
            in1 => \N__64582\,
            in2 => \N__41328\,
            in3 => \N__42837\,
            lcout => \s_paddr_I2C_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65634\,
            ce => \N__50076\,
            sr => \N__64995\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_11_LC_19_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110000000"
        )
    port map (
            in0 => \N__64581\,
            in1 => \N__41298\,
            in2 => \N__47403\,
            in3 => \N__43050\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65634\,
            ce => \N__50076\,
            sr => \N__64995\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_9_LC_19_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101010110000000"
        )
    port map (
            in0 => \N__47379\,
            in1 => \N__64583\,
            in2 => \N__41313\,
            in3 => \N__43068\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.s_paddr_I2C_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65634\,
            ce => \N__50076\,
            sr => \N__64995\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIIP1Q6_13_LC_19_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__64713\,
            in1 => \N__55794\,
            in2 => \N__56250\,
            in3 => \N__55988\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1113_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_0_LC_19_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100010111001010"
        )
    port map (
            in0 => \N__55989\,
            in1 => \N__64485\,
            in2 => \N__41316\,
            in3 => \N__46756\,
            lcout => \s_paddr_I2C_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65634\,
            ce => \N__50076\,
            sr => \N__64995\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_0_LC_19_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48292\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.s_addr1_o_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_1_LC_19_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__48157\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.s_addr1_o_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_2_LC_19_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48106\,
            lcout => \I2C_top_level_inst1.s_addr1_o_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_3_LC_19_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48048\,
            lcout => \I2C_top_level_inst1.s_addr1_o_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_4_LC_19_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41378\,
            lcout => \I2C_top_level_inst1.s_addr1_o_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_5_LC_19_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41807\,
            lcout => \I2C_top_level_inst1.s_addr1_o_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_6_LC_19_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41752\,
            lcout => \I2C_top_level_inst1.s_addr1_o_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr1_reg_inst.c_addr1_7_LC_19_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41690\,
            lcout => \I2C_top_level_inst1.s_addr1_o_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47990\,
            ce => \N__41420\,
            sr => \N__62859\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_0_LC_19_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48293\,
            lcout => \I2C_top_level_inst1.s_addr0_o_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_1_LC_19_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48158\,
            lcout => \I2C_top_level_inst1.s_addr0_o_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_2_LC_19_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48107\,
            lcout => \I2C_top_level_inst1.s_addr0_o_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_3_LC_19_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48049\,
            lcout => \I2C_top_level_inst1.s_addr0_o_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_4_LC_19_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41379\,
            lcout => \I2C_top_level_inst1.s_addr0_o_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_5_LC_19_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41808\,
            lcout => \I2C_top_level_inst1.s_addr0_o_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_6_LC_19_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41753\,
            lcout => \I2C_top_level_inst1.s_addr0_o_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.addr0_reg_inst.c_addr0_7_LC_19_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41691\,
            lcout => \I2C_top_level_inst1.s_addr0_o_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47992\,
            ce => \N__43739\,
            sr => \N__62853\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_0_LC_19_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000111110101"
        )
    port map (
            in0 => \N__44142\,
            in1 => \N__47055\,
            in2 => \N__48330\,
            in3 => \N__41619\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_304_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_2_LC_19_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__66769\,
            in1 => \N__56661\,
            in2 => \N__41598\,
            in3 => \N__56818\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_0_LC_19_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__64374\,
            in1 => \N__56376\,
            in2 => \N__41583\,
            in3 => \N__41541\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNOZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_LC_19_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110000001100"
        )
    port map (
            in0 => \N__56181\,
            in1 => \N__41563\,
            in2 => \N__41580\,
            in3 => \N__56594\,
            lcout => \I2C_top_level_inst1.s_no_restart\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65676\,
            ce => 'H',
            sr => \N__65007\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_1_LC_19_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__64794\,
            in1 => \N__48325\,
            in2 => \N__44151\,
            in3 => \N__44141\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_address52_3_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_LC_19_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__66867\,
            in1 => \N__64803\,
            in2 => \N__41517\,
            in3 => \N__41535\,
            lcout => \I2C_top_level_inst1.s_ack\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65685\,
            ce => 'H',
            sr => \N__65011\
        );

    \serializer_mod_inst.shift_reg_6_LC_19_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45461\,
            in1 => \N__41838\,
            in2 => \_gnd_net_\,
            in3 => \N__45040\,
            lcout => \serializer_mod_inst.shift_regZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65700\,
            ce => 'H',
            sr => \N__62836\
        );

    \serializer_mod_inst.shift_reg_64_LC_19_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45039\,
            in1 => \N__44199\,
            in2 => \_gnd_net_\,
            in3 => \N__45460\,
            lcout => \serializer_mod_inst.shift_regZ0Z_64\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65700\,
            ce => 'H',
            sr => \N__62836\
        );

    \serializer_mod_inst.shift_reg_5_LC_19_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011001100"
        )
    port map (
            in0 => \N__41820\,
            in1 => \N__45045\,
            in2 => \_gnd_net_\,
            in3 => \N__45456\,
            lcout => \serializer_mod_inst.shift_regZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65718\,
            ce => 'H',
            sr => \N__62833\
        );

    \serializer_mod_inst.shift_reg_3_LC_19_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47730\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41832\,
            lcout => \serializer_mod_inst.shift_regZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65718\,
            ce => 'H',
            sr => \N__62833\
        );

    \serializer_mod_inst.shift_reg_4_LC_19_24_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41826\,
            in2 => \_gnd_net_\,
            in3 => \N__47731\,
            lcout => \serializer_mod_inst.shift_regZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65718\,
            ce => 'H',
            sr => \N__62833\
        );

    \serializer_mod_inst.shift_reg_28_LC_19_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47729\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41949\,
            lcout => \serializer_mod_inst.shift_regZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65718\,
            ce => 'H',
            sr => \N__62833\
        );

    \serializer_mod_inst.shift_reg_126_LC_19_24_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41886\,
            in2 => \_gnd_net_\,
            in3 => \N__47728\,
            lcout => \serializer_mod_inst.shift_regZ0Z_126\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65718\,
            ce => 'H',
            sr => \N__62833\
        );

    \serializer_mod_inst.shift_reg_24_LC_19_25_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45454\,
            in1 => \N__41937\,
            in2 => \_gnd_net_\,
            in3 => \N__45043\,
            lcout => \serializer_mod_inst.shift_regZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65727\,
            ce => 'H',
            sr => \N__62826\
        );

    \serializer_mod_inst.shift_reg_21_LC_19_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45041\,
            in1 => \N__41904\,
            in2 => \_gnd_net_\,
            in3 => \N__45452\,
            lcout => \serializer_mod_inst.shift_regZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65727\,
            ce => 'H',
            sr => \N__62826\
        );

    \serializer_mod_inst.shift_reg_27_LC_19_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010110001000"
        )
    port map (
            in0 => \N__45455\,
            in1 => \N__41853\,
            in2 => \_gnd_net_\,
            in3 => \N__45044\,
            lcout => \serializer_mod_inst.shift_regZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65727\,
            ce => 'H',
            sr => \N__62826\
        );

    \serializer_mod_inst.shift_reg_23_LC_19_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010010101010"
        )
    port map (
            in0 => \N__45042\,
            in1 => \N__41943\,
            in2 => \_gnd_net_\,
            in3 => \N__45453\,
            lcout => \serializer_mod_inst.shift_regZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65727\,
            ce => 'H',
            sr => \N__62826\
        );

    \serializer_mod_inst.shift_reg_109_LC_19_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41931\,
            in2 => \_gnd_net_\,
            in3 => \N__47706\,
            lcout => \serializer_mod_inst.shift_regZ0Z_109\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65727\,
            ce => 'H',
            sr => \N__62826\
        );

    \serializer_mod_inst.shift_reg_20_LC_19_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47707\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41913\,
            lcout => \serializer_mod_inst.shift_regZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65727\,
            ce => 'H',
            sr => \N__62826\
        );

    \serializer_mod_inst.shift_reg_124_LC_19_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41865\,
            in2 => \_gnd_net_\,
            in3 => \N__47646\,
            lcout => \serializer_mod_inst.shift_regZ0Z_124\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65737\,
            ce => 'H',
            sr => \N__62821\
        );

    \serializer_mod_inst.shift_reg_25_LC_19_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41898\,
            in2 => \_gnd_net_\,
            in3 => \N__47648\,
            lcout => \serializer_mod_inst.shift_regZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65737\,
            ce => 'H',
            sr => \N__62821\
        );

    \serializer_mod_inst.shift_reg_125_LC_19_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47647\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41892\,
            lcout => \serializer_mod_inst.shift_regZ0Z_125\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65737\,
            ce => 'H',
            sr => \N__62821\
        );

    \serializer_mod_inst.shift_reg_123_LC_19_26_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__41877\,
            in2 => \_gnd_net_\,
            in3 => \N__47645\,
            lcout => \serializer_mod_inst.shift_regZ0Z_123\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65737\,
            ce => 'H',
            sr => \N__62821\
        );

    \serializer_mod_inst.shift_reg_26_LC_19_26_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47649\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__41859\,
            lcout => \serializer_mod_inst.shift_regZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65737\,
            ce => 'H',
            sr => \N__62821\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_27_LC_20_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__42144\,
            in1 => \N__52771\,
            in2 => \N__42126\,
            in3 => \N__52526\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_27_LC_20_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000011110000"
        )
    port map (
            in0 => \N__49143\,
            in1 => \_gnd_net_\,
            in2 => \N__42105\,
            in3 => \N__52231\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_27_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_27_LC_20_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__42102\,
            in1 => \N__42096\,
            in2 => \N__42084\,
            in3 => \N__42060\,
            lcout => \I2C_top_level_inst1_s_data_oreg_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65534\,
            ce => \N__54500\,
            sr => \N__65023\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_27_LC_20_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100000000"
        )
    port map (
            in0 => \N__51921\,
            in1 => \N__42081\,
            in2 => \N__48504\,
            in3 => \N__42072\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_16_LC_20_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__52998\,
            in1 => \N__53524\,
            in2 => \N__53323\,
            in3 => \N__54207\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_16_LC_20_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__42054\,
            in1 => \N__52745\,
            in2 => \N__42036\,
            in3 => \N__52492\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_16_LC_20_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52187\,
            in2 => \N__42015\,
            in3 => \N__42012\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_16_LC_20_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__44432\,
            in1 => \N__41988\,
            in2 => \N__63134\,
            in3 => \N__44658\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_16_LC_20_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__41970\,
            in1 => \N__51922\,
            in2 => \N__41952\,
            in3 => \N__51657\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_16_LC_20_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__42336\,
            in1 => \N__42327\,
            in2 => \N__42321\,
            in3 => \N__42318\,
            lcout => \I2C_top_level_inst1_s_data_oreg_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65554\,
            ce => \N__54497\,
            sr => \N__65018\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_24_LC_20_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__42312\,
            in1 => \N__44657\,
            in2 => \N__57608\,
            in3 => \N__44431\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_22_LC_20_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59587\,
            in1 => \N__61348\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_3_LC_20_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59589\,
            in2 => \_gnd_net_\,
            in3 => \N__63940\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_4_LC_20_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59727\,
            in2 => \_gnd_net_\,
            in3 => \N__63827\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_5_LC_20_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59590\,
            in2 => \_gnd_net_\,
            in3 => \N__63687\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_6_LC_20_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59588\,
            in1 => \N__63581\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_7_LC_20_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59591\,
            in2 => \_gnd_net_\,
            in3 => \N__63483\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_17_LC_20_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59726\,
            in2 => \_gnd_net_\,
            in3 => \N__57392\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_9_LC_20_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59592\,
            in2 => \_gnd_net_\,
            in3 => \N__46500\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65566\,
            ce => \N__58880\,
            sr => \N__62934\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIQQQI1_LC_20_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__46597\,
            in1 => \N__55249\,
            in2 => \N__42608\,
            in3 => \N__55449\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNID06H2_LC_20_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__55056\,
            in1 => \N__46598\,
            in2 => \N__54835\,
            in3 => \N__42604\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8D7_LC_20_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53993\,
            in1 => \N__53371\,
            in2 => \N__42387\,
            in3 => \N__45546\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIMN8DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI1RPF7_LC_20_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53714\,
            in2 => \N__42384\,
            in3 => \N__42381\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15_LC_20_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__42375\,
            in1 => \_gnd_net_\,
            in2 => \N__42369\,
            in3 => \N__55724\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net\,
            ce => \N__55570\,
            sr => \N__62925\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8D7_LC_20_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53960\,
            in1 => \N__54206\,
            in2 => \N__42366\,
            in3 => \N__45540\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIRS8DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI60QF7_LC_20_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53715\,
            in1 => \_gnd_net_\,
            in2 => \N__42357\,
            in3 => \N__42354\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_16_LC_20_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55725\,
            in1 => \_gnd_net_\,
            in2 => \N__42348\,
            in3 => \N__42345\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_15C_net\,
            ce => \N__55570\,
            sr => \N__62925\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_1_LC_20_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61860\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_2_LC_20_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61745\,
            in2 => \_gnd_net_\,
            in3 => \N__59511\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_3_LC_20_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__63945\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_4_LC_20_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__63789\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59512\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_9_LC_20_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59516\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__46530\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_10_LC_20_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58796\,
            in2 => \_gnd_net_\,
            in3 => \N__59509\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_11_LC_20_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59513\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58691\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_20_LC_20_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59510\,
            in2 => \_gnd_net_\,
            in3 => \N__61546\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65589\,
            ce => \N__48724\,
            sr => \N__62917\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_20_LC_20_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59428\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61547\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_12_LC_20_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__58590\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59430\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_21_LC_20_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59429\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61437\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_22_LC_20_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61356\,
            in2 => \_gnd_net_\,
            in3 => \N__59424\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_22,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_14_LC_20_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59426\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58499\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_23_LC_20_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61248\,
            in2 => \_gnd_net_\,
            in3 => \N__59425\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_15_LC_20_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59427\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57535\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_16_LC_20_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57618\,
            in2 => \_gnd_net_\,
            in3 => \N__59423\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65601\,
            ce => \N__45571\,
            sr => \N__62909\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNISMV43_LC_20_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__46064\,
            in1 => \N__46369\,
            in2 => \N__45921\,
            in3 => \N__42550\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238D7_LC_20_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__42514\,
            in1 => \N__54003\,
            in2 => \N__42489\,
            in3 => \N__42825\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI238DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID6PF7_LC_20_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__46115\,
            in1 => \_gnd_net_\,
            in2 => \N__42828\,
            in3 => \N__53673\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5O5H2_LC_20_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__54781\,
            in1 => \N__42940\,
            in2 => \N__55052\,
            in3 => \N__42905\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_11_LC_20_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__58701\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59431\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65609\,
            ce => \N__45569\,
            sr => \N__62899\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI9S5H2_LC_20_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55022\,
            in1 => \N__54782\,
            in2 => \N__46159\,
            in3 => \N__42793\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_13_LC_20_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58376\,
            in2 => \_gnd_net_\,
            in3 => \N__59432\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65609\,
            ce => \N__45569\,
            sr => \N__62899\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIB08H2_LC_20_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__54780\,
            in1 => \N__49480\,
            in2 => \N__55053\,
            in3 => \N__49453\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIGGQI1_LC_20_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55231\,
            in1 => \N__55427\,
            in2 => \N__42728\,
            in3 => \N__42751\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3M5H2_LC_20_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__42724\,
            in1 => \N__55020\,
            in2 => \N__42758\,
            in3 => \N__54818\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_10_LC_20_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59422\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58797\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_10,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65622\,
            ce => \N__49063\,
            sr => \N__62888\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNII6FN1_LC_20_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55429\,
            in1 => \N__55232\,
            in2 => \N__43004\,
            in3 => \N__42964\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_2_LC_20_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59421\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61719\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65622\,
            ce => \N__49063\,
            sr => \N__62888\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI5CQL2_LC_20_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55021\,
            in1 => \N__54817\,
            in2 => \N__43003\,
            in3 => \N__42965\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIIIQI1_LC_20_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55230\,
            in1 => \N__55428\,
            in2 => \N__42944\,
            in3 => \N__42904\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_11_LC_20_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59420\,
            in2 => \_gnd_net_\,
            in3 => \N__58700\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65622\,
            ce => \N__49063\,
            sr => \N__62888\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_c_0_LC_20_17_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__55982\,
            in2 => \N__46763\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_20_17_0_\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_1_LC_20_17_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46824\,
            in2 => \_gnd_net_\,
            in3 => \N__42873\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_1\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_0\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_2_LC_20_17_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46907\,
            in2 => \_gnd_net_\,
            in3 => \N__42855\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_2\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_1\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_LUT4_0_LC_20_17_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54338\,
            in2 => \_gnd_net_\,
            in3 => \N__42840\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_2\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_4_LC_20_17_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47197\,
            in2 => \_gnd_net_\,
            in3 => \N__42831\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_4\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_3\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_5_LC_20_17_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47247\,
            in2 => \_gnd_net_\,
            in3 => \N__43104\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_5\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_4\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_6_LC_20_17_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47170\,
            in2 => \_gnd_net_\,
            in3 => \N__43089\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_6\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_5\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_7_LC_20_17_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47118\,
            in2 => \_gnd_net_\,
            in3 => \N__43074\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_7\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_6\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_LUT4_0_LC_20_18_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56122\,
            in2 => \_gnd_net_\,
            in3 => \N__43071\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_20_18_0_\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_9_LC_20_18_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47008\,
            in2 => \_gnd_net_\,
            in3 => \N__43062\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_9\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_8\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_10_LC_20_18_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47037\,
            in2 => \_gnd_net_\,
            in3 => \N__43053\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_10\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_9\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_11_LC_20_18_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__46942\,
            in2 => \_gnd_net_\,
            in3 => \N__43044\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_11\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_10\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_12_LC_20_18_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43041\,
            in2 => \_gnd_net_\,
            in3 => \N__43008\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_12\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_11\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_13_LC_20_18_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43275\,
            in2 => \_gnd_net_\,
            in3 => \N__43245\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_13\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_12\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_14_LC_20_18_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43242\,
            in2 => \_gnd_net_\,
            in3 => \N__43212\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_14\,
            ltout => OPEN,
            carryin => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_13\,
            carryout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_15_LC_20_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43209\,
            in2 => \_gnd_net_\,
            in3 => \N__43188\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_s_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_13_LC_20_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__56621\,
            in1 => \N__66264\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_103_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_2_LC_20_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43158\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_1_LC_20_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43152\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_q_0_LC_20_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43746\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.start_inter_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65661\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIABID_21_LC_20_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__56232\,
            in1 => \N__43619\,
            in2 => \_gnd_net_\,
            in3 => \N__43146\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_291\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_291_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_0_LC_20_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001010000"
        )
    port map (
            in0 => \N__66794\,
            in1 => \N__56620\,
            in2 => \N__43119\,
            in3 => \N__57237\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_new_address_RNO_0_LC_20_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__43747\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43669\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.un1_c_state_6_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_FSM_inst.c_state_RNO_0_0_LC_20_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011011101"
        )
    port map (
            in0 => \N__43670\,
            in1 => \N__50886\,
            in2 => \_gnd_net_\,
            in3 => \N__43836\,
            lcout => \I2C_top_level_inst1.I2C_FSM_inst.N_1378\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI5MGJ_2_LC_20_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__65871\,
            in1 => \N__56361\,
            in2 => \N__64789\,
            in3 => \N__56816\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.m24_i_a3_LC_20_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000101"
        )
    port map (
            in0 => \N__56817\,
            in1 => \N__66273\,
            in2 => \N__65986\,
            in3 => \N__65872\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_op_inst1.N_1676_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_2_LC_20_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__66165\,
            in1 => \N__64343\,
            in2 => \N__43626\,
            in3 => \N__62455\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65677\,
            ce => 'H',
            sr => \N__65008\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_22_LC_20_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001000100010"
        )
    port map (
            in0 => \N__43623\,
            in1 => \N__66164\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65677\,
            ce => 'H',
            sr => \N__65008\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIEVJ7_22_LC_20_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65974\,
            in2 => \_gnd_net_\,
            in3 => \N__56815\,
            lcout => \c_state_RNIEVJ7_22\,
            ltout => \c_state_RNIEVJ7_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASSA_22_LC_20_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__43587\,
            in3 => \N__43513\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_77_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF6Q22_14_LC_20_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__57123\,
            in1 => \N__57089\,
            in2 => \N__43299\,
            in3 => \N__64432\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_0_LC_20_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__43955\,
            in1 => \N__43905\,
            in2 => \_gnd_net_\,
            in3 => \N__48290\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_2_1_4_LC_20_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48195\,
            in2 => \_gnd_net_\,
            in3 => \N__50112\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1606_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_2_LC_20_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__43767\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_0_LC_20_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__43857\,
            in1 => \N__43829\,
            in2 => \_gnd_net_\,
            in3 => \N__43794\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_2_LC_20_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43755\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_ready_slave_addr_q_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_1_LC_20_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43773\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_15_LC_20_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__66150\,
            in1 => \N__48310\,
            in2 => \_gnd_net_\,
            in3 => \N__44140\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_607\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_q_1_LC_20_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43761\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.ready_slave_addr_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65686\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI1I79_18_LC_20_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__47563\,
            in1 => \N__50536\,
            in2 => \_gnd_net_\,
            in3 => \N__56584\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_294\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_4_LC_20_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47562\,
            in2 => \_gnd_net_\,
            in3 => \N__56729\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_0_1_LC_20_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56583\,
            in2 => \_gnd_net_\,
            in3 => \N__50113\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1353_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_RNISHA8_2_LC_20_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__50537\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50933\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_305_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_0_LC_20_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48291\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65701\,
            ce => \N__44061\,
            sr => \N__65019\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rx_1_LC_20_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48156\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_data_rxZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65701\,
            ce => \N__44061\,
            sr => \N__65019\
        );

    \serializer_mod_inst.shift_reg_65_LC_20_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110001000"
        )
    port map (
            in0 => \N__44025\,
            in1 => \N__45446\,
            in2 => \_gnd_net_\,
            in3 => \N__45046\,
            lcout => \serializer_mod_inst.shift_regZ0Z_65\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65719\,
            ce => 'H',
            sr => \N__62842\
        );

    \serializer_mod_inst.shift_reg_128_LC_20_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47814\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__43968\,
            lcout => \serializer_mod_inst.shift_regZ0Z_128\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65719\,
            ce => 'H',
            sr => \N__62842\
        );

    \serializer_mod_inst.shift_reg_127_LC_20_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43974\,
            in2 => \_gnd_net_\,
            in3 => \N__47813\,
            lcout => \serializer_mod_inst.shift_regZ0Z_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65719\,
            ce => 'H',
            sr => \N__62842\
        );

    \serializer_mod_inst.shift_reg_29_LC_20_24_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__43962\,
            in2 => \_gnd_net_\,
            in3 => \N__47724\,
            lcout => \serializer_mod_inst.shift_regZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65728\,
            ce => 'H',
            sr => \N__62837\
        );

    \serializer_mod_inst.shift_reg_62_LC_20_24_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47726\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44175\,
            lcout => \serializer_mod_inst.shift_regZ0Z_62\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65728\,
            ce => 'H',
            sr => \N__62837\
        );

    \serializer_mod_inst.shift_reg_30_LC_20_24_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44220\,
            lcout => \serializer_mod_inst.shift_regZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65728\,
            ce => 'H',
            sr => \N__62837\
        );

    \serializer_mod_inst.shift_reg_63_LC_20_24_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44205\,
            lcout => \serializer_mod_inst.shift_regZ0Z_63\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65728\,
            ce => 'H',
            sr => \N__62837\
        );

    \serializer_mod_inst.shift_reg_58_LC_20_25_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44157\,
            in2 => \_gnd_net_\,
            in3 => \N__47651\,
            lcout => \serializer_mod_inst.shift_regZ0Z_58\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65738\,
            ce => 'H',
            sr => \N__62834\
        );

    \serializer_mod_inst.shift_reg_59_LC_20_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44193\,
            lcout => \serializer_mod_inst.shift_regZ0Z_59\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65738\,
            ce => 'H',
            sr => \N__62834\
        );

    \serializer_mod_inst.shift_reg_60_LC_20_25_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44187\,
            in2 => \_gnd_net_\,
            in3 => \N__47653\,
            lcout => \serializer_mod_inst.shift_regZ0Z_60\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65738\,
            ce => 'H',
            sr => \N__62834\
        );

    \serializer_mod_inst.shift_reg_61_LC_20_25_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__47654\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__44181\,
            lcout => \serializer_mod_inst.shift_regZ0Z_61\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65738\,
            ce => 'H',
            sr => \N__62834\
        );

    \serializer_mod_inst.shift_reg_57_LC_20_25_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__44169\,
            in2 => \_gnd_net_\,
            in3 => \N__47650\,
            lcout => \serializer_mod_inst.shift_regZ0Z_57\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65738\,
            ce => 'H',
            sr => \N__62834\
        );

    \serializer_mod_inst.current_state_RNIVDDK_0_0_LC_20_26_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__45201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__45035\,
            lcout => \serializer_mod_inst.current_state_RNIVDDK_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.current_state_RNO_1_0_LC_20_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48430\,
            in2 => \_gnd_net_\,
            in3 => \N__48478\,
            lcout => OPEN,
            ltout => \serializer_mod_inst.un22_next_state_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.current_state_RNO_0_0_LC_20_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__48616\,
            in1 => \N__48458\,
            in2 => \N__45501\,
            in3 => \N__48489\,
            lcout => \serializer_mod_inst.un22_next_state\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.current_state_RNIVDDK_0_LC_20_27_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__45402\,
            in2 => \_gnd_net_\,
            in3 => \N__45088\,
            lcout => \serializer_mod_inst.next_state32_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_0_LC_21_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__44244\,
            in1 => \N__44250\,
            in2 => \N__44721\,
            in3 => \N__44706\,
            lcout => \I2C_top_level_inst1_s_data_oreg_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65535\,
            ce => \N__54501\,
            sr => \N__65028\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_5_0_LC_21_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__44691\,
            in1 => \N__44676\,
            in2 => \N__44454\,
            in3 => \N__44433\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_0_LC_21_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__44274\,
            in1 => \N__51920\,
            in2 => \N__44253\,
            in3 => \N__58256\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_0_LC_21_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__58227\,
            in1 => \N__53014\,
            in2 => \N__53310\,
            in3 => \N__60645\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_25_LC_21_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__61018\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59717\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf4_c_data_system_o_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65567\,
            ce => \N__45573\,
            sr => \N__62946\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_17_LC_21_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__57412\,
            in1 => \_gnd_net_\,
            in2 => \N__59729\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65567\,
            ce => \N__45573\,
            sr => \N__62946\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_26_LC_21_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59718\,
            in2 => \_gnd_net_\,
            in3 => \N__60905\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_3Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65567\,
            ce => \N__45573\,
            sr => \N__62946\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_18_LC_21_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__59844\,
            in1 => \_gnd_net_\,
            in2 => \N__59730\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65567\,
            ce => \N__45573\,
            sr => \N__62946\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_19_LC_21_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59716\,
            in2 => \_gnd_net_\,
            in3 => \N__61644\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65567\,
            ce => \N__45573\,
            sr => \N__62946\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf4.c_data_system_o_0_LC_21_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59719\,
            in1 => \N__61930\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkstopmask_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65567\,
            ce => \N__45573\,
            sr => \N__62946\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI4VV43_LC_21_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__45903\,
            in1 => \N__46056\,
            in2 => \N__48565\,
            in3 => \N__46198\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI61053_LC_21_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__46054\,
            in1 => \N__45904\,
            in2 => \N__53525\,
            in3 => \N__51652\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI6LK93_LC_21_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__46057\,
            in1 => \N__45530\,
            in2 => \N__45919\,
            in3 => \N__48745\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIA5053_LC_21_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__46055\,
            in1 => \N__45905\,
            in2 => \N__51434\,
            in3 => \N__51364\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIAPK93_LC_21_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__45906\,
            in1 => \N__46052\,
            in2 => \N__49382\,
            in3 => \N__49819\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIC7053_LC_21_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__46053\,
            in1 => \N__45907\,
            in2 => \N__51505\,
            in3 => \N__57323\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIO6K93_LC_21_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010001011110011"
        )
    port map (
            in0 => \N__46058\,
            in1 => \N__60641\,
            in2 => \N__45920\,
            in3 => \N__58246\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIQ8K93_LC_21_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__46051\,
            in1 => \N__45908\,
            in2 => \N__60709\,
            in3 => \N__57826\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIUUQI1_LC_21_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55262\,
            in1 => \N__55450\,
            in2 => \N__46556\,
            in3 => \N__45613\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNI83053_LC_21_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__45902\,
            in1 => \N__46059\,
            in2 => \N__51588\,
            in3 => \N__51610\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029D7_LC_21_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53961\,
            in1 => \N__54152\,
            in2 => \N__45645\,
            in3 => \N__45594\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI029DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIB5QF7_LC_21_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53721\,
            in2 => \N__45642\,
            in3 => \N__45639\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17_LC_21_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55744\,
            in1 => \_gnd_net_\,
            in2 => \N__45633\,
            in3 => \N__45630\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net\,
            ce => \N__55558\,
            sr => \N__62935\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIH46H2_LC_21_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111100100011"
        )
    port map (
            in0 => \N__54816\,
            in1 => \N__46552\,
            in2 => \N__45618\,
            in3 => \N__55055\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_0_LC_21_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__55742\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48878\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net\,
            ce => \N__55558\,
            sr => \N__62935\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_11_LC_21_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__46686\,
            in1 => \N__55743\,
            in2 => \_gnd_net_\,
            in3 => \N__46116\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_17C_net\,
            ce => \N__55558\,
            sr => \N__62935\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIS1692_17_LC_21_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__57981\,
            in1 => \N__58179\,
            in2 => \N__45743\,
            in3 => \N__45763\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LH5_LC_21_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60597\,
            in1 => \N__46306\,
            in2 => \N__46089\,
            in3 => \N__46074\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNII5LHZ0Z5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIKMSI1_LC_21_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55254\,
            in1 => \N__55444\,
            in2 => \N__45674\,
            in3 => \N__45691\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_21_LC_21_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59508\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61435\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65602\,
            ce => \N__49093\,
            sr => \N__62926\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_6_RNIUQ153_LC_21_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110101"
        )
    port map (
            in0 => \N__46307\,
            in1 => \N__46060\,
            in2 => \N__45870\,
            in3 => \N__45764\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_2_21_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDD7_LC_21_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__45742\,
            in1 => \N__53966\,
            in2 => \N__45711\,
            in3 => \N__45651\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI7DDDZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI7S7H2_LC_21_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__54806\,
            in1 => \N__45692\,
            in2 => \N__55019\,
            in3 => \N__45670\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_11_LC_21_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__58696\,
            in2 => \_gnd_net_\,
            in3 => \N__59416\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_11,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_12_LC_21_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59412\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58591\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_12,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_21_LC_21_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61434\,
            in2 => \_gnd_net_\,
            in3 => \N__59418\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_21,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_30_LC_21_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__59415\,
            in1 => \_gnd_net_\,
            in2 => \N__62183\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_13_LC_21_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__58364\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59417\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_25_LC_21_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59414\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61019\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_31_LC_21_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62072\,
            in2 => \_gnd_net_\,
            in3 => \N__59419\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_15_LC_21_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59413\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57536\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65610\,
            ce => \N__58868\,
            sr => \N__62918\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_13_LC_21_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59433\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58377\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_13,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_31_LC_21_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59439\,
            in2 => \_gnd_net_\,
            in3 => \N__62073\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_23_LC_21_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59435\,
            in1 => \N__61254\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_15_LC_21_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59437\,
            in2 => \_gnd_net_\,
            in3 => \N__57540\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_24_LC_21_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59436\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61117\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_25_LC_21_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59438\,
            in2 => \_gnd_net_\,
            in3 => \N__61013\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_17_LC_21_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59434\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57414\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_9_LC_21_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59440\,
            in2 => \_gnd_net_\,
            in3 => \N__46526\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_9,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65623\,
            ce => \N__49071\,
            sr => \N__62910\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSL7_LC_21_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53967\,
            in1 => \N__49427\,
            in2 => \N__46419\,
            in3 => \N__46614\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILBSLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI0FDO7_LC_21_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53674\,
            in2 => \N__46404\,
            in3 => \N__46401\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9_LC_21_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55727\,
            in1 => \_gnd_net_\,
            in2 => \N__46395\,
            in3 => \N__46392\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net\,
            ce => \N__55571\,
            sr => \N__62900\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7D7_LC_21_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010111111111"
        )
    port map (
            in0 => \N__46725\,
            in1 => \N__53968\,
            in2 => \N__49344\,
            in3 => \N__46710\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITT7DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI81PF7_LC_21_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53675\,
            in1 => \_gnd_net_\,
            in2 => \N__46704\,
            in3 => \N__46701\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_10_LC_21_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__46695\,
            in1 => \_gnd_net_\,
            in2 => \N__46689\,
            in3 => \N__55726\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_9C_net\,
            ce => \N__55571\,
            sr => \N__62900\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI0LFN1_LC_21_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55255\,
            in1 => \N__55430\,
            in2 => \N__46667\,
            in3 => \N__46627\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJQQL2_LC_21_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__46660\,
            in1 => \N__55036\,
            in2 => \N__46634\,
            in3 => \N__54834\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_0_4_LC_21_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__47168\,
            in1 => \N__47244\,
            in2 => \N__47122\,
            in3 => \N__47207\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_93_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_3_LC_21_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111110101"
        )
    port map (
            in0 => \N__56127\,
            in1 => \N__56057\,
            in2 => \N__46608\,
            in3 => \N__54335\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1590_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_2_LC_21_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__50545\,
            in1 => \N__56128\,
            in2 => \_gnd_net_\,
            in3 => \N__55916\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_1_LC_21_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101001100"
        )
    port map (
            in0 => \N__54402\,
            in1 => \N__55868\,
            in2 => \N__46965\,
            in3 => \N__55796\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIOK81_4_LC_21_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__47169\,
            in1 => \N__47245\,
            in2 => \N__47123\,
            in3 => \N__47208\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_1_LC_21_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__47171\,
            in1 => \N__46980\,
            in2 => \N__47124\,
            in3 => \N__47061\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIOFAP_9_LC_21_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__47041\,
            in2 => \_gnd_net_\,
            in3 => \N__47012\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_o2_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_ack_RNO_3_LC_21_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__46813\,
            in1 => \N__46762\,
            in2 => \N__46908\,
            in3 => \N__54337\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_n_no_restart_2_sqmuxa_i_a3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_LC_21_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__46761\,
            in1 => \N__46892\,
            in2 => \_gnd_net_\,
            in3 => \N__46812\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1577_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIB9ER2_0_3_LC_21_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46974\,
            in1 => \N__56129\,
            in2 => \N__46968\,
            in3 => \N__54336\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1586_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_11_LC_21_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__46956\,
            in1 => \N__46946\,
            in2 => \N__46914\,
            in3 => \N__47468\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1591_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIG4FU_0_0_LC_21_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__46891\,
            in1 => \N__46811\,
            in2 => \_gnd_net_\,
            in3 => \N__46760\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1575_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIKPI66_9_LC_21_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__47478\,
            in1 => \N__50192\,
            in2 => \_gnd_net_\,
            in3 => \N__47469\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_394\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIGUM51_1_LC_21_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010101010101"
        )
    port map (
            in0 => \N__64679\,
            in1 => \N__56574\,
            in2 => \N__48222\,
            in3 => \N__55857\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_935_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNICOOV_1_LC_21_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__55853\,
            in1 => \_gnd_net_\,
            in2 => \N__56591\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_8_LC_21_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101111"
        )
    port map (
            in0 => \N__47445\,
            in1 => \_gnd_net_\,
            in2 => \N__47436\,
            in3 => \N__47426\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_8_LC_21_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101000111100010"
        )
    port map (
            in0 => \N__56123\,
            in1 => \N__47413\,
            in2 => \N__47328\,
            in3 => \N__47325\,
            lcout => \s_paddr_I2C_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65678\,
            ce => \N__50052\,
            sr => \N__65009\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_1_LC_21_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111110101010"
        )
    port map (
            in0 => \N__47319\,
            in1 => \_gnd_net_\,
            in2 => \N__48220\,
            in3 => \N__55855\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1651\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_1_2_LC_21_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100100010"
        )
    port map (
            in0 => \N__55854\,
            in1 => \N__48209\,
            in2 => \_gnd_net_\,
            in3 => \N__47286\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1652\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_4_LC_21_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010101010"
        )
    port map (
            in0 => \N__64472\,
            in1 => \_gnd_net_\,
            in2 => \N__48221\,
            in3 => \N__55856\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_4_LC_21_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__56489\,
            in1 => \N__50681\,
            in2 => \N__47250\,
            in3 => \N__56469\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_14_LC_21_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101011111"
        )
    port map (
            in0 => \N__47493\,
            in1 => \N__56027\,
            in2 => \N__66609\,
            in3 => \N__48205\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_14_LC_21_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__66125\,
            in1 => \N__64696\,
            in2 => \_gnd_net_\,
            in3 => \N__50137\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_0_1_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_17_LC_21_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101010101"
        )
    port map (
            in0 => \N__64697\,
            in1 => \N__66324\,
            in2 => \_gnd_net_\,
            in3 => \N__65914\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_279_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_17_LC_21_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010000000101"
        )
    port map (
            in0 => \N__66129\,
            in1 => \N__66325\,
            in2 => \N__47487\,
            in3 => \N__66607\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65687\,
            ce => 'H',
            sr => \N__65012\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_7_LC_21_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__66375\,
            in1 => \N__62406\,
            in2 => \N__66156\,
            in3 => \N__50138\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_0_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_7_LC_21_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__55862\,
            in1 => \N__56028\,
            in2 => \N__47484\,
            in3 => \N__66376\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65687\,
            ce => 'H',
            sr => \N__65012\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_20_LC_21_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__55861\,
            in1 => \N__50682\,
            in2 => \N__48219\,
            in3 => \N__64473\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65687\,
            ce => 'H',
            sr => \N__65012\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_9_LC_21_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__50544\,
            in1 => \N__50930\,
            in2 => \N__56520\,
            in3 => \N__57287\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_268_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_9_LC_21_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__66603\,
            in1 => \N__50643\,
            in2 => \N__47481\,
            in3 => \N__50166\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65702\,
            ce => 'H',
            sr => \N__65020\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_10_LC_21_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50642\,
            in2 => \_gnd_net_\,
            in3 => \N__66602\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_10_LC_21_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111010100110000"
        )
    port map (
            in0 => \N__66109\,
            in1 => \N__47510\,
            in2 => \N__47571\,
            in3 => \N__66755\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65702\,
            ce => 'H',
            sr => \N__65020\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_18_LC_21_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111001100"
        )
    port map (
            in0 => \N__50721\,
            in1 => \N__47564\,
            in2 => \_gnd_net_\,
            in3 => \N__50543\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_18_LC_21_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__66110\,
            in1 => \_gnd_net_\,
            in2 => \N__47568\,
            in3 => \N__50932\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65702\,
            ce => 'H',
            sr => \N__65020\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_8_LC_21_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__50931\,
            in1 => \N__66111\,
            in2 => \_gnd_net_\,
            in3 => \N__47565\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65702\,
            ce => 'H',
            sr => \N__65020\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_o2_26_LC_21_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011000000000"
        )
    port map (
            in0 => \N__51078\,
            in1 => \N__51052\,
            in2 => \N__51023\,
            in3 => \N__51121\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1605_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_0_0_LC_21_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__48181\,
            in1 => \N__51076\,
            in2 => \_gnd_net_\,
            in3 => \N__47526\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_burst16_0_o2_LC_21_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__51013\,
            in1 => \N__51048\,
            in2 => \_gnd_net_\,
            in3 => \N__51118\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_107_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_14_LC_21_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__48183\,
            in1 => \N__64433\,
            in2 => \N__47520\,
            in3 => \N__51079\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_a3_1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNI68137_11_LC_21_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__56173\,
            in1 => \N__50004\,
            in2 => \_gnd_net_\,
            in3 => \N__48182\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1600_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.un1_command_1_i_i_o2_LC_21_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__51119\,
            in1 => \N__51014\,
            in2 => \N__51054\,
            in3 => \N__51075\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_315_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_o4_1_1_a3_0_o2_4_LC_21_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__51120\,
            in1 => \N__51015\,
            in2 => \_gnd_net_\,
            in3 => \N__51077\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_403_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_0_LC_21_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48294\,
            lcout => \I2C_top_level_inst1.s_command_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47996\,
            ce => \N__47931\,
            sr => \N__62848\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_1_LC_21_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48162\,
            lcout => \I2C_top_level_inst1.s_command_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47996\,
            ce => \N__47931\,
            sr => \N__62848\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_2_LC_21_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48111\,
            lcout => \I2C_top_level_inst1.s_command_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47996\,
            ce => \N__47931\,
            sr => \N__62848\
        );

    \I2C_top_level_inst1.command_reg_inst.c_command_3_LC_21_23_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__48056\,
            lcout => \I2C_top_level_inst1.s_command_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__47996\,
            ce => \N__47931\,
            sr => \N__62848\
        );

    \serializer_mod_inst.counter_sr_RNIO9BB_0_LC_21_25_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__48357\,
            in1 => \N__48435\,
            in2 => \_gnd_net_\,
            in3 => \N__48483\,
            lcout => \serializer_mod_inst.un1_counter_srlto6_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.counter_sr_RNIDF4F_1_LC_21_26_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48374\,
            in1 => \N__48392\,
            in2 => \N__48459\,
            in3 => \N__48410\,
            lcout => OPEN,
            ltout => \serializer_mod_inst.un1_counter_srlto6_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.counter_sr_RNIREMI1_7_LC_21_26_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101010111111111"
        )
    port map (
            in0 => \N__48617\,
            in1 => \N__47892\,
            in2 => \N__47886\,
            in3 => \N__47644\,
            lcout => \serializer_mod_inst.counter_sre_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.current_state_RNO_2_0_LC_21_26_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__48373\,
            in1 => \N__48391\,
            in2 => \N__48356\,
            in3 => \N__48409\,
            lcout => \serializer_mod_inst.un22_next_state_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \serializer_mod_inst.counter_sr_0_LC_21_27_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48651\,
            in1 => \N__48482\,
            in2 => \_gnd_net_\,
            in3 => \N__48462\,
            lcout => \serializer_mod_inst.counter_srZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_21_27_0_\,
            carryout => \serializer_mod_inst.counter_sr_cry_0\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_1_LC_21_27_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48638\,
            in1 => \N__48457\,
            in2 => \_gnd_net_\,
            in3 => \N__48438\,
            lcout => \serializer_mod_inst.counter_srZ0Z_1\,
            ltout => OPEN,
            carryin => \serializer_mod_inst.counter_sr_cry_0\,
            carryout => \serializer_mod_inst.counter_sr_cry_1\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_2_LC_21_27_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48652\,
            in1 => \N__48434\,
            in2 => \_gnd_net_\,
            in3 => \N__48414\,
            lcout => \serializer_mod_inst.counter_srZ0Z_2\,
            ltout => OPEN,
            carryin => \serializer_mod_inst.counter_sr_cry_1\,
            carryout => \serializer_mod_inst.counter_sr_cry_2\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_3_LC_21_27_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48639\,
            in1 => \N__48411\,
            in2 => \_gnd_net_\,
            in3 => \N__48396\,
            lcout => \serializer_mod_inst.counter_srZ0Z_3\,
            ltout => OPEN,
            carryin => \serializer_mod_inst.counter_sr_cry_2\,
            carryout => \serializer_mod_inst.counter_sr_cry_3\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_4_LC_21_27_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48653\,
            in1 => \N__48393\,
            in2 => \_gnd_net_\,
            in3 => \N__48378\,
            lcout => \serializer_mod_inst.counter_srZ0Z_4\,
            ltout => OPEN,
            carryin => \serializer_mod_inst.counter_sr_cry_3\,
            carryout => \serializer_mod_inst.counter_sr_cry_4\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_5_LC_21_27_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48640\,
            in1 => \N__48375\,
            in2 => \_gnd_net_\,
            in3 => \N__48360\,
            lcout => \serializer_mod_inst.counter_srZ0Z_5\,
            ltout => OPEN,
            carryin => \serializer_mod_inst.counter_sr_cry_4\,
            carryout => \serializer_mod_inst.counter_sr_cry_5\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_6_LC_21_27_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48654\,
            in1 => \N__48355\,
            in2 => \_gnd_net_\,
            in3 => \N__48333\,
            lcout => \serializer_mod_inst.counter_srZ0Z_6\,
            ltout => OPEN,
            carryin => \serializer_mod_inst.counter_sr_cry_5\,
            carryout => \serializer_mod_inst.counter_sr_cry_6\,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \serializer_mod_inst.counter_sr_7_LC_21_27_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__48641\,
            in1 => \N__48618\,
            in2 => \_gnd_net_\,
            in3 => \N__48621\,
            lcout => \serializer_mod_inst.counter_srZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65754\,
            ce => \N__48600\,
            sr => \N__62827\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_15_LC_22_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__57524\,
            in2 => \_gnd_net_\,
            in3 => \N__59708\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_24_LC_22_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59712\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61113\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_16_LC_22_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59709\,
            in2 => \_gnd_net_\,
            in3 => \N__57627\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_25_LC_22_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59713\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60981\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_17_LC_22_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59710\,
            in2 => \_gnd_net_\,
            in3 => \N__57413\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_26_LC_22_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60897\,
            lcout => \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.c_data_system_o_2Z0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_18_LC_22_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59711\,
            in2 => \_gnd_net_\,
            in3 => \N__59865\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_27_LC_22_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__60786\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65568\,
            ce => \N__48726\,
            sr => \N__62955\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_19_LC_22_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61645\,
            in2 => \_gnd_net_\,
            in3 => \N__59593\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65580\,
            ce => \N__48725\,
            sr => \N__62952\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_28_LC_22_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59596\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62367\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65580\,
            ce => \N__48725\,
            sr => \N__62952\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_29_LC_22_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__62262\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59597\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf5_c_data_system_o_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65580\,
            ce => \N__48725\,
            sr => \N__62952\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_0_LC_22_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59595\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61943\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65580\,
            ce => \N__48725\,
            sr => \N__62952\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf5.c_data_system_o_7_LC_22_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63482\,
            in2 => \_gnd_net_\,
            in3 => \N__59594\,
            lcout => cemf_module_64ch_ctrl_inst1_data_interrupts_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65580\,
            ce => \N__48725\,
            sr => \N__62952\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI23RI1_LC_22_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55228\,
            in1 => \N__55455\,
            in2 => \N__48677\,
            in3 => \N__48694\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIL86H2_LC_22_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100001101"
        )
    port map (
            in0 => \N__48670\,
            in1 => \N__55057\,
            in2 => \N__48701\,
            in3 => \N__54832\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_19_LC_22_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61646\,
            in2 => \_gnd_net_\,
            in3 => \N__59599\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65591\,
            ce => \N__49095\,
            sr => \N__62947\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIE2FN1_LC_22_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55454\,
            in1 => \N__55229\,
            in2 => \N__48914\,
            in3 => \N__48934\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_0_LC_22_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__61969\,
            in2 => \_gnd_net_\,
            in3 => \N__59598\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65591\,
            ce => \N__49095\,
            sr => \N__62947\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI18QL2_LC_22_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__54833\,
            in1 => \N__48935\,
            in2 => \N__55062\,
            in3 => \N__48910\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQL7_LC_22_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100111111"
        )
    port map (
            in0 => \N__54006\,
            in1 => \N__48891\,
            in2 => \N__48885\,
            in3 => \N__58223\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI8TQLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIJ0CO7_LC_22_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53718\,
            in1 => \_gnd_net_\,
            in2 => \N__48882\,
            in3 => \N__48879\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNI01RI1_LC_22_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55263\,
            in1 => \N__55445\,
            in2 => \N__48867\,
            in3 => \N__49156\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNIJ66H2_LC_22_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111101000101"
        )
    port map (
            in0 => \N__48866\,
            in1 => \N__55058\,
            in2 => \N__49163\,
            in3 => \N__54837\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579D7_LC_22_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53962\,
            in1 => \N__51395\,
            in2 => \N__48837\,
            in3 => \N__48834\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNI579DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIGAQF7_LC_22_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53716\,
            in2 => \N__48828\,
            in3 => \N__48825\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18_LC_22_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__48819\,
            in2 => \N__48813\,
            in3 => \N__55745\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net\,
            ce => \N__55559\,
            sr => \N__62941\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9D7_LC_22_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53948\,
            in1 => \N__51476\,
            in2 => \N__48810\,
            in3 => \N__48801\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIAC9DZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNILFQF7_LC_22_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53717\,
            in1 => \_gnd_net_\,
            in2 => \N__49209\,
            in3 => \N__49206\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_19_LC_22_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55746\,
            in1 => \_gnd_net_\,
            in2 => \N__49200\,
            in3 => \N__49197\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_18C_net\,
            ce => \N__55559\,
            sr => \N__62941\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_18_LC_22_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59505\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59853\,
            lcout => cemf_module_64ch_ctrl_inst1_data_clkctrovf_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65611\,
            ce => \N__49094\,
            sr => \N__62936\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_27_LC_22_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59504\,
            in2 => \_gnd_net_\,
            in3 => \N__60806\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65611\,
            ce => \N__49094\,
            sr => \N__62936\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_28_LC_22_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59506\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62356\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65611\,
            ce => \N__49094\,
            sr => \N__62936\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf3.c_data_system_o_29_LC_22_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__62263\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59507\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf3_c_data_system_o_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65611\,
            ce => \N__49094\,
            sr => \N__62936\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI06692_17_LC_22_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__57926\,
            in1 => \N__58184\,
            in2 => \N__49008\,
            in3 => \N__51241\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLH5_LC_22_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60598\,
            in1 => \N__48975\,
            in2 => \N__48945\,
            in3 => \N__49437\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNISFLHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNITTFV5_LC_22_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60379\,
            in1 => \_gnd_net_\,
            in2 => \N__49572\,
            in3 => \N__49569\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23_LC_22_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49503\,
            in2 => \N__49563\,
            in3 => \N__60196\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.dout_conf\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net\,
            ce => \N__60023\,
            sr => \N__62927\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIOOFV5_LC_22_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__60378\,
            in1 => \N__49527\,
            in2 => \N__49539\,
            in3 => \_gnd_net_\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_22_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_22_LC_22_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49521\,
            in2 => \N__49506\,
            in3 => \N__60195\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_23C_net\,
            ce => \N__60023\,
            sr => \N__62927\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIOQSI1_LC_22_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__55453\,
            in1 => \N__55156\,
            in2 => \N__49493\,
            in3 => \N__49454\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI81C92_17_LC_22_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__58182\,
            in1 => \N__57989\,
            in2 => \N__49431\,
            in3 => \N__49378\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOR392_17_LC_22_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__57990\,
            in1 => \N__58183\,
            in2 => \N__49339\,
            in3 => \N__49308\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFH5_LC_22_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60618\,
            in1 => \N__49268\,
            in2 => \N__49233\,
            in3 => \N__49230\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI8MFHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI94AV5_LC_22_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60377\,
            in1 => \_gnd_net_\,
            in2 => \N__49218\,
            in3 => \N__49215\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10_LC_22_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60193\,
            in1 => \_gnd_net_\,
            in2 => \N__49860\,
            in3 => \N__49758\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net\,
            ce => \N__60022\,
            sr => \N__62919\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044Q5_LC_22_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60617\,
            in1 => \N__49832\,
            in2 => \N__49803\,
            in3 => \N__49791\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI044QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI1IU76_LC_22_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60376\,
            in2 => \N__49785\,
            in3 => \N__49782\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_9_LC_22_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49776\,
            in2 => \N__49761\,
            in3 => \N__60194\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_10C_net\,
            ce => \N__60022\,
            sr => \N__62919\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIQIB92_17_LC_22_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58013\,
            in1 => \N__58110\,
            in2 => \N__53793\,
            in3 => \N__49751\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNISKB92_17_LC_22_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58111\,
            in1 => \N__58014\,
            in2 => \N__49718\,
            in3 => \N__49677\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253Q5_LC_22_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60605\,
            in1 => \N__49637\,
            in2 => \N__49599\,
            in3 => \N__49596\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI253QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI3JT76_LC_22_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60374\,
            in2 => \N__49581\,
            in3 => \N__49578\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3_LC_22_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__49905\,
            in2 => \N__49986\,
            in3 => \N__60167\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net\,
            ce => \N__60018\,
            sr => \N__62911\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2Q5_LC_22_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60612\,
            in1 => \N__49961\,
            in2 => \N__49935\,
            in3 => \N__49926\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNITV2QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIUDT76_LC_22_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60375\,
            in1 => \_gnd_net_\,
            in2 => \N__49917\,
            in3 => \N__49914\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_2_LC_22_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60166\,
            in1 => \_gnd_net_\,
            in2 => \N__49908\,
            in3 => \N__60657\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_3C_net\,
            ce => \N__60018\,
            sr => \N__62911\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_2_LC_22_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101001100"
        )
    port map (
            in0 => \N__54403\,
            in1 => \N__56726\,
            in2 => \N__50196\,
            in3 => \N__56447\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_6_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_2_LC_22_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__50218\,
            in1 => \N__50611\,
            in2 => \N__49893\,
            in3 => \N__50050\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65662\,
            ce => 'H',
            sr => \N__65004\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_3_LC_22_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111011110000000"
        )
    port map (
            in0 => \N__50051\,
            in1 => \N__50219\,
            in2 => \N__54231\,
            in3 => \N__55943\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65662\,
            ce => 'H',
            sr => \N__65004\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_15_LC_22_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110101"
        )
    port map (
            in0 => \N__56725\,
            in1 => \N__50015\,
            in2 => \N__54405\,
            in3 => \N__49890\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_15_LC_22_17_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000011110000"
        )
    port map (
            in0 => \N__50140\,
            in1 => \N__50175\,
            in2 => \N__49878\,
            in3 => \N__56446\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_1_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_1_LC_22_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010110011001100"
        )
    port map (
            in0 => \N__54237\,
            in1 => \N__55964\,
            in2 => \N__50220\,
            in3 => \N__50049\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65662\,
            ce => 'H',
            sr => \N__65004\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_3_LC_22_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50191\,
            in2 => \_gnd_net_\,
            in3 => \N__54398\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1593_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIMJR28_26_LC_22_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__55864\,
            in1 => \N__56448\,
            in2 => \N__50169\,
            in3 => \N__50139\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_842_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIJU6F7_23_LC_22_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__50016\,
            in1 => \N__54404\,
            in2 => \_gnd_net_\,
            in3 => \N__56718\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_267\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_267_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAOTPE_26_LC_22_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000001"
        )
    port map (
            in0 => \N__50154\,
            in1 => \N__56439\,
            in2 => \N__50148\,
            in3 => \N__50141\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_321_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIIC372_3_LC_22_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__54251\,
            in1 => \N__56056\,
            in2 => \_gnd_net_\,
            in3 => \N__54342\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_a3_1_1_i_m2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIDH244_3_LC_22_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100000100"
        )
    port map (
            in0 => \N__54343\,
            in1 => \N__54419\,
            in2 => \N__50019\,
            in3 => \N__56130\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_101\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_2_LC_22_18_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110000000000"
        )
    port map (
            in0 => \N__49997\,
            in1 => \N__56360\,
            in2 => \N__64737\,
            in3 => \N__55929\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1802\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_0_2_LC_22_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__50714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66118\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_904\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_0_LC_22_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__56358\,
            in1 => \_gnd_net_\,
            in2 => \N__66155\,
            in3 => \N__64420\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_1_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_0_LC_22_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000101"
        )
    port map (
            in0 => \N__56512\,
            in1 => \N__50551\,
            in2 => \N__50469\,
            in3 => \N__57209\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3TI11_2_LC_22_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__56357\,
            in1 => \_gnd_net_\,
            in2 => \N__66154\,
            in3 => \N__50715\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_316_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_7_14_LC_22_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64316\,
            in2 => \N__50466\,
            in3 => \N__64265\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_372_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_14_LC_22_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__50581\,
            in1 => \N__50226\,
            in2 => \N__50463\,
            in3 => \N__50460\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_412_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_14_LC_22_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101110111011"
        )
    port map (
            in0 => \N__50766\,
            in1 => \N__50427\,
            in2 => \N__50418\,
            in3 => \N__50415\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65688\,
            ce => 'H',
            sr => \N__65013\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_14_LC_22_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101111111"
        )
    port map (
            in0 => \N__56359\,
            in1 => \N__56511\,
            in2 => \N__50386\,
            in3 => \N__64421\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_0_o2_1_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_25_LC_22_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__50923\,
            in1 => \N__50631\,
            in2 => \N__57014\,
            in3 => \N__66453\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65703\,
            ce => 'H',
            sr => \N__65021\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_RNISQP11_2_LC_22_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__65852\,
            in1 => \N__50666\,
            in2 => \N__65932\,
            in3 => \N__66020\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_87_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9FLC_24_LC_22_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50921\,
            in2 => \_gnd_net_\,
            in3 => \N__57029\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1596_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_25_LC_22_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__66560\,
            in1 => \N__57002\,
            in2 => \N__50634\,
            in3 => \N__66691\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_24_LC_22_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101111"
        )
    port map (
            in0 => \N__66608\,
            in1 => \N__50922\,
            in2 => \N__57013\,
            in3 => \N__57030\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_24_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_24_LC_22_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0100111100001111"
        )
    port map (
            in0 => \N__50621\,
            in1 => \N__50585\,
            in2 => \N__50565\,
            in3 => \N__55920\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65703\,
            ce => 'H',
            sr => \N__65021\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_14_LC_22_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__65926\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__66021\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_86_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_11_LC_22_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66093\,
            in2 => \_gnd_net_\,
            in3 => \N__66554\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_0_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_11_LC_22_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000001000000"
        )
    port map (
            in0 => \N__50717\,
            in1 => \N__50538\,
            in2 => \N__50562\,
            in3 => \N__64788\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_11_LC_22_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001100000"
        )
    port map (
            in0 => \N__50539\,
            in1 => \N__66680\,
            in2 => \N__50493\,
            in3 => \N__66503\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_1_LC_22_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50727\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_14_LC_22_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__66105\,
            in1 => \N__65848\,
            in2 => \N__50775\,
            in3 => \N__50667\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_95_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_0_LC_22_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50757\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.stop_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_RNI3DKR_2_LC_22_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__50716\,
            in2 => \_gnd_net_\,
            in3 => \N__66094\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_844_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_2_LC_22_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50655\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65720\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_i_o2_LC_22_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__51080\,
            in1 => \N__51044\,
            in2 => \N__51024\,
            in3 => \N__51122\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1594_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_1_LC_22_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57642\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_2_LC_22_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50649\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_1_LC_22_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51129\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQUIH_10_LC_22_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66095\,
            in2 => \_gnd_net_\,
            in3 => \N__64787\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1754_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.stop_q_2_LC_22_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51213\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_stop_q_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.scl_q_0_LC_22_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51206\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.scl_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65729\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6_0_a2_LC_22_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__51123\,
            in1 => \N__51081\,
            in2 => \N__51053\,
            in3 => \N__51022\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_no_restart6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_0_LC_22_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50993\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_1_LC_22_23_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__50955\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_q_2_LC_22_23_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50949\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.load_wdata_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_1_LC_22_23_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__66383\,
            in1 => \N__66789\,
            in2 => \N__66693\,
            in3 => \N__66412\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_2_LC_22_23_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__51309\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_q_0_LC_22_23_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__50882\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.start_I2C_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65739\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_6_0_LC_22_23_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000001"
        )
    port map (
            in0 => \N__66790\,
            in1 => \N__66382\,
            in2 => \N__66419\,
            in3 => \N__66504\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_122_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_1_LC_22_24_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51285\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_q_0_LC_22_24_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__51303\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.r_w_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65747\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_18_LC_23_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59672\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59864\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_18,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65581\,
            ce => \N__54123\,
            sr => \N__62958\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_27_LC_23_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59675\,
            in2 => \_gnd_net_\,
            in3 => \N__60787\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65581\,
            ce => \N__54123\,
            sr => \N__62958\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_19_LC_23_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59673\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61631\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65581\,
            ce => \N__54123\,
            sr => \N__62958\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_25_LC_23_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__60980\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__59676\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65581\,
            ce => \N__54123\,
            sr => \N__62958\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_29_LC_23_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__62246\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65581\,
            ce => \N__54123\,
            sr => \N__62958\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_23_LC_23_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59671\,
            in2 => \_gnd_net_\,
            in3 => \N__61242\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_23,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65581\,
            ce => \N__54123\,
            sr => \N__62958\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HH5_LC_23_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__57319\,
            in1 => \N__60614\,
            in2 => \N__51447\,
            in3 => \N__51543\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIL4HHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIMIBV5_LC_23_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60385\,
            in1 => \_gnd_net_\,
            in2 => \N__51537\,
            in3 => \N__51534\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_19_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19_LC_23_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60207\,
            in1 => \_gnd_net_\,
            in2 => \N__51528\,
            in3 => \N__51315\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net\,
            ce => \N__60017\,
            sr => \N__62956\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIAE492_17_LC_23_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__58006\,
            in1 => \N__58199\,
            in2 => \N__51506\,
            in3 => \N__51463\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI8C492_17_LC_23_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58200\,
            in1 => \N__58007\,
            in2 => \N__51430\,
            in3 => \N__51382\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGH5_LC_23_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60613\,
            in1 => \N__51369\,
            in2 => \N__51342\,
            in3 => \N__51339\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIGVGHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIHDBV5_LC_23_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60384\,
            in2 => \N__51327\,
            in3 => \N__51324\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_18_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_18_LC_23_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53535\,
            in2 => \N__51318\,
            in3 => \N__60206\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_19C_net\,
            ce => \N__60017\,
            sr => \N__62956\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_1_25_LC_23_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011101110111"
        )
    port map (
            in0 => \N__53340\,
            in1 => \N__53266\,
            in2 => \N__53034\,
            in3 => \N__53009\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_4_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_4_25_LC_23_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__52803\,
            in1 => \N__52782\,
            in2 => \N__52548\,
            in3 => \N__52525\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_1_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_0_25_LC_23_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__52254\,
            in2 => \N__52239\,
            in3 => \N__52235\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_3_25_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_25_LC_23_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__51984\,
            in1 => \N__51975\,
            in2 => \N__51969\,
            in3 => \N__51663\,
            lcout => \I2C_top_level_inst1_s_data_oreg_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65604\,
            ce => \N__54495\,
            sr => \N__65024\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_RNO_3_25_LC_23_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__51966\,
            in1 => \N__51923\,
            in2 => \N__51684\,
            in3 => \N__51672\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_data32_1_6_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI48492_17_LC_23_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58196\,
            in1 => \N__57991\,
            in2 => \N__51656\,
            in3 => \N__54193\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNI6A492_17_LC_23_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__57992\,
            in1 => \N__58197\,
            in2 => \N__51620\,
            in3 => \N__54142\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGH5_LC_23_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__51587\,
            in1 => \N__60590\,
            in2 => \N__51555\,
            in3 => \N__51552\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIBQGHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIC8BV5_LC_23_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60383\,
            in2 => \N__53547\,
            in3 => \N__53544\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_17_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17_LC_23_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60163\,
            in1 => \_gnd_net_\,
            in2 => \N__53538\,
            in3 => \N__53454\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net\,
            ce => \N__60016\,
            sr => \N__62948\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGH5_LC_23_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60589\,
            in1 => \N__53526\,
            in2 => \N__53496\,
            in3 => \N__53481\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNI6LGHZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNI73BV5_LC_23_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60382\,
            in1 => \_gnd_net_\,
            in2 => \N__53475\,
            in3 => \N__53472\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_16_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_16_LC_23_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \N__53466\,
            in1 => \_gnd_net_\,
            in2 => \N__53457\,
            in3 => \N__60162\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_17C_net\,
            ce => \N__60016\,
            sr => \N__62948\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_31_LC_23_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62059\,
            in2 => \_gnd_net_\,
            in3 => \N__59602\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_14_LC_23_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59603\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__58489\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_14,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_0_LC_23_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59607\,
            in2 => \_gnd_net_\,
            in3 => \N__61968\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_15_LC_23_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59604\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57534\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_15,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_24_LC_23_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59600\,
            in2 => \_gnd_net_\,
            in3 => \N__61124\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_16_LC_23_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59605\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57628\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_16,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_28_LC_23_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59601\,
            in2 => \_gnd_net_\,
            in3 => \N__62357\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf1_c_data_system_o_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf1.c_data_system_o_17_LC_23_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59606\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__57418\,
            lcout => cemf_module_64ch_ctrl_inst1_data_config_17,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65625\,
            ce => \N__54118\,
            sr => \N__62942\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RL7_LC_23_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53992\,
            in1 => \N__57801\,
            in2 => \N__54048\,
            in3 => \N__54576\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNID2RLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNIO5CO7_LC_23_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__53719\,
            in2 => \N__54030\,
            in3 => \N__54027\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1_LC_23_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__54021\,
            in2 => \N__54009\,
            in3 => \N__55740\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net\,
            ce => \N__55572\,
            sr => \N__62937\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RL7_LC_23_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__53991\,
            in1 => \N__53788\,
            in2 => \N__53745\,
            in3 => \N__53730\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNII7RLZ0Z7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_7_RNITACO7_LC_23_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__53720\,
            in1 => \_gnd_net_\,
            in2 => \N__55755\,
            in3 => \N__55752\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_2_LC_23_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__55741\,
            in1 => \_gnd_net_\,
            in2 => \N__55596\,
            in3 => \N__55593\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_dataZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.ser_data_1C_net\,
            ce => \N__55572\,
            sr => \N__62937\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_5_RNIG4FN1_LC_23_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010111011"
        )
    port map (
            in0 => \N__55452\,
            in1 => \N__54634\,
            in2 => \N__55192\,
            in3 => \N__54598\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.c_state_ret_3_RNI3AQL2_LC_23_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__55054\,
            in1 => \N__54825\,
            in2 => \N__54638\,
            in3 => \N__54599\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_b.spi_conf_inst1.data_1_iv_i_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_data32_26_LC_23_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__54570\,
            in1 => \N__54558\,
            in2 => \N__54546\,
            in3 => \N__64266\,
            lcout => \I2C_top_level_inst1_s_data_oreg_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65651\,
            ce => \N__54494\,
            sr => \N__65010\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNIBPUN4_3_LC_23_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__54423\,
            in1 => \N__54380\,
            in2 => \_gnd_net_\,
            in3 => \N__54344\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_230\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_230_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_1_LC_23_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__56145\,
            in1 => \N__54258\,
            in2 => \N__54240\,
            in3 => \N__56727\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNO_0_3_LC_23_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__56728\,
            in1 => \N__56146\,
            in2 => \N__56040\,
            in3 => \N__56070\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_err_state_2_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNII6J06_8_LC_23_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__56144\,
            in1 => \N__56069\,
            in2 => \_gnd_net_\,
            in3 => \N__56036\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1604_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_4_LC_23_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__62402\,
            in2 => \N__56013\,
            in3 => \N__66174\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_365_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_4_LC_23_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111010111010101"
        )
    port map (
            in0 => \N__56010\,
            in1 => \N__55869\,
            in2 => \N__55998\,
            in3 => \N__55800\,
            lcout => \I2C_top_level_inst1_I2C_Interpreter_inst_c_state_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65663\,
            ce => 'H',
            sr => \N__65001\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQQ5F_13_LC_23_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__56248\,
            in1 => \N__64705\,
            in2 => \N__56353\,
            in3 => \N__56560\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.un1_c_state_4_0_a2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI4NN21_13_LC_23_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__55995\,
            in3 => \N__64496\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_676_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIFO0G5_7_LC_23_17_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__55761\,
            in1 => \N__55767\,
            in2 => \N__55992\,
            in3 => \N__55875\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_address\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_err_state_RNISM8F1_3_LC_23_17_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010011001100"
        )
    port map (
            in0 => \N__55960\,
            in1 => \N__56336\,
            in2 => \N__55944\,
            in3 => \N__55928\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_2_sqmuxa_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI05EA2_7_LC_23_17_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000101010"
        )
    port map (
            in0 => \N__64704\,
            in1 => \N__55863\,
            in2 => \N__57291\,
            in3 => \N__55795\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1565_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIF5IJ_13_LC_23_17_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56247\,
            in2 => \_gnd_net_\,
            in3 => \N__66244\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_799_0_i_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_16_LC_23_17_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__56660\,
            in2 => \N__56364\,
            in3 => \N__57208\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_115\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_7_0_LC_23_18_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__65897\,
            in1 => \N__64706\,
            in2 => \N__57015\,
            in3 => \N__56350\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_6_0_LC_23_18_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__64707\,
            in1 => \N__62472\,
            in2 => \_gnd_net_\,
            in3 => \N__56351\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_5_0_LC_23_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__66290\,
            in1 => \N__64802\,
            in2 => \_gnd_net_\,
            in3 => \N__64407\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_0_LC_23_18_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__56748\,
            in1 => \N__56853\,
            in2 => \N__56283\,
            in3 => \N__56280\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_0_LC_23_18_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100110011001100"
        )
    port map (
            in0 => \N__56274\,
            in1 => \N__56262\,
            in2 => \N__56253\,
            in3 => \N__57132\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65689\,
            ce => 'H',
            sr => \N__65014\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIASHJ_14_LC_23_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__64406\,
            in1 => \N__56700\,
            in2 => \N__57216\,
            in3 => \N__56441\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_691\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_23_LC_23_19_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__66251\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__56249\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_a3_0_23_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_23_LC_23_19_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110101111"
        )
    port map (
            in0 => \N__66166\,
            in1 => \N__56180\,
            in2 => \N__56154\,
            in3 => \N__56559\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_0_i_0_0_0_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIAAHD_16_LC_23_19_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__56649\,
            in1 => \N__64457\,
            in2 => \_gnd_net_\,
            in3 => \N__57736\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_288\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_288_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9QGJ_23_LC_23_19_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__56742\,
            in3 => \N__56701\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_231\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_23_LC_23_19_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001110110011"
        )
    port map (
            in0 => \N__57012\,
            in1 => \N__56739\,
            in2 => \N__66449\,
            in3 => \N__66692\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65704\,
            ce => 'H',
            sr => \N__65022\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_16_LC_23_19_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000100000000"
        )
    port map (
            in0 => \N__66167\,
            in1 => \N__56670\,
            in2 => \N__57227\,
            in3 => \N__56627\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65704\,
            ce => 'H',
            sr => \N__65022\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_1_LC_23_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000001010"
        )
    port map (
            in0 => \N__56650\,
            in1 => \_gnd_net_\,
            in2 => \N__56631\,
            in3 => \N__66168\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65704\,
            ce => 'H',
            sr => \N__65022\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_3_LC_23_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000111110001000"
        )
    port map (
            in0 => \N__64458\,
            in1 => \N__56516\,
            in2 => \N__56493\,
            in3 => \N__56468\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65704\,
            ce => 'H',
            sr => \N__65022\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI046R_4_LC_23_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__56442\,
            in1 => \N__56908\,
            in2 => \N__56844\,
            in3 => \N__56946\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.un30_i_a2_9_a2_4_a2_0_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNISICG1_25_LC_23_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__56994\,
            in1 => \N__57056\,
            in2 => \N__56379\,
            in3 => \N__64686\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1446_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIPVAM1_12_LC_23_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__57060\,
            in3 => \N__56885\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI59N81_25_LC_23_20_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__56993\,
            in1 => \N__56770\,
            in2 => \N__57057\,
            in3 => \N__64685\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un40_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIKLID_24_LC_23_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__57028\,
            in1 => \N__66019\,
            in2 => \_gnd_net_\,
            in3 => \N__65978\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_232\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_232_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBFN81_25_LC_23_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__56995\,
            in1 => \N__56964\,
            in2 => \N__56955\,
            in3 => \N__64687\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_a2_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIQ47E3_25_LC_23_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__56771\,
            in1 => \N__57124\,
            in2 => \N__56952\,
            in3 => \N__57082\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_o2_1_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_4_0_LC_23_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__56947\,
            in1 => \N__56909\,
            in2 => \N__66333\,
            in3 => \N__56886\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_a2_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_0_LC_23_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__57255\,
            in1 => \N__57066\,
            in2 => \N__56757\,
            in3 => \N__57300\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65730\,
            ce => 'H',
            sr => \N__65025\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_8_0_LC_23_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__66779\,
            in1 => \N__56843\,
            in2 => \N__64801\,
            in3 => \N__56829\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_3_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_0_LC_23_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__56787\,
            in1 => \N__57146\,
            in2 => \N__56778\,
            in3 => \N__56775\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_212\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_0_LC_23_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__66780\,
            in1 => \_gnd_net_\,
            in2 => \N__57147\,
            in3 => \N__65800\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_2_LC_23_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010011110111"
        )
    port map (
            in0 => \N__65819\,
            in1 => \N__66493\,
            in2 => \N__65807\,
            in3 => \N__57744\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1653_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_2_LC_23_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010000000000"
        )
    port map (
            in0 => \N__57753\,
            in1 => \N__66675\,
            in2 => \N__57294\,
            in3 => \N__66699\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65730\,
            ce => 'H',
            sr => \N__65025\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_0_LC_23_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__66548\,
            in1 => \N__66653\,
            in2 => \_gnd_net_\,
            in3 => \N__66492\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_255_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_0_LC_23_22_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000001010"
        )
    port map (
            in0 => \N__66851\,
            in1 => \N__66674\,
            in2 => \N__57267\,
            in3 => \N__66559\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_208\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNI9PI7_14_LC_23_22_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100010001"
        )
    port map (
            in0 => \N__57223\,
            in1 => \N__64425\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1601_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNI6FAA_0_LC_23_22_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__57150\,
            in3 => \N__66497\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_239\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_239_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_0_LC_23_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010000"
        )
    port map (
            in0 => \N__66788\,
            in1 => \N__66411\,
            in2 => \N__57135\,
            in3 => \N__66378\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_a3_1_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_0_LC_23_22_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__57131\,
            in1 => \N__57705\,
            in2 => \N__57093\,
            in3 => \N__57090\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_2_2_LC_23_22_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__66673\,
            in1 => \N__66431\,
            in2 => \_gnd_net_\,
            in3 => \N__65783\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1776\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNINS3G1_8_LC_23_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__66410\,
            in1 => \N__66377\,
            in2 => \_gnd_net_\,
            in3 => \N__66787\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_90_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_5_0_LC_23_22_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__66498\,
            in1 => \N__66850\,
            in2 => \N__57747\,
            in3 => \N__57743\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_209\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_q_0_LC_23_23_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__57686\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.sda_i_qZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65748\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16_LC_24_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63341\,
            in1 => \N__57435\,
            in2 => \_gnd_net_\,
            in3 => \N__57620\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net\,
            ce => \N__63030\,
            sr => \N__62959\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_15_LC_24_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58386\,
            in1 => \N__63342\,
            in2 => \_gnd_net_\,
            in3 => \N__57496\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net\,
            ce => \N__63030\,
            sr => \N__62959\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_17_LC_24_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__57429\,
            in1 => \N__63343\,
            in2 => \_gnd_net_\,
            in3 => \N__57419\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_16C_net\,
            ce => \N__63030\,
            sr => \N__62959\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_19_LC_24_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__59652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61640\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_19,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65613\,
            ce => \N__58884\,
            sr => \N__62957\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_29_LC_24_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__59651\,
            in2 => \_gnd_net_\,
            in3 => \N__62260\,
            lcout => \cemf_module_64ch_ctrl_inst1_top_cemf_module_64ch_reg_inst_I2C_Register_conf2_c_data_system_o_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65613\,
            ce => \N__58884\,
            sr => \N__62957\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.I2C_Register_conf2.c_data_system_o_0_LC_24_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0100010001000100"
        )
    port map (
            in0 => \N__59653\,
            in1 => \N__61959\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => cemf_module_64ch_ctrl_inst1_data_coarseovf_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65613\,
            ce => \N__58884\,
            sr => \N__62957\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10_LC_24_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58818\,
            in1 => \N__63353\,
            in2 => \_gnd_net_\,
            in3 => \N__58795\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\,
            ce => \N__63025\,
            sr => \N__62953\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_11_LC_24_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63352\,
            in1 => \N__58707\,
            in2 => \_gnd_net_\,
            in3 => \N__58684\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\,
            ce => \N__63025\,
            sr => \N__62953\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_12_LC_24_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58602\,
            in1 => \N__63354\,
            in2 => \_gnd_net_\,
            in3 => \N__58592\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\,
            ce => \N__63025\,
            sr => \N__62953\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_14_LC_24_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__58263\,
            in1 => \N__63355\,
            in2 => \_gnd_net_\,
            in3 => \N__58473\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\,
            ce => \N__63025\,
            sr => \N__62953\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_13_LC_24_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__58348\,
            in1 => \_gnd_net_\,
            in2 => \N__63376\,
            in3 => \N__58269\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_10C_net\,
            ce => \N__63025\,
            sr => \N__62953\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIMEB92_17_LC_24_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000101011001111"
        )
    port map (
            in0 => \N__57987\,
            in1 => \N__58180\,
            in2 => \N__58257\,
            in3 => \N__58211\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_0_RNIOGB92_17_LC_24_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110010101111"
        )
    port map (
            in0 => \N__58181\,
            in1 => \N__57988\,
            in2 => \N__57833\,
            in3 => \N__57799\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_iv_i_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2Q5_LC_24_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100111111111111"
        )
    port map (
            in0 => \N__60616\,
            in1 => \N__60714\,
            in2 => \N__60678\,
            in3 => \N__60675\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIOQ2QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIP8T76_LC_24_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__60387\,
            in2 => \N__60669\,
            in3 => \N__60666\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1_LC_24_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__60205\,
            in1 => \_gnd_net_\,
            in2 => \N__60660\,
            in3 => \N__60030\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net\,
            ce => \N__60024\,
            sr => \N__62949\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2Q5_LC_24_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111111111111"
        )
    port map (
            in0 => \N__60640\,
            in1 => \N__60615\,
            in2 => \N__60411\,
            in3 => \N__60393\,
            lcout => OPEN,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_11_RNIJL2QZ0Z5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.c_state_ret_13_RNIK3T76_LC_24_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__60386\,
            in1 => \_gnd_net_\,
            in2 => \N__60219\,
            in3 => \N__60216\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0\,
            ltout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.data_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_0_LC_24_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__60210\,
            in3 => \N__60204\,
            lcout => \cemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_dataZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVcemf_module_64ch_ctrl_inst1.spi_top_inst1.tdc_inst_a.spi_conf_inst1.ser_data_1C_net\,
            ce => \N__60024\,
            sr => \N__62949\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18_LC_24_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__59863\,
            in1 => \N__59763\,
            in2 => \_gnd_net_\,
            in3 => \N__63348\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_18\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_19_LC_24_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63344\,
            in1 => \N__59754\,
            in2 => \_gnd_net_\,
            in3 => \N__61647\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_20_LC_24_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__61551\,
            in1 => \N__61461\,
            in2 => \_gnd_net_\,
            in3 => \N__63349\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_21_LC_24_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63345\,
            in1 => \N__61455\,
            in2 => \_gnd_net_\,
            in3 => \N__61447\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_22_LC_24_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__61362\,
            in1 => \N__63350\,
            in2 => \_gnd_net_\,
            in3 => \N__61355\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_22\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_23_LC_24_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63346\,
            in1 => \N__61260\,
            in2 => \_gnd_net_\,
            in3 => \N__61229\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_24_LC_24_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__61137\,
            in1 => \N__63351\,
            in2 => \_gnd_net_\,
            in3 => \N__61130\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_24\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_25_LC_24_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63347\,
            in1 => \N__61026\,
            in2 => \_gnd_net_\,
            in3 => \N__61000\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_25\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_18C_net\,
            ce => \N__63003\,
            sr => \N__62943\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26_LC_24_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__60927\,
            in1 => \N__63298\,
            in2 => \_gnd_net_\,
            in3 => \N__60849\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_26\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_27_LC_24_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63295\,
            in1 => \N__60822\,
            in2 => \_gnd_net_\,
            in3 => \N__60798\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_27\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_28_LC_24_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__62382\,
            in1 => \N__63299\,
            in2 => \_gnd_net_\,
            in3 => \N__62368\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_29_LC_24_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63296\,
            in1 => \N__62271\,
            in2 => \_gnd_net_\,
            in3 => \N__62261\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_30_LC_24_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63300\,
            in1 => \N__62190\,
            in2 => \_gnd_net_\,
            in3 => \N__62169\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_31_LC_24_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63297\,
            in1 => \N__62079\,
            in2 => \_gnd_net_\,
            in3 => \N__62071\,
            lcout => \I2C_top_level_inst1.s_sda_o_reg\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_i_LC_24_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__63293\,
            in2 => \_gnd_net_\,
            in3 => \N__62421\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.un1_enable_desp_1_0_iZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_0_LC_24_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__63294\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__61970\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_26C_net\,
            ce => \N__63002\,
            sr => \N__62938\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1_LC_24_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__61878\,
            in1 => \N__63381\,
            in2 => \_gnd_net_\,
            in3 => \N__61872\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_2_LC_24_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63377\,
            in1 => \N__61752\,
            in2 => \_gnd_net_\,
            in3 => \N__61746\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_3_LC_24_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__63951\,
            in1 => \N__63382\,
            in2 => \_gnd_net_\,
            in3 => \N__63944\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_4_LC_24_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63378\,
            in1 => \N__63837\,
            in2 => \_gnd_net_\,
            in3 => \N__63826\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_5_LC_24_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__63708\,
            in1 => \N__63383\,
            in2 => \_gnd_net_\,
            in3 => \N__63701\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_6_LC_24_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63379\,
            in1 => \N__63591\,
            in2 => \_gnd_net_\,
            in3 => \N__63585\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_7_LC_24_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__63489\,
            in1 => \N__63384\,
            in2 => \_gnd_net_\,
            in3 => \N__63477\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_8_LC_24_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__63380\,
            in1 => \N__63156\,
            in2 => \_gnd_net_\,
            in3 => \N__63118\,
            lcout => \I2C_top_level_inst1.TX_Shift_Register_inst.c_data_inZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVI2C_top_level_inst1.TX_Shift_Register_inst.c_data_in_1C_net\,
            ce => \N__63015\,
            sr => \N__62928\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_LC_24_17_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011111111"
        )
    port map (
            in0 => \N__66866\,
            in1 => \N__66243\,
            in2 => \_gnd_net_\,
            in3 => \N__64605\,
            lcout => \I2C_top_level_inst1_s_burst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65690\,
            ce => 'H',
            sr => \N__65015\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_load_rdata2_LC_24_17_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011111111"
        )
    port map (
            in0 => \N__62420\,
            in1 => \N__64359\,
            in2 => \_gnd_net_\,
            in3 => \N__62480\,
            lcout => \I2C_top_level_inst1.s_load_rdata2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65690\,
            ce => 'H',
            sr => \N__65015\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIBMR9_7_LC_24_18_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__64712\,
            in1 => \N__66593\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1610_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_0_LC_24_18_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__64708\,
            in1 => \N__64629\,
            in2 => \N__64617\,
            in3 => \N__66561\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1609_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_address_RNO_0_0_LC_24_18_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000111000000"
        )
    port map (
            in0 => \N__64599\,
            in1 => \N__64551\,
            in2 => \N__64515\,
            in3 => \N__64497\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_address_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNIG0J7_19_LC_24_19_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__65892\,
            in2 => \_gnd_net_\,
            in3 => \N__66017\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_295\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_295_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_0_19_LC_24_19_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100011"
        )
    port map (
            in0 => \N__65991\,
            in1 => \N__64323\,
            in2 => \N__64476\,
            in3 => \N__64355\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_ns_i_i_1_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_no_restart_RNO_3_LC_24_20_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__64465\,
            in1 => \N__65893\,
            in2 => \N__64437\,
            in3 => \N__66326\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1386_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.load_rdata_q_RNI63VI_2_LC_24_20_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__66327\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__65933\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_81_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_3_19_LC_24_20_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__64344\,
            in1 => \N__66018\,
            in2 => \N__65987\,
            in3 => \N__66328\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_277\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \cemf_module_64ch_ctrl_inst1.top_cemf_module_64ch_reg_inst.pready_i_i2_i_i_o2_i_a2_LC_24_20_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__64299\,
            in2 => \_gnd_net_\,
            in3 => \N__64269\,
            lcout => OPEN,
            ltout => \N_73_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_1_19_LC_24_20_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000001000100"
        )
    port map (
            in0 => \N__66329\,
            in1 => \N__66291\,
            in2 => \N__66279\,
            in3 => \N__66255\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_274_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_19_LC_24_20_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__66201\,
            in1 => \N__65829\,
            in2 => \N__66195\,
            in3 => \N__66163\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_stateZ0Z_19\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65731\,
            ce => 'H',
            sr => \N__65026\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_state_RNO_2_19_LC_24_20_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__65985\,
            in1 => \N__65934\,
            in2 => \N__65898\,
            in3 => \N__65856\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_276\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_1_1_LC_24_21_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__66553\,
            in1 => \N__65820\,
            in2 => \N__65808\,
            in3 => \N__66687\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1669_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_1_LC_24_21_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000100000001100"
        )
    port map (
            in0 => \N__65787\,
            in1 => \N__64809\,
            in2 => \N__65772\,
            in3 => \N__64722\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.c_contZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__65740\,
            ce => 'H',
            sr => \N__65027\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_1_LC_24_21_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001000"
        )
    port map (
            in0 => \N__66853\,
            in1 => \N__66658\,
            in2 => \N__64824\,
            in3 => \N__66496\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_burst_RNO_3_LC_24_21_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__64790\,
            in1 => \N__64721\,
            in2 => \_gnd_net_\,
            in3 => \N__66549\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.un38_i_a2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIRCF5_0_LC_24_21_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66654\,
            in2 => \_gnd_net_\,
            in3 => \N__66494\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0\,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1607_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_3_2_LC_24_21_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66852\,
            in2 => \N__66825\,
            in3 => \N__66551\,
            lcout => OPEN,
            ltout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_0_2_LC_24_21_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010110000"
        )
    port map (
            in0 => \N__66552\,
            in1 => \N__66339\,
            in2 => \N__66822\,
            in3 => \N__66798\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.n_cont_i_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNIQ478_0_LC_24_21_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101000000000"
        )
    port map (
            in0 => \N__66495\,
            in1 => \_gnd_net_\,
            in2 => \N__66676\,
            in3 => \N__66550\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_80_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNISDF5_0_LC_24_22_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66555\,
            in2 => \_gnd_net_\,
            in3 => \N__66502\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1602_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \I2C_top_level_inst1.I2C_Interpreter_inst.c_cont_RNO_4_2_LC_24_22_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__66420\,
            in2 => \_gnd_net_\,
            in3 => \N__66384\,
            lcout => \I2C_top_level_inst1.I2C_Interpreter_inst.N_1666_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );
end \INTERFACE\;
